** sch_path: /home/ahmedreda/Project/AR_BGR/testbench/full_ldo/fullldox_v2-tb/noise.sch
**.subckt noise
vdd1 vdd1 vss 3.3 ac=1
.save i(vdd1)
vss2 vss GND 0
.save i(vss2)
Vbias net1 biasbgr 0
.save i(vbias)
vtot vdd1 vdd 0
.save i(vtot)
R2 net1 vdd 450000 m=1
R3 net2 vdd 300000 m=1
Vbiasldo net2 biasldo 0
.save i(vbiasldo)
C3 vo net3 47u m=1
R4 net3 vss 0.1 m=1
R5 vo net4 18 m=1
Vl net4 vss 0
.save i(vl)
x1 biasldo biasbgr vss vss vss vdd vss vss vss vss vss vss vss vss vss vss vss vss vo vdd vss fullldom

**** begin user architecture code


.options RSHUNT=1e15
.options savecurrents
.option TEMP=27
.option TNOM=27
.control
**set filetype=binary
set filetype=ascii
set color0=white
set color1=black
set color3=blue
set xbrushwidth=3
run
op
save all
noise v(vo) vdd1 dec 10 10 0.001MEG
setplot noise1
plot inoise_spectrum
plot onoise_spectrum


setplot noise2
print inoise_total onoise_total


.endc




.lib /home/ahmedreda/PDK/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include fullldom.spice




.GLOBAL GND
.end
