magic
tech sky130A
magscale 1 2
timestamp 1681430344
<< metal1 >>
rect -2978 8070 -1510 8102
rect -3058 7876 2974 8070
rect -32794 6460 -29382 7070
rect -3058 6764 -2880 7876
rect -1638 7570 2974 7876
rect -1638 6764 -1348 7570
rect -3058 6570 -1348 6764
rect -32656 6440 -29382 6460
rect 10698 160 14212 718
<< via1 >>
rect -2880 6764 -1638 7876
<< metal2 >>
rect -33230 20702 25682 23448
rect -2 20650 25660 20702
rect 10158 12476 24710 14948
rect -28390 8086 -28150 8252
rect -3058 7876 -1348 8070
rect -32794 6996 -29382 7070
rect -32794 6514 -32708 6996
rect -31874 6514 -29382 6996
rect -3058 6764 -2880 7876
rect -1638 6764 -1348 7876
rect -3058 6570 -1348 6764
rect -32794 6460 -29382 6514
rect -32656 6440 -29382 6460
rect -8544 6288 -7494 6402
rect -8544 6244 -8458 6288
rect -9478 6040 -8458 6244
rect -7546 6040 -7494 6288
rect -9478 6014 -7494 6040
rect -8544 5986 -7494 6014
rect -24838 5612 -24758 5760
rect -23784 5598 -23692 5776
rect -22718 5600 -22636 5760
rect -21660 5622 -21578 5762
rect -20602 5598 -20518 5760
rect -19546 5606 -19450 5762
rect -18478 5606 -18394 5734
rect -17426 5582 -17338 5694
rect 2300 4026 2928 4116
rect 2300 3666 2380 4026
rect 2854 3924 2928 4026
rect 2854 3830 6344 3924
rect 6840 3840 7204 3896
rect 2854 3666 2928 3830
rect 2300 3552 2928 3666
rect -24838 1998 -24756 2104
rect -23780 1998 -23698 2126
rect -22720 2000 -22638 2136
rect -21658 2002 -21578 2124
rect -20598 1998 -20516 2134
rect -19538 2000 -19456 2146
rect -18478 2002 -18396 2142
rect -17430 2002 -17308 2150
rect 5766 1720 5978 1834
<< via2 >>
rect -32708 6514 -31874 6996
rect -8458 6040 -7546 6288
rect 2380 3666 2854 4026
<< metal3 >>
rect -33230 20702 25682 23448
rect -2 20650 25660 20702
rect -32754 19396 -31750 20280
rect -32754 16476 -32644 19396
rect -31842 19246 -31750 19396
rect -31842 18592 -31802 19246
rect -31842 16554 -31750 18592
rect -31842 16476 -31768 16554
rect -32754 16416 -31768 16476
rect -32754 16024 -31876 16416
rect -32754 15818 -31768 16024
rect -32754 6996 -31750 15818
rect -5992 15602 -5796 15682
rect -2558 13200 1184 15070
rect 10158 12476 24710 14948
rect -2034 10756 -1214 10762
rect -5988 10702 -1214 10756
rect -5988 10076 -1976 10702
rect -1278 10076 -1214 10702
rect -5988 9980 -1214 10076
rect -5988 9978 -1826 9980
rect -32754 6514 -32708 6996
rect -31874 6514 -31750 6996
rect -32754 20 -31750 6514
rect -8544 6366 -7494 6402
rect -8544 6288 -8424 6366
rect -8544 6040 -8458 6288
rect -7538 6060 -7494 6366
rect -7546 6040 -7494 6060
rect -8544 5986 -7494 6040
rect 2300 4050 2928 4116
rect 2300 3604 2332 4050
rect 2884 3604 2928 4050
rect 2300 3552 2928 3604
<< via3 >>
rect -32644 16476 -31842 19396
rect -1976 10076 -1278 10702
rect -8424 6288 -7538 6366
rect -8424 6060 -7546 6288
rect -7546 6060 -7538 6288
rect 2332 4026 2884 4050
rect 2332 3666 2380 4026
rect 2380 3666 2854 4026
rect 2854 3666 2884 4026
rect 2332 3604 2884 3666
rect 1356 2664 1958 3222
<< metal4 >>
rect -33230 20702 25682 23448
rect -2 20650 25660 20702
rect -32804 20348 -31660 20364
rect -32804 20340 -30186 20348
rect -32828 19562 -30186 20340
rect -32828 19396 -31594 19562
rect -32828 16476 -32644 19396
rect -31842 17788 -31594 19396
rect -2044 19180 -1206 19186
rect -2452 18734 -1206 19180
rect -31842 17184 -30178 17788
rect -31842 16476 -31594 17184
rect -2028 16928 -1206 18734
rect -2048 16644 -1206 16928
rect -32828 15908 -31594 16476
rect -2436 16046 -1200 16644
rect -32774 15900 -31768 15908
rect -2028 10702 -1206 16046
rect 10158 12476 24710 14948
rect -2028 10076 -1976 10702
rect -1278 10076 -1206 10702
rect -2028 9978 -1206 10076
rect -8518 6800 -7522 6804
rect -8518 6366 2940 6800
rect -8518 6060 -8424 6366
rect -7538 6360 2940 6366
rect -7538 6060 -7522 6360
rect -8518 6006 -7522 6060
rect 2304 4906 2940 6360
rect 2300 4872 3994 4906
rect 2294 4856 3994 4872
rect 2294 4574 4000 4856
rect 2300 4530 4000 4574
rect 2304 4050 2940 4530
rect 2304 3604 2332 4050
rect 2884 3604 2940 4050
rect 3480 4138 4000 4530
rect 3480 4032 3972 4138
rect 2304 3524 2940 3604
rect 1262 3222 2112 3364
rect 1262 2664 1356 3222
rect 1958 2996 2112 3222
rect 1958 2774 4286 2996
rect 1958 2664 2112 2774
rect 1262 2554 2112 2664
use bandgapmd  bandgapmd_0
timestamp 1677883869
transform 1 0 -30388 0 1 20086
box -1026 -20046 30079 -4982
use cap_mim_m3_1_2x12  cap_mim_m3_1_2x12_0
timestamp 1681424555
transform 0 -1 -16304 1 0 17712
box -2492 -13920 2492 13920
use ldomc  ldomc_0
timestamp 1681424353
transform 1 0 2102 0 1 152
box -2078 -10 27574 23408
use sky130_fd_pr__cap_mim_m3_1_H9XL9H  sky130_fd_pr__cap_mim_m3_1_H9XL9H_0
timestamp 1681425679
transform 0 -1 3756 -1 0 3538
box -686 -540 686 540
<< labels >>
flabel metal1 13060 340 13402 520 0 FreeSans 4800 0 0 0 vss
port 4 nsew
flabel metal2 5822 1774 5890 1818 0 FreeSans 1600 0 0 0 biasldo
port 15 nsew
flabel metal2 -28338 8118 -28272 8198 0 FreeSans 800 0 0 0 biasbgr
port 20 nsew
flabel metal2 -24806 5688 -24796 5706 0 FreeSans 160 0 0 0 trim[0]
port 23 nsew
flabel metal2 -23760 5734 -23740 5750 0 FreeSans 160 0 0 0 trim[2]
port 26 nsew
flabel metal2 -22694 5704 -22670 5736 0 FreeSans 160 0 0 0 trim[4]
port 28 nsew
flabel metal2 -21626 5706 -21598 5740 0 FreeSans 160 0 0 0 trim[6]
port 30 nsew
flabel metal2 -20574 5708 -20544 5734 0 FreeSans 160 0 0 0 trim[8]
port 32 nsew
flabel metal2 -19512 5716 -19474 5750 0 FreeSans 160 0 0 0 trim[10]
port 34 nsew
flabel metal2 -18446 5670 -18428 5718 0 FreeSans 160 0 0 0 trim[12]
port 36 nsew
flabel metal2 -17406 5664 -17372 5682 0 FreeSans 160 0 0 0 trim[14]
port 38 nsew
flabel metal2 -17390 2020 -17374 2040 0 FreeSans 160 0 0 0 trim[15]
port 39 nsew
flabel metal2 -18450 2020 -18434 2040 0 FreeSans 160 0 0 0 trim[13]
port 41 nsew
flabel metal2 -19512 2016 -19492 2038 0 FreeSans 160 0 0 0 trim[11]
port 43 nsew
flabel metal2 -20568 2022 -20546 2044 0 FreeSans 160 0 0 0 trim[9]
port 45 nsew
flabel metal2 -21640 2020 -21626 2032 0 FreeSans 160 0 0 0 trim[7]
port 47 nsew
flabel metal2 -22696 2012 -22674 2032 0 FreeSans 160 0 0 0 trim[5]
port 49 nsew
flabel metal2 -23758 2012 -23734 2028 0 FreeSans 160 0 0 0 trim[3]
port 51 nsew
flabel metal2 -24806 2010 -24794 2022 0 FreeSans 160 0 0 0 trim[1]
port 53 nsew
flabel metal4 19218 21896 20338 22656 0 FreeSans 4800 0 0 0 vdd
port 54 nsew
flabel metal4 16746 13596 17486 14482 0 FreeSans 4800 0 0 0 out
port 56 nsew
<< end >>
