**.subckt dcsweep
vdd1 vdd1 vss 3.3
.save i(vdd1)
vss2 vss GND 0
.save i(vss2)
Vbias net1 biasbgr 0
.save i(vbias)
vtot vdd1 vdd 0
.save i(vtot)
R3 net4 vdd 300000 m=1
C3 vo net2 47u m=1
R4 net2 vss 0.1 m=1
R5 vo net3 1800 m=1
Vl net3 vss 0
.save i(vl)
Vbiasldo net4 biasldo 0
.save i(vbiasldo)
R2 net1 vdd 450000 m=1
**x1 vss vss vss vss vss vss vss vss vss vdd vss vss vss vss vss vss vss biasbgr vdd biasldo vo fullldoxcc

**x1 vo biasldo biasbgr vss vss vss vdd vss vss vss vss vss vss vss vss vss vss vss vss vss vdd fullldomcc

**x1 biasldo biasbgr vss vss vss vdd vss vss vss vss vss vss vss vss vss vss vss vss vo vdd vss fullldomf  -->no rc spice file


x1 biasldo biasbgr vss vss vss vdd vss vss vss vss vss vss vss vss vss vss vss vss vo vdd vss fullldom

**.subckt fullldom biasldo biasbgr trim[0] trim[2] trim[4] trim[6] trim[8] trim[10]
**+ trim[12] trim[14] trim[15] trim[13] trim[11] trim[9] trim[7] trim[5] trim[3] trim[1]
**+ out vdd vss



**** begin user architecture code


.lib /home/ahmedreda/PDK/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.include fullldom.spice


.options RSHUNT=1e15
.options savecurrents
.option TEMP=27
.option TNOM=27
.control
**set filetype=binary
set filetype=ascii
set color0=white
set color1=black
set color3=blue
set xbrushwidth=3
save all
OP
dc vdd1 0 5 0.1
meas DC vo_nom FIND vo AT=3.3

let ibias=vbias#branch
let itot=vtot#branch
let il=vl#branch
let ibldo=vbiasldo#branch

print  vo_nom
plot ibias itot il ibldo
plot vdd1 vo
plot vdd1-vo

meas DC vonom FIND vo AT=3.3
meas DC vo1 FIND vo AT=2.97
meas DC vo2 FIND vo AT=3.63
let lr=mag(vo1-vo2)/0.66
let lrPer=(mag(vo1-vo2)/0.66)*100

print lr
print lrPer

.endc



.GLOBAL GND
.end
