* NGSPICE file created from fullldom.ext - technology: sky130A

.subckt fullldom biasldo biasbgr trim[0] trim[2] trim[4] trim[6] trim[8] trim[10]
+ trim[12] trim[14] trim[15] trim[13] trim[11] trim[9] trim[7] trim[5] trim[3] trim[1]
+ out vdd vss
X0 vss.t210 vss.t207 vss.t209 vss.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1 vss.t84 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosrm_0.outn.t15 vss.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff vdd.t324 sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+13p pd=2.145e+08u as=0p ps=0u w=4e+06u l=1e+06u
X3 vdd.t98 ldomc_0.otaldom_0.pmosrm_0.out out.t65 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X4 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmosrm_0.outn vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.22e+12p pd=4.122e+07u as=4.64e+12p ps=3.896e+07u w=2e+06u l=4e+06u
X5 vss vss.t202 vss vss.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=3.712e+13p pd=2.9776e+08u as=0p ps=0u w=1e+06u l=1e+06u
X6 out.t64 ldomc_0.otaldom_0.pmosrm_0.out vdd vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4.5066e+14p ps=3.15498e+09u w=5e+07u l=500000u
X7 ldomc_0.otaldom_0.pcascodeupm_0.o1.t7 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t314 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.22e+12p ps=4.122e+07u w=2e+06u l=4e+06u
X8 vdd.t240 vdd.t238 vdd.t239 vdd.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=4.64e+12p pd=3.896e+07u as=5.22e+12p ps=4.122e+07u w=2e+06u l=4e+06u
X10 vss.t304 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosrm_0.outn vss.t303 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X11 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t82 vss.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X12 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t80 vss.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X13 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff vdd.t323 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X14 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t302 vss.t301 sky130_fd_pr__nfet_g5v0d10v5 ad=4.64e+12p pd=3.722e+07u as=0p ps=0u w=1e+06u l=1e+06u
X15 out.t63 ldomc_0.otaldom_0.pmosrm_0.out vdd.t96 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X16 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inp.t2 bandgapmd_0.otam_1.nmoslm_0.outp vdd.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+13p pd=2.145e+08u as=5.8e+12p ps=4.29e+07u w=4e+06u l=1e+06u
X17 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t78 vss.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X18 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff vdd.t248 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X19 bandgapmd_0.otam_1.nmosrm_0.outn.t33 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.pcsm_0.diff vdd.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X20 out.t66 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X21 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X22 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff vdd.t322 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X23 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 vdd.t313 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64e+12p pd=3.432e+07u as=8.12e+12p ps=6.006e+07u w=4e+06u l=1e+06u
X24 a_n7846_4436# bandgapmd_0.bg_stupm_0.vs2.t1 vdd.t139 vdd.t138 sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X25 vdd ldomc_0.otaldom_0.pmosrm_0.out out.t62 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X26 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t35 vdd.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64e+12p pd=3.664e+07u as=0p ps=0u w=2e+06u l=4e+06u
X27 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmosrm_0.outn vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X28 a_n24544_2674# a_n24956_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X29 ldomc_0.otaldom_0.nmosrm_0.outn bandgapmd_0.bg_pmosm_0.vbg.t3 ldomc_0.otaldom_0.pcsm_0.diff vdd.t283 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.29e+07u as=0p ps=0u w=4e+06u l=1e+06u
X30 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t175 vdd.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X31 vdd.t93 ldomc_0.otaldom_0.pmosrm_0.out out.t61 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X32 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X33 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t312 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X34 vdd.t92 ldomc_0.otaldom_0.pmosrm_0.out out.t60 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X35 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t272 sky130_fd_pr__pfet_g5v0d10v5 ad=8.12e+12p pd=6.006e+07u as=4.64e+12p ps=3.432e+07u w=4e+06u l=1e+06u
X36 a_8404_8048# a_8284_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X37 vss vss.t196 vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X38 a_n22428_2672# a_n22834_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X39 a_n24544_2674# a_n23894_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X40 bandgapmd_0.otam_1.pmosrm_0.out vss.t354 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X41 vdd.t91 ldomc_0.otaldom_0.pmosrm_0.out out.t59 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X42 bandgapmd_0.otam_1.nmosrm_0.outn.t32 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.pcsm_0.diff vdd.t281 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X43 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmoslm_0.outp vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.22e+12p pd=4.122e+07u as=4.64e+12p ps=3.896e+07u w=2e+06u l=4e+06u
X44 bandgapmd_0.otam_1.pmosrm_0.out vss.t353 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X45 vss vss.t198 bandgapmd_0.bg_trimmup_0.bot sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X46 bandgapmd_0.otam_1.nmosrm_0.outn.t31 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.pcsm_0.diff vdd.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X47 vdd.t173 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.diff vdd.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X48 bandgapmd_0.otam_1.pcascodeupm_0.o1.t7 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t33 vdd.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X49 a_n22428_2672# a_n21774_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X50 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o1.t15 vdd.t271 sky130_fd_pr__pfet_g5v0d10v5 ad=5.22e+12p pd=4.122e+07u as=0p ps=0u w=2e+06u l=4e+06u
X51 vss vss.t192 vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X52 vss.t309 vss.t310 vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X53 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t171 vdd.t170 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X54 bandgapmd_0.otam_1.pmosrm_0.out vss.t352 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X55 out.t67 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X56 a_8524_8048# a_9124_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X57 ldomc_0.otaldom_0.nmosrm_0.outn bandgapmd_0.bg_pmosm_0.vbg.t4 ldomc_0.otaldom_0.pcsm_0.diff vdd.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X58 ldomc_0.otaldom_0.pcascodeupm_0.o1.t15 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t388 vdd.t387 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X59 bandgapmd_0.otam_1.pmosrm_0.out vss.t351 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X60 vdd.t237 vdd.t235 vdd.t236 vdd.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X61 out.t58 ldomc_0.otaldom_0.pmosrm_0.out vdd.t90 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X62 bandgapmd_0.bg_stupm_0.vs2 vss.t221 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X63 bandgapmd_0.otam_1.pmosrm_0.out vss.t350 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X64 vss vss.t187 vss vss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X65 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.nmoslm_0.outp vdd.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+12p ps=4.29e+07u w=4e+06u l=1e+06u
X66 out.t57 ldomc_0.otaldom_0.pmosrm_0.out vdd.t89 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X67 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X68 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.nmosrm_0.outn.t30 vdd.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X69 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o1.t6 vdd.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X70 a_n11444_2076# bandgapmd_0.bg_pmosm_0.comp.t0 vss.t313 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X71 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmoslm_0.outp vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X72 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmosrm_0.outn.t23 vss sky130_fd_pr__nfet_g5v0d10v5 ad=5.51e+12p pd=4.38e+07u as=0p ps=0u w=2e+06u l=4e+06u
X73 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.nmosrm_0.outn.t29 vdd.t278 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X74 vss vss.t183 vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X75 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t169 vdd.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X76 bandgapmd_0.bg_stupm_0.vs2 vss.t220 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X77 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcsm_0.diff vdd.t334 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X78 vss vss.t174 bandgapmd_0.bg_trimmup_0.bot sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X79 a_n14486_2076# a_n13784_5108# vss.t318 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X80 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t31 vdd.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X81 vdd.t29 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o2 vdd.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X82 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o1.t14 vdd.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X83 ldomc_0.otaldom_0.pmosrm_0.out out.t21 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X84 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X85 ldomc_0.otaldom_0.pdiffm_0.inp a_8284_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X86 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o1.t5 vdd.t310 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X87 bandgapmd_0.bg_pmosm_0.vbg.t1 bandgapmd_0.otam_1.pmosrm_0.out vdd.t343 vdd.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X88 vss.t6 biasbgr.t4 bandgapmd_0.otam_1.pmosrm_0.bias1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+07u
X89 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmoslm_0.outp vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X90 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff vdd.t247 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X91 ldomc_0.otaldom_0.pmosrm_0.out out.t20 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X92 vdd.t137 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.vbn2 vdd.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u w=4e+06u l=1e+06u
X93 out.t56 ldomc_0.otaldom_0.pmosrm_0.out vdd vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X94 a_n13316_2076# a_n12848_5108# vss.t226 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X95 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X96 vdd.t234 vdd.t232 vdd.t233 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X97 vss.t300 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosrm_0.outn vss.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X98 out.t68 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X99 vss.t358 biasldo.t2 biasldo.t3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+07u
X100 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X101 a_n23460_2674# a_n23894_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X102 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t76 vss.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X103 out.t55 ldomc_0.otaldom_0.pmosrm_0.out vdd.t86 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X104 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o1.t4 vdd.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X105 ldomc_0.otaldom_0.pcascodeupm_0.o1.t14 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t386 vdd.t385 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X106 bandgapmd_0.otam_1.pmosrm_0.out vss.t349 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X107 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t135 vdd.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X108 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t133 vdd.t132 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X109 vdd.t231 vdd.t229 vdd.t230 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X110 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.out vdd.t269 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.22e+12p ps=4.122e+07u w=2e+06u l=4e+06u
X111 bandgapmd_0.bg_stupm_0.vs2 vss.t219 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X112 vdd vdd.t224 vdd vdd.t225 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X113 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t298 vss.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X114 a_n21356_2676# a_n21774_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X115 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 vdd.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X116 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcsm_0.vbn2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X117 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t296 vss.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X118 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t294 vss.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X119 vss.t74 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmoslm_0.outp vss.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X120 vss.t72 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmoslm_0.outp vss.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X121 vdd.t26 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o1.t6 vdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X122 vdd.t131 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.diff vdd.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X123 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X124 ldomc_0.otaldom_0.pcascodeupm_0.o2.t15 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t384 vdd.t383 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X125 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X126 vss.t70 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmoslm_0.outp vss.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X127 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X128 vdd.t129 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X129 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X130 a_8524_8048# a_8164_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X131 vss.t292 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmoslm_0.outp vss.t291 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X132 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcsm_0.vbn2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=4.64e+12p pd=3.722e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X133 bandgapmd_0.bg_stupm_0.vs2 vss.t218 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X134 a_n20290_2674# a_n19654_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X135 vss.t290 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmoslm_0.outp vss.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X136 bandgapmd_0.otam_1.nmosrm_0.outn.t14 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t68 vss.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X137 bandgapmd_0.otam_1.nmosrm_0.outn.t13 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t66 vss.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X138 vdd.t167 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.diff vdd.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X139 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X140 bandgapmd_0.otam_1.nmosrm_0.outn.t12 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t64 vss.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X141 vss vss.t178 vss vss.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X142 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t288 vss.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X143 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 vdd.t267 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X144 ldomc_0.otaldom_0.pcascodeupm_0.o2.t7 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.out vdd.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.22e+12p ps=4.122e+07u w=2e+06u l=4e+06u
X145 vss vss.t172 bandgapmd_0.bg_trimmup_0.bot sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X146 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t286 vss.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X147 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t284 vss.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X148 a_n18160_2676# a_n17534_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X149 vss vss.t176 bandgapmd_0.otam_1.pdiffm_0.inn sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X150 vss.t62 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosrm_0.outn.t11 vss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X151 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X152 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o2 vdd.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X153 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 vdd.t265 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X154 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t282 vss.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X155 a_n11444_2076# a_n11678_5108# vss.t11 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X156 bandgapmd_0.bg_trimmup_0.bot trim[0].t0 a_n24956_4148# vss.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=9.28e+12p pd=7.328e+07u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X157 vss.t60 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosrm_0.outn.t10 vss.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X158 ldomc_0.otaldom_0.pmosrm_0.out out.t19 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X159 a_8404_8048# a_9244_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X160 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t307 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X161 vdd.t21 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o2 vdd.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X162 bandgapmd_0.otam_1.pmosrm_0.out vss.t348 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X163 vss.t58 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X164 a_n14486_2076# a_n14720_5108# vss.t330 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X165 vss.t327 vss.t328 vss.t326 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X166 vdd.t101 bandgapmd_0.bg_stupm_0.vs2.t0 bandgapmd_0.bg_stupm_0.vs2 vdd.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=1e+06u
X167 vdd.t382 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o1.t13 vdd.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X168 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o1.t13 vdd.t264 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X169 bandgapmd_0.otam_1.nmosrm_0.outn.t22 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X170 a_n7846_4436# bandgapmd_0.bg_pmosm_0.vbg.t5 vss.t315 vss.t314 sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X171 ldomc_0.otaldom_0.nmosrm_0.outn bandgapmd_0.bg_pmosm_0.vbg.t6 ldomc_0.otaldom_0.pcsm_0.diff vdd.t285 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X172 bandgapmd_0.otam_1.pmosrm_0.out vss.t347 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X173 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pdiffm_0.inp.t3 bandgapmd_0.otam_1.pcsm_0.diff vdd.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X174 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X175 vdd.t342 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.bg_pmosm_0.comp.t2 vdd.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X176 ldomc_0.otaldom_0.pcascodeupm_0.o1.t3 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t306 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X177 a_n13550_2076# a_n13784_5108# vss.t212 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X178 vdd.t380 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o1.t12 vdd.t379 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X179 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t127 vdd.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X180 vdd vdd.t219 vdd vdd.t220 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X181 vss.t280 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X182 vss vss.t170 bandgapmd_0.bg_trimmup_0.bot sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X183 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff vdd.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X184 vdd.t165 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.diff vdd.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X185 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.nmoslm_0.outp vdd.t333 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X186 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 vdd.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X187 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X188 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o2 vdd.t263 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X189 bandgapmd_0.bg_pmosm_0.vbg.t7 vss.t316 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X190 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X191 vss.t5 biasbgr.t2 biasbgr.t3 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+07u
X192 bandgapmd_0.otam_1.pmosrm_0.out vss.t346 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X193 a_n24544_2674# trim[1].t0 bandgapmd_0.bg_trimmup_0.bot vss.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X194 vdd.t378 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o2.t14 vdd.t377 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X195 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcsm_0.diff vdd.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X196 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pdiffm_0.inp.t4 bandgapmd_0.otam_1.pcsm_0.diff vdd.t346 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X197 out.t69 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X198 bandgapmd_0.otam_1.pmosrm_0.out vss.t345 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X199 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcsm_0.diff vdd.t331 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X200 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X201 a_n19218_2674# a_n19654_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X202 vdd.t19 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o1.t5 vdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X203 a_n20290_2674# a_n20714_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X204 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff vdd.t245 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X205 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t278 vss.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X206 bandgapmd_0.otam_1.pmosrm_0.out vss.t344 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X207 out.t70 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X208 vdd.t376 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o1.t11 vdd.t375 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X209 ldomc_0.otaldom_0.pcsm_0.diff bandgapmd_0.bg_pmosm_0.vbg.t8 ldomc_0.otaldom_0.nmosrm_0.outn vdd.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X210 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff vdd.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X211 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff vdd.t244 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X212 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmosrm_0.outn vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X213 bandgapmd_0.bg_resm_0.trimup bandgapmd_0.otam_1.pdiffm_0.inp vss.t217 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X214 bandgapmd_0.bg_resm_0.trimup a_n17534_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X215 a_n19218_2674# a_n18594_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X216 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X217 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff vdd.t243 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X218 ldomc_0.otaldom_0.pdiffm_0.inp a_8644_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X219 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X220 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inp.t5 bandgapmd_0.otam_1.nmoslm_0.outp vdd.t347 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X221 a_n12146_2076# a_n12848_5108# vss.t321 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X222 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o2.t6 vdd.t304 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X223 vss.t230 vss.t231 vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X224 ldomc_0.otaldom_0.pmosrm_0.out out.t18 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X225 ldomc_0.otaldom_0.pcascodeupm_0.o2.t13 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t373 vdd.t372 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X226 vdd.t17 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o2 vdd.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X227 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t371 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X228 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff vdd.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X229 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t163 vdd.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X230 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t125 vdd.t124 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X231 vss vss.t168 bandgapmd_0.bg_trimmup_0.bot sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X232 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X233 a_n15188_2076# bandgapmd_0.otam_1.pdiffm_0.inp.t0 vss.t216 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X234 ldomc_0.otaldom_0.pmosrm_0.out out.t17 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X235 a_n11210_2076# a_n11912_5108# vss.t214 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X236 bandgapmd_0.otam_1.pmosrm_0.out vss.t343 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X237 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 vdd.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X238 vss.t276 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosrm_0.outn vss.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X239 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o2.t5 vdd.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X240 vdd.t218 vdd.t216 vdd.t217 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X241 bandgapmd_0.bg_trimmup_0.bot a_n24956_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X242 out.t1 a_9244_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X243 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcsm_0.vbn2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X244 vdd.t369 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o2.t12 vdd.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X245 vdd.t123 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.diff vdd.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X246 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.nmosrm_0.outn.t28 vdd.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X247 vdd vdd.t211 vdd vdd.t212 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X248 out.t71 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X249 vdd.t210 vdd.t208 vdd.t209 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X250 vss.t274 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosrm_0.outn vss.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X251 bandgapmd_0.otam_1.nmosrm_0.outn.t27 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.pcsm_0.diff vdd.t276 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X252 vdd.t207 vdd.t205 vdd.t206 vdd.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X253 vdd.t161 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X254 vss.t272 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosrm_0.outn vss.t271 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X255 ldomc_0.otaldom_0.pmosrm_0.out out.t16 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X256 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t56 vss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X257 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t15 vdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X258 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmoslm_0.outp vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X259 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o2 vdd.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X260 bandgapmd_0.otam_1.pmosrm_0.out vss.t342 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X261 bandgapmd_0.bg_stupm_0.vs2 vdd.t203 vss.t361 vdd.t204 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X262 vdd.t159 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.vbn2 vdd.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u w=4e+06u l=1e+06u
X263 vdd.t13 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o1.t4 vdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X264 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmoslm_0.outp vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X265 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X266 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t270 vss.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X267 a_n12146_2076# a_n11912_5108# vss.t8 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X268 vdd.t202 vdd.t199 vdd.t201 vdd.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X269 vss.t54 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmoslm_0.outp vss.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X270 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X271 ldomc_0.otaldom_0.pmosrm_0.bias1 biasldo.t4 vss.t322 vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+07u
X272 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out vdd.t341 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X273 vss vss.t166 bandgapmd_0.bg_trimmup_0.bot sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X274 a_n15188_2076# a_n14954_5108# vss.t3 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X275 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o1.t2 vdd.t302 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X276 a_n18160_2676# a_n18594_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X277 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmoslm_0.outp vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X278 ldomc_0.otaldom_0.pmosrm_0.out out.t15 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X279 bandgapmd_0.otam_1.nmosrm_0.outn.t9 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t52 vss.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X280 vss.t268 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmoslm_0.outp vss.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X281 vdd.t121 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.diff vdd.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X282 vss.t165 vss.t162 vss.t164 vss.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X283 ldomc_0.otaldom_0.pmosrm_0.out out.t14 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X284 ldomc_0.otaldom_0.pcascodeupm_0.o2.t11 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t367 vdd.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X285 bandgapmd_0.otam_1.nmosrm_0.outn.t8 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t50 vss.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X286 vss.t228 vss.t229 vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X287 vdd.t157 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.diff vdd.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X288 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.nmosrm_0.outn.t26 vdd.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X289 vss.t48 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X290 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X291 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t155 vdd.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X292 bandgapmd_0.otam_1.pmosrm_0.out vss.t341 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X293 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o2 vdd.t260 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X294 a_n19218_2674# trim[11].t0 bandgapmd_0.bg_trimmup_0.bot vss.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X295 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t266 vss.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X296 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X297 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t153 vdd.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X298 ldomc_0.otaldom_0.pcascodeupm_0.o1.t10 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t365 vdd.t364 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X299 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t46 vss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X300 vss.t44 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosrm_0.outn.t7 vss.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X301 vss.t42 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosrm_0.outn.t6 vss.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X302 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X303 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t119 vdd.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X304 vdd.t11 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o2 vdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X305 vss vss.t157 vss vss.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X306 vdd vdd.t194 vdd vdd.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X307 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcsm_0.vbn2 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X308 out.t72 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X309 vdd vdd.t189 vdd vdd.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X310 bandgapmd_0.bg_trimmup_0.bot trim[2].t0 a_n23894_4148# vss.t319 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X311 ldomc_0.otaldom_0.pcascodeupm_0.o2.t4 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.out vdd.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X312 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t40 vss.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X313 vdd.t117 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.diff vdd.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X314 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t151 vdd.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X315 vss vss.t152 vss vss.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X316 ldomc_0.otaldom_0.pcascodeupm_0.o1.t9 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t363 vdd.t362 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X317 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X318 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t38 vss.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X319 ldomc_0.otaldom_0.nmosrm_0.outn bandgapmd_0.bg_pmosm_0.vbg.t9 ldomc_0.otaldom_0.pcsm_0.diff vdd.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X320 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 vdd.t300 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X321 a_8764_8048# a_8644_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X322 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t149 vdd.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X323 vdd.t188 vdd.t185 vdd.t187 vdd.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X324 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.out vdd.t259 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X325 out.t73 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X326 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X327 ldomc_0.otaldom_0.pcascodeupm_0.o2.t3 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.out vdd.t299 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X328 vdd vdd.t180 vdd vdd.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X329 vss.t151 vss.t149 vss.t150 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X330 out.t74 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X331 bandgapmd_0.bg_trimmup_0.bot trim[4].t0 a_n22834_4148# vss.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X332 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X333 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.nmoslm_0.outp vdd.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X334 bandgapmd_0.otam_1.pmosrm_0.out vss.t340 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X335 vss vss.t147 bandgapmd_0.bg_trimmup_0.bot sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X336 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t9 vdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X337 bandgapmd_0.otam_1.pmosrm_0.out vss.t339 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X338 out.t0 a_9124_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X339 a_n13550_2076# a_n12614_5108# vss.t215 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X340 vdd ldomc_0.otaldom_0.pmosrm_0.out out.t54 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X341 vdd.t147 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.vbn2 vdd.t146 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X342 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X343 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out vdd.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X344 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X345 ldomc_0.otaldom_0.pcascodeupm_0.o1.t1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X346 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 vdd.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X347 vss vss.t143 vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X348 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X349 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out vdd.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X350 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pdiffm_0.inp.t6 bandgapmd_0.otam_1.pcsm_0.diff vdd.t348 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X351 vdd.t81 ldomc_0.otaldom_0.pmosrm_0.out out.t53 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X352 vdd.t179 vdd.t176 vdd.t178 vdd.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X353 vss.t1 vss.t2 vss.t0 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X354 vdd.t361 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o2.t10 vdd.t360 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X355 bandgapmd_0.otam_1.pmosrm_0.out vss.t338 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X356 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out vdd.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X357 ldomc_0.otaldom_0.pcsm_0.diff bandgapmd_0.bg_pmosm_0.vbg.t10 ldomc_0.otaldom_0.nmosrm_0.outn vdd.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X358 biasbgr.t1 biasbgr.t0 vss.t4 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+07u
X359 vss.t142 vss.t140 vss.t141 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X360 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X361 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X362 out.t52 ldomc_0.otaldom_0.pmosrm_0.out vdd.t79 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X363 ldomc_0.otaldom_0.pmosrm_0.out out.t13 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X364 a_n15422_2076# a_n14720_5108# vss.t12 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X365 ldomc_0.otaldom_0.pcascodeupm_0.o2.t2 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.out vdd.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X366 bandgapmd_0.bg_trimmup_0.bot trim[14].t0 a_n17534_4148# vss.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X367 vss.t305 vss.t306 vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X368 vss.t264 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmoslm_0.outp vss.t263 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X369 out.t75 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X370 ldomc_0.otaldom_0.pmosrm_0.out out.t12 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X371 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff vdd.t319 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X372 out.t51 ldomc_0.otaldom_0.pmosrm_0.out vdd.t78 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X373 bandgapmd_0.otam_1.pcascodeupm_0.o1.t3 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t7 vdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X374 out.t76 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X375 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t115 vdd.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X376 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t262 vss.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X377 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inp.t7 bandgapmd_0.otam_1.nmoslm_0.outp vdd.t349 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X378 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X379 out.t77 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X380 a_n22428_2672# trim[5].t0 bandgapmd_0.bg_trimmup_0.bot vss.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X381 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X382 bandgapmd_0.otam_1.nmosrm_0.outn.t21 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X383 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X384 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff vdd.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X385 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X386 ldomc_0.otaldom_0.pmosrm_0.out out.t11 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X387 bandgapmd_0.bg_trimmup_0.bot trim[10].t0 a_n19654_4148# vss.t355 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X388 bandgapmd_0.otam_1.pmosrm_0.out vss.t337 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X389 vdd.t113 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X390 ldomc_0.otaldom_0.pcsm_0.diff bandgapmd_0.bg_pmosm_0.vbg.t11 ldomc_0.otaldom_0.nmosrm_0.outn vdd.t289 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X391 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X392 bandgapmd_0.bg_pmosm_0.comp.t1 bandgapmd_0.otam_1.pmosrm_0.out vdd.t340 vdd.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X393 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out vdd.t339 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X394 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X395 vss.t260 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosrm_0.outn vss.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X396 vdd.t77 ldomc_0.otaldom_0.pmosrm_0.out out.t50 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X397 a_n14252_2076# a_n14954_5108# vss.t307 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X398 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inp.t8 bandgapmd_0.otam_1.nmoslm_0.outp vdd.t350 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X399 a_n20290_2674# trim[9].t0 bandgapmd_0.bg_trimmup_0.bot vss.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X400 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t111 vdd.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X401 out.t49 ldomc_0.otaldom_0.pmosrm_0.out vdd.t76 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X402 a_8764_8048# a_8884_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X403 vdd.t75 ldomc_0.otaldom_0.pmosrm_0.out out.t48 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X404 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t258 vss.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X405 vss vss.t135 vss vss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X406 a_n13316_2076# a_n14018_5108# vss.t227 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X407 out.t47 ldomc_0.otaldom_0.pmosrm_0.out vdd.t74 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X408 vdd.t145 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X409 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t256 vss.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X410 vss.t36 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmoslm_0.outp vss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X411 ldomc_0.otaldom_0.pmosrm_0.out out.t10 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X412 vdd.t109 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.vbn2 vdd.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X413 vss.t34 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmoslm_0.outp vss.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X414 vss vss.t130 vss vss.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X415 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff vdd.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X416 vss.t32 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmoslm_0.outp vss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X417 vss.t30 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmoslm_0.outp vss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X418 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t28 vss.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X419 vss.t254 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmoslm_0.outp vss.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X420 a_n11210_2076# bandgapmd_0.bg_pmosm_0.vbg.t2 vss.t356 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X421 vdd ldomc_0.otaldom_0.pmosrm_0.out out.t46 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X422 bandgapmd_0.otam_1.nmosrm_0.outn.t25 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.pcsm_0.diff vdd.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X423 out.t78 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X424 ldomc_0.otaldom_0.pmosrm_0.out out.t9 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X425 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmosrm_0.outn vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X426 vss.t252 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmoslm_0.outp vss.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X427 vss.t250 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmoslm_0.outp vss.t249 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X428 bandgapmd_0.otam_1.pmosrm_0.out vss.t336 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X429 bandgapmd_0.otam_1.nmosrm_0.outn.t5 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t26 vss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X430 bandgapmd_0.otam_1.pcascodeupm_0.o1.t12 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X431 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o2.t1 vdd.t295 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X432 out.t45 ldomc_0.otaldom_0.pmosrm_0.out vdd vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X433 bandgapmd_0.otam_1.nmosrm_0.outn.t4 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t24 vss.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X434 vdd.t69 ldomc_0.otaldom_0.pmosrm_0.out out.t44 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X435 bandgapmd_0.otam_1.pcascodeupm_0.o1.t11 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X436 ldomc_0.otaldom_0.pmosrm_0.out out.t8 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X437 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t143 vdd.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X438 out.t43 ldomc_0.otaldom_0.pmosrm_0.out vdd.t67 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X439 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t248 vss.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X440 out.t42 ldomc_0.otaldom_0.pmosrm_0.out vdd vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X441 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t246 vss.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X442 vss.t22 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosrm_0.outn.t3 vss.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X443 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 vdd.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X444 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o2.t0 vdd.t294 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X445 vss.t20 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosrm_0.outn.t2 vss.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X446 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmoslm_0.outp vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X447 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmosrm_0.outn.t20 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X448 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 vdd.t255 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X449 out.t41 ldomc_0.otaldom_0.pmosrm_0.out vdd.t65 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X450 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 vdd.t293 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X451 ldomc_0.otaldom_0.pmosrm_0.out out.t7 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X452 vss vss.t125 vss vss.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X453 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.nmosrm_0.outn.t24 vdd.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X454 bandgapmd_0.otam_1.pmosrm_0.out a_n7846_4436# vss.t10 vss.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X455 ldomc_0.otaldom_0.nmosrm_0.outn bandgapmd_0.bg_pmosm_0.vbg.t12 ldomc_0.otaldom_0.pcsm_0.diff vdd.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X456 bandgapmd_0.otam_1.pmosrm_0.bias1 biasbgr.t5 vss.t7 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+07u
X457 vdd.t64 ldomc_0.otaldom_0.pmosrm_0.out out.t40 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X458 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmoslm_0.outp vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X459 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmosrm_0.outn.t19 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X460 bandgapmd_0.otam_1.pcascodeupm_0.o1.t10 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X461 out.t79 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X462 out.t39 ldomc_0.otaldom_0.pmosrm_0.out vdd vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X463 bandgapmd_0.otam_1.pmosrm_0.out vss.t335 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X464 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t107 vdd.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X465 bandgapmd_0.bg_resm_0.trimup trim[15].t0 bandgapmd_0.bg_trimmup_0.bot vss.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X466 vdd.t61 ldomc_0.otaldom_0.pmosrm_0.out out.t38 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X467 vdd.t141 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.diff vdd.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X468 a_n18160_2676# trim[13].t0 bandgapmd_0.bg_trimmup_0.bot vss.t317 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X469 bandgapmd_0.bg_trimmup_0.bot trim[6].t0 a_n21774_4148# vss.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X470 vdd ldomc_0.otaldom_0.pmosrm_0.out out.t37 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X471 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcsm_0.vbp1 vdd.t253 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X472 out.t80 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X473 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.nmoslm_0.outp vdd.t329 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X474 out.t36 ldomc_0.otaldom_0.pmosrm_0.out vdd.t58 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X475 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.nmoslm_0.outp vdd.t328 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X476 vdd.t57 ldomc_0.otaldom_0.pmosrm_0.out out.t35 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X477 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.out vdd.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X478 a_n23460_2674# trim[3].t0 bandgapmd_0.bg_trimmup_0.bot vss.t324 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X479 bandgapmd_0.otam_1.pmosrm_0.out vss.t334 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X480 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pmosrm_0.bias1 vdd.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X481 vdd.t338 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.bg_pmosm_0.vbg.t0 vdd.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X482 a_n14252_2076# a_n14018_5108# vss.t312 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X483 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcsm_0.diff vdd.t327 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X484 vss vss.t121 vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X485 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcsm_0.diff vdd.t326 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X486 out.t34 ldomc_0.otaldom_0.pmosrm_0.out vdd.t55 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X487 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out vdd.t337 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X488 ldomc_0.otaldom_0.pmosrm_0.out out.t6 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X489 vdd ldomc_0.otaldom_0.pmosrm_0.out out.t33 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X490 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o1.t9 vdd.t252 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X491 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t359 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X492 a_n12380_2076# a_n11678_5108# vss.t211 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X493 out.t32 ldomc_0.otaldom_0.pmosrm_0.out vdd.t52 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X494 out.t81 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X495 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmosrm_0.outn.t18 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X496 ldomc_0.otaldom_0.pcsm_0.diff bandgapmd_0.bg_pmosm_0.vbg.t13 ldomc_0.otaldom_0.nmosrm_0.outn vdd.t315 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X497 bandgapmd_0.bg_trimmup_0.bot trim[8].t0 a_n20714_4148# vss.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X498 bandgapmd_0.otam_1.pmosrm_0.out vss.t333 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X499 vdd.t51 ldomc_0.otaldom_0.pmosrm_0.out out.t31 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X500 vdd ldomc_0.otaldom_0.pmosrm_0.out out.t30 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X501 bandgapmd_0.otam_1.pcascodeupm_0.o1.t2 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t5 vdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X502 out.t82 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X503 vdd.t48 ldomc_0.otaldom_0.pmosrm_0.out out.t29 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X504 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.diff vdd.t241 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X505 out.t83 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X506 bandgapmd_0.otam_1.pmosrm_0.out vss.t332 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X507 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.out vdd.t251 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X508 vss vss.t116 vss vss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X509 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X510 out.t84 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X511 biasldo.t1 biasldo.t0 vss.t357 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+07u
X512 out.t28 ldomc_0.otaldom_0.pmosrm_0.out vdd vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X513 ldomc_0.otaldom_0.pcascodeupm_0.o2.t9 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t358 vdd.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X514 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.vbp1 vdd.t105 vdd.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X515 vdd.t45 ldomc_0.otaldom_0.pmosrm_0.out out.t27 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X516 vss vss.t112 vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X517 out.t26 ldomc_0.otaldom_0.pmosrm_0.out vdd.t44 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X518 vss.t244 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosrm_0.outn vss.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X519 out.t25 ldomc_0.otaldom_0.pmosrm_0.out vdd vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X520 ldomc_0.otaldom_0.pcsm_0.diff bandgapmd_0.bg_pmosm_0.vbg.t14 ldomc_0.otaldom_0.nmosrm_0.outn vdd.t316 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X521 vdd.t41 ldomc_0.otaldom_0.pmosrm_0.out out.t24 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X522 bandgapmd_0.otam_1.pcascodeupm_0.o1.t8 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t250 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X523 vdd.t103 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.diff vdd.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X524 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X525 vss vss.t110 bandgapmd_0.bg_trimmup_0.bot sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1
X526 out.t23 ldomc_0.otaldom_0.pmosrm_0.out vdd.t40 vdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X527 vss.t242 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosrm_0.outn vss.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X528 vss vss.t105 vss vss.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X529 vss vss.t100 vss vss.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X530 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X531 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out vdd.t336 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X532 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t18 vss.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X533 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pdiffm_0.inp.t9 bandgapmd_0.otam_1.pcsm_0.diff vdd.t351 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X534 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.diff vdd.t317 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X535 vss.t359 a_8884_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X536 bandgapmd_0.otam_1.nmosrm_0.outn.t17 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X537 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X538 ldomc_0.otaldom_0.pmosrm_0.out out.t5 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X539 a_n21356_2676# trim[7].t0 bandgapmd_0.bg_trimmup_0.bot vss.t329 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X540 bandgapmd_0.otam_1.pmosrm_0.out vss.t331 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X541 vss.t99 vss.t96 vss.t98 vss.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X542 ldomc_0.otaldom_0.pcascodeupm_0.o1.t0 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.vg vdd.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X543 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.out vdd.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X544 ldomc_0.otaldom_0.pmosrm_0.out out.t4 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X545 a_n23460_2674# a_n22834_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X546 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X547 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X548 vss vss.t91 vss vss.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X549 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t240 vss.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X550 ldomc_0.otaldom_0.pmosrm_0.out out.t3 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X551 vdd.t356 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o1.t8 vdd.t355 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X552 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.vg vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X553 out.t85 ldomc_0.otaldom_0.pdiffm_0.inp sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X554 vss.t238 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmoslm_0.outp vss.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X555 a_n12380_2076# a_n12614_5108# vss.t232 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
X556 a_n21356_2676# a_n20714_4148# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X557 bandgapmd_0.otam_1.pcascodeupm_0.o1.t1 bandgapmd_0.otam_1.pcascodeupm_0.vg vdd.t3 vdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X558 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pdiffm_0.inp.t10 bandgapmd_0.otam_1.pcsm_0.diff vdd.t352 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X559 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t236 vss.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X560 bandgapmd_0.otam_1.nmosrm_0.outn.t1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss.t16 vss.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X561 vss.t90 vss.t87 vss.t89 vss.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X562 bandgapmd_0.bg_trimmup_0.bot trim[12].t0 a_n18594_4148# vss.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X563 vdd.t1 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o1.t0 vdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X564 vdd.t354 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o2.t8 vdd.t353 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X565 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inp.t11 bandgapmd_0.otam_1.nmoslm_0.outp vdd.t325 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X566 bandgapmd_0.otam_1.nmosrm_0.outn.t16 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pmosrm_0.out vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X567 ldomc_0.otaldom_0.pdiffm_0.inp a_8164_10248# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X568 vss.t323 biasldo.t5 ldomc_0.otaldom_0.pmosrm_0.bias1 vss sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+07u
X569 vdd ldomc_0.otaldom_0.pmosrm_0.out out.t22 vdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+07u l=500000u
X570 vss.t14 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.otam_1.nmosrm_0.outn.t0 vss.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X571 ldomc_0.otaldom_0.pmosrm_0.out out.t2 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X572 vss.t234 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X573 a_n15422_2076# bandgapmd_0.otam_1.pdiffm_0.inn vss.t325 sky130_fd_pr__res_xhigh_po_0p69 l=1.3e+07u
R0 vss.n2 vss.n17626 10.418
R1 vss.n20295 vss.n0 10.418
R2 vss.n6 vss.n4236 10.418
R3 vss.n6905 vss.n4 10.418
R4 vss.n20408 vss.n17547 13786.1
R5 vss.n7018 vss.n4157 13786.1
R6 vss.n20411 vss.n20410 7649.77
R7 vss.n7021 vss.n7020 7649.77
R8 vss.n20410 vss.n20409 6102.55
R9 vss.n7020 vss.n7019 6102.55
R10 vss.n20409 vss.n17548 2614.68
R11 vss.n7019 vss.n4158 2614.68
R12 vss.n20294 vss.n17619 1534.21
R13 vss.n20283 vss.n20282 1534.21
R14 vss.n20282 vss.n19036 1534.21
R15 vss.n20275 vss.n20274 1534.21
R16 vss.n20268 vss.n20267 1534.21
R17 vss.n20256 vss.n19050 1534.21
R18 vss.n20254 vss.n19060 1534.21
R19 vss.n20245 vss.n20244 1534.21
R20 vss.n20233 vss.n19070 1534.21
R21 vss.n20231 vss.n19079 1534.21
R22 vss.n20211 vss.n19101 1534.21
R23 vss.n20209 vss.n19102 1534.21
R24 vss.n20198 vss.n20197 1534.21
R25 vss.n20188 vss.n19120 1534.21
R26 vss.n20186 vss.n19121 1534.21
R27 vss.n20175 vss.n20174 1534.21
R28 vss.n20165 vss.n19139 1534.21
R29 vss.n20163 vss.n19140 1534.21
R30 vss.n20157 vss.n19140 1534.21
R31 vss.n20155 vss.n19145 1534.21
R32 vss.n20144 vss.n20143 1534.21
R33 vss.n20137 vss.n20136 1534.21
R34 vss.n20125 vss.n19160 1534.21
R35 vss.n20123 vss.n19170 1534.21
R36 vss.n20114 vss.n20113 1534.21
R37 vss.n20102 vss.n19180 1534.21
R38 vss.n20089 vss.n19196 1534.21
R39 vss.n20077 vss.n19208 1534.21
R40 vss.n20075 vss.n19209 1534.21
R41 vss.n20064 vss.n20063 1534.21
R42 vss.n20054 vss.n19227 1534.21
R43 vss.n20052 vss.n19228 1534.21
R44 vss.n20041 vss.n20040 1534.21
R45 vss.n20033 vss.n19245 1534.21
R46 vss.n20033 vss.n20032 1534.21
R47 vss.n19256 vss.n19246 1534.21
R48 vss.n20021 vss.n20020 1534.21
R49 vss.n20009 vss.n19258 1534.21
R50 vss.n20007 vss.n19267 1534.21
R51 vss.n19998 vss.n19997 1534.21
R52 vss.n19986 vss.n19277 1534.21
R53 vss.n19984 vss.n19286 1534.21
R54 vss.n19964 vss.n19308 1534.21
R55 vss.n19962 vss.n19309 1534.21
R56 vss.n19951 vss.n19950 1534.21
R57 vss.n19941 vss.n19327 1534.21
R58 vss.n19939 vss.n19328 1534.21
R59 vss.n19928 vss.n19927 1534.21
R60 vss.n19918 vss.n19346 1534.21
R61 vss.n19916 vss.n19347 1534.21
R62 vss.n19910 vss.n19347 1534.21
R63 vss.n19908 vss.n19352 1534.21
R64 vss.n19897 vss.n19896 1534.21
R65 vss.n19890 vss.n19889 1534.21
R66 vss.n19878 vss.n19367 1534.21
R67 vss.n19876 vss.n19377 1534.21
R68 vss.n19867 vss.n19866 1534.21
R69 vss.n19855 vss.n19387 1534.21
R70 vss.n19842 vss.n19403 1534.21
R71 vss.n19830 vss.n19415 1534.21
R72 vss.n19828 vss.n19416 1534.21
R73 vss.n19817 vss.n19816 1534.21
R74 vss.n19807 vss.n19434 1534.21
R75 vss.n19805 vss.n19435 1534.21
R76 vss.n19794 vss.n19793 1534.21
R77 vss.n19786 vss.n19452 1534.21
R78 vss.n19786 vss.n19785 1534.21
R79 vss.n19463 vss.n19453 1534.21
R80 vss.n19774 vss.n19773 1534.21
R81 vss.n19762 vss.n19465 1534.21
R82 vss.n19760 vss.n19474 1534.21
R83 vss.n19751 vss.n19750 1534.21
R84 vss.n19739 vss.n19484 1534.21
R85 vss.n19737 vss.n19493 1534.21
R86 vss.n19717 vss.n19515 1534.21
R87 vss.n19715 vss.n19516 1534.21
R88 vss.n19704 vss.n19703 1534.21
R89 vss.n19694 vss.n19534 1534.21
R90 vss.n19692 vss.n19535 1534.21
R91 vss.n19681 vss.n19680 1534.21
R92 vss.n19671 vss.n19553 1534.21
R93 vss.n19669 vss.n19554 1534.21
R94 vss.n19663 vss.n19554 1534.21
R95 vss.n19661 vss.n19559 1534.21
R96 vss.n19650 vss.n19649 1534.21
R97 vss.n19643 vss.n19642 1534.21
R98 vss.n19631 vss.n19574 1534.21
R99 vss.n19629 vss.n19584 1534.21
R100 vss.n19601 vss.n19596 1534.21
R101 vss.n19609 vss.n19608 1534.21
R102 vss.n20349 vss.n20348 1534.21
R103 vss.n20342 vss.n17597 1534.21
R104 vss.n20340 vss.n17599 1534.21
R105 vss.n20334 vss.n17601 1534.21
R106 vss.n20328 vss.n20327 1534.21
R107 vss.n20323 vss.n20322 1534.21
R108 vss.n17613 vss.n17606 1534.21
R109 vss.n20312 vss.n20311 1534.21
R110 vss.n20311 vss.n20310 1534.21
R111 vss.n20300 vss.n20299 1534.21
R112 vss.n19019 vss.n17627 1534.21
R113 vss.n19017 vss.n17634 1534.21
R114 vss.n19011 vss.n17634 1534.21
R115 vss.n19009 vss.n17638 1534.21
R116 vss.n18998 vss.n18997 1534.21
R117 vss.n18991 vss.n18990 1534.21
R118 vss.n18979 vss.n17653 1534.21
R119 vss.n18977 vss.n17663 1534.21
R120 vss.n18968 vss.n18967 1534.21
R121 vss.n18956 vss.n17673 1534.21
R122 vss.n18943 vss.n17689 1534.21
R123 vss.n18931 vss.n17701 1534.21
R124 vss.n18929 vss.n17702 1534.21
R125 vss.n18918 vss.n18917 1534.21
R126 vss.n18908 vss.n17720 1534.21
R127 vss.n18906 vss.n17721 1534.21
R128 vss.n18895 vss.n18894 1534.21
R129 vss.n18887 vss.n17738 1534.21
R130 vss.n18887 vss.n18886 1534.21
R131 vss.n17749 vss.n17739 1534.21
R132 vss.n18875 vss.n18874 1534.21
R133 vss.n18863 vss.n17751 1534.21
R134 vss.n18861 vss.n17760 1534.21
R135 vss.n18852 vss.n18851 1534.21
R136 vss.n18840 vss.n17770 1534.21
R137 vss.n18838 vss.n17779 1534.21
R138 vss.n18818 vss.n17801 1534.21
R139 vss.n18816 vss.n17802 1534.21
R140 vss.n18805 vss.n18804 1534.21
R141 vss.n18795 vss.n17820 1534.21
R142 vss.n18793 vss.n17821 1534.21
R143 vss.n18782 vss.n18781 1534.21
R144 vss.n18772 vss.n17839 1534.21
R145 vss.n18770 vss.n17840 1534.21
R146 vss.n17849 vss.n17840 1534.21
R147 vss.n18762 vss.n18761 1534.21
R148 vss.n18750 vss.n17851 1534.21
R149 vss.n18748 vss.n17860 1534.21
R150 vss.n18739 vss.n18738 1534.21
R151 vss.n18727 vss.n17870 1534.21
R152 vss.n18725 vss.n17879 1534.21
R153 vss.n18716 vss.n18715 1534.21
R154 vss.n18702 vss.n17902 1534.21
R155 vss.n18688 vss.n17915 1534.21
R156 vss.n18677 vss.n18676 1534.21
R157 vss.n18667 vss.n17933 1534.21
R158 vss.n18665 vss.n17934 1534.21
R159 vss.n18654 vss.n18653 1534.21
R160 vss.n18646 vss.n17951 1534.21
R161 vss.n18646 vss.n18645 1534.21
R162 vss.n17962 vss.n17952 1534.21
R163 vss.n18634 vss.n18633 1534.21
R164 vss.n18622 vss.n17964 1534.21
R165 vss.n18620 vss.n17973 1534.21
R166 vss.n18611 vss.n18610 1534.21
R167 vss.n18599 vss.n17983 1534.21
R168 vss.n18597 vss.n17992 1534.21
R169 vss.n18577 vss.n18014 1534.21
R170 vss.n18575 vss.n18015 1534.21
R171 vss.n18564 vss.n18563 1534.21
R172 vss.n18554 vss.n18033 1534.21
R173 vss.n18552 vss.n18034 1534.21
R174 vss.n18541 vss.n18540 1534.21
R175 vss.n18531 vss.n18052 1534.21
R176 vss.n18529 vss.n18053 1534.21
R177 vss.n18062 vss.n18053 1534.21
R178 vss.n18521 vss.n18520 1534.21
R179 vss.n18509 vss.n18064 1534.21
R180 vss.n18507 vss.n18073 1534.21
R181 vss.n18498 vss.n18497 1534.21
R182 vss.n18486 vss.n18083 1534.21
R183 vss.n18484 vss.n18092 1534.21
R184 vss.n18475 vss.n18474 1534.21
R185 vss.n18461 vss.n18115 1534.21
R186 vss.n18449 vss.n18127 1534.21
R187 vss.n18447 vss.n18128 1534.21
R188 vss.n18436 vss.n18435 1534.21
R189 vss.n18426 vss.n18146 1534.21
R190 vss.n18424 vss.n18147 1534.21
R191 vss.n18413 vss.n18412 1534.21
R192 vss.n18405 vss.n18164 1534.21
R193 vss.n18405 vss.n18404 1534.21
R194 vss.n18175 vss.n18165 1534.21
R195 vss.n18393 vss.n18392 1534.21
R196 vss.n18381 vss.n18177 1534.21
R197 vss.n18379 vss.n18186 1534.21
R198 vss.n18370 vss.n18369 1534.21
R199 vss.n18358 vss.n18196 1534.21
R200 vss.n18356 vss.n18205 1534.21
R201 vss.n18336 vss.n18227 1534.21
R202 vss.n18334 vss.n18228 1534.21
R203 vss.n18323 vss.n18322 1534.21
R204 vss.n18313 vss.n18246 1534.21
R205 vss.n18311 vss.n18247 1534.21
R206 vss.n18300 vss.n18299 1534.21
R207 vss.n18290 vss.n18265 1534.21
R208 vss.n18288 vss.n18266 1534.21
R209 vss.n18277 vss.n18266 1534.21
R210 vss.n18280 vss.n18279 1534.21
R211 vss.n6904 vss.n4229 1534.21
R212 vss.n6893 vss.n6892 1534.21
R213 vss.n6892 vss.n5646 1534.21
R214 vss.n6885 vss.n6884 1534.21
R215 vss.n6878 vss.n6877 1534.21
R216 vss.n6866 vss.n5660 1534.21
R217 vss.n6864 vss.n5670 1534.21
R218 vss.n6855 vss.n6854 1534.21
R219 vss.n6843 vss.n5680 1534.21
R220 vss.n6841 vss.n5689 1534.21
R221 vss.n6821 vss.n5711 1534.21
R222 vss.n6819 vss.n5712 1534.21
R223 vss.n6808 vss.n6807 1534.21
R224 vss.n6798 vss.n5730 1534.21
R225 vss.n6796 vss.n5731 1534.21
R226 vss.n6785 vss.n6784 1534.21
R227 vss.n6775 vss.n5749 1534.21
R228 vss.n6773 vss.n5750 1534.21
R229 vss.n6767 vss.n5750 1534.21
R230 vss.n6765 vss.n5755 1534.21
R231 vss.n6754 vss.n6753 1534.21
R232 vss.n6747 vss.n6746 1534.21
R233 vss.n6735 vss.n5770 1534.21
R234 vss.n6733 vss.n5780 1534.21
R235 vss.n6724 vss.n6723 1534.21
R236 vss.n6712 vss.n5790 1534.21
R237 vss.n6699 vss.n5806 1534.21
R238 vss.n6687 vss.n5818 1534.21
R239 vss.n6685 vss.n5819 1534.21
R240 vss.n6674 vss.n6673 1534.21
R241 vss.n6664 vss.n5837 1534.21
R242 vss.n6662 vss.n5838 1534.21
R243 vss.n6651 vss.n6650 1534.21
R244 vss.n6643 vss.n5855 1534.21
R245 vss.n6643 vss.n6642 1534.21
R246 vss.n5866 vss.n5856 1534.21
R247 vss.n6631 vss.n6630 1534.21
R248 vss.n6619 vss.n5868 1534.21
R249 vss.n6617 vss.n5877 1534.21
R250 vss.n6608 vss.n6607 1534.21
R251 vss.n6596 vss.n5887 1534.21
R252 vss.n6594 vss.n5896 1534.21
R253 vss.n6574 vss.n5918 1534.21
R254 vss.n6572 vss.n5919 1534.21
R255 vss.n6561 vss.n6560 1534.21
R256 vss.n6551 vss.n5937 1534.21
R257 vss.n6549 vss.n5938 1534.21
R258 vss.n6538 vss.n6537 1534.21
R259 vss.n6528 vss.n5956 1534.21
R260 vss.n6526 vss.n5957 1534.21
R261 vss.n6520 vss.n5957 1534.21
R262 vss.n6518 vss.n5962 1534.21
R263 vss.n6507 vss.n6506 1534.21
R264 vss.n6500 vss.n6499 1534.21
R265 vss.n6488 vss.n5977 1534.21
R266 vss.n6486 vss.n5987 1534.21
R267 vss.n6477 vss.n6476 1534.21
R268 vss.n6465 vss.n5997 1534.21
R269 vss.n6452 vss.n6013 1534.21
R270 vss.n6440 vss.n6025 1534.21
R271 vss.n6438 vss.n6026 1534.21
R272 vss.n6427 vss.n6426 1534.21
R273 vss.n6417 vss.n6044 1534.21
R274 vss.n6415 vss.n6045 1534.21
R275 vss.n6404 vss.n6403 1534.21
R276 vss.n6396 vss.n6062 1534.21
R277 vss.n6396 vss.n6395 1534.21
R278 vss.n6073 vss.n6063 1534.21
R279 vss.n6384 vss.n6383 1534.21
R280 vss.n6372 vss.n6075 1534.21
R281 vss.n6370 vss.n6084 1534.21
R282 vss.n6361 vss.n6360 1534.21
R283 vss.n6349 vss.n6094 1534.21
R284 vss.n6347 vss.n6103 1534.21
R285 vss.n6327 vss.n6125 1534.21
R286 vss.n6325 vss.n6126 1534.21
R287 vss.n6314 vss.n6313 1534.21
R288 vss.n6304 vss.n6144 1534.21
R289 vss.n6302 vss.n6145 1534.21
R290 vss.n6291 vss.n6290 1534.21
R291 vss.n6281 vss.n6163 1534.21
R292 vss.n6279 vss.n6164 1534.21
R293 vss.n6273 vss.n6164 1534.21
R294 vss.n6271 vss.n6169 1534.21
R295 vss.n6260 vss.n6259 1534.21
R296 vss.n6253 vss.n6252 1534.21
R297 vss.n6241 vss.n6184 1534.21
R298 vss.n6239 vss.n6194 1534.21
R299 vss.n6211 vss.n6206 1534.21
R300 vss.n6219 vss.n6218 1534.21
R301 vss.n6959 vss.n6958 1534.21
R302 vss.n6952 vss.n4207 1534.21
R303 vss.n6950 vss.n4209 1534.21
R304 vss.n6944 vss.n4211 1534.21
R305 vss.n6938 vss.n6937 1534.21
R306 vss.n6933 vss.n6932 1534.21
R307 vss.n4223 vss.n4216 1534.21
R308 vss.n6922 vss.n6921 1534.21
R309 vss.n6921 vss.n6920 1534.21
R310 vss.n6910 vss.n6909 1534.21
R311 vss.n5629 vss.n4237 1534.21
R312 vss.n5627 vss.n4244 1534.21
R313 vss.n5621 vss.n4244 1534.21
R314 vss.n5619 vss.n4248 1534.21
R315 vss.n5608 vss.n5607 1534.21
R316 vss.n5601 vss.n5600 1534.21
R317 vss.n5589 vss.n4263 1534.21
R318 vss.n5587 vss.n4273 1534.21
R319 vss.n5578 vss.n5577 1534.21
R320 vss.n5566 vss.n4283 1534.21
R321 vss.n5553 vss.n4299 1534.21
R322 vss.n5541 vss.n4311 1534.21
R323 vss.n5539 vss.n4312 1534.21
R324 vss.n5528 vss.n5527 1534.21
R325 vss.n5518 vss.n4330 1534.21
R326 vss.n5516 vss.n4331 1534.21
R327 vss.n5505 vss.n5504 1534.21
R328 vss.n5497 vss.n4348 1534.21
R329 vss.n5497 vss.n5496 1534.21
R330 vss.n4359 vss.n4349 1534.21
R331 vss.n5485 vss.n5484 1534.21
R332 vss.n5473 vss.n4361 1534.21
R333 vss.n5471 vss.n4370 1534.21
R334 vss.n5462 vss.n5461 1534.21
R335 vss.n5450 vss.n4380 1534.21
R336 vss.n5448 vss.n4389 1534.21
R337 vss.n5428 vss.n4411 1534.21
R338 vss.n5426 vss.n4412 1534.21
R339 vss.n5415 vss.n5414 1534.21
R340 vss.n5405 vss.n4430 1534.21
R341 vss.n5403 vss.n4431 1534.21
R342 vss.n5392 vss.n5391 1534.21
R343 vss.n5382 vss.n4449 1534.21
R344 vss.n5380 vss.n4450 1534.21
R345 vss.n4459 vss.n4450 1534.21
R346 vss.n5372 vss.n5371 1534.21
R347 vss.n5360 vss.n4461 1534.21
R348 vss.n5358 vss.n4470 1534.21
R349 vss.n5349 vss.n5348 1534.21
R350 vss.n5337 vss.n4480 1534.21
R351 vss.n5335 vss.n4489 1534.21
R352 vss.n5326 vss.n5325 1534.21
R353 vss.n5312 vss.n4512 1534.21
R354 vss.n5298 vss.n4525 1534.21
R355 vss.n5287 vss.n5286 1534.21
R356 vss.n5277 vss.n4543 1534.21
R357 vss.n5275 vss.n4544 1534.21
R358 vss.n5264 vss.n5263 1534.21
R359 vss.n5256 vss.n4561 1534.21
R360 vss.n5256 vss.n5255 1534.21
R361 vss.n4572 vss.n4562 1534.21
R362 vss.n5244 vss.n5243 1534.21
R363 vss.n5232 vss.n4574 1534.21
R364 vss.n5230 vss.n4583 1534.21
R365 vss.n5221 vss.n5220 1534.21
R366 vss.n5209 vss.n4593 1534.21
R367 vss.n5207 vss.n4602 1534.21
R368 vss.n5187 vss.n4624 1534.21
R369 vss.n5185 vss.n4625 1534.21
R370 vss.n5174 vss.n5173 1534.21
R371 vss.n5164 vss.n4643 1534.21
R372 vss.n5162 vss.n4644 1534.21
R373 vss.n5151 vss.n5150 1534.21
R374 vss.n5141 vss.n4662 1534.21
R375 vss.n5139 vss.n4663 1534.21
R376 vss.n4672 vss.n4663 1534.21
R377 vss.n5131 vss.n5130 1534.21
R378 vss.n5119 vss.n4674 1534.21
R379 vss.n5117 vss.n4683 1534.21
R380 vss.n5108 vss.n5107 1534.21
R381 vss.n5096 vss.n4693 1534.21
R382 vss.n5094 vss.n4702 1534.21
R383 vss.n5085 vss.n5084 1534.21
R384 vss.n5071 vss.n4725 1534.21
R385 vss.n5059 vss.n4737 1534.21
R386 vss.n5057 vss.n4738 1534.21
R387 vss.n5046 vss.n5045 1534.21
R388 vss.n5036 vss.n4756 1534.21
R389 vss.n5034 vss.n4757 1534.21
R390 vss.n5023 vss.n5022 1534.21
R391 vss.n5015 vss.n4774 1534.21
R392 vss.n5015 vss.n5014 1534.21
R393 vss.n4785 vss.n4775 1534.21
R394 vss.n5003 vss.n5002 1534.21
R395 vss.n4991 vss.n4787 1534.21
R396 vss.n4989 vss.n4796 1534.21
R397 vss.n4980 vss.n4979 1534.21
R398 vss.n4968 vss.n4806 1534.21
R399 vss.n4966 vss.n4815 1534.21
R400 vss.n4946 vss.n4837 1534.21
R401 vss.n4944 vss.n4838 1534.21
R402 vss.n4933 vss.n4932 1534.21
R403 vss.n4923 vss.n4856 1534.21
R404 vss.n4921 vss.n4857 1534.21
R405 vss.n4910 vss.n4909 1534.21
R406 vss.n4900 vss.n4875 1534.21
R407 vss.n4898 vss.n4876 1534.21
R408 vss.n4887 vss.n4876 1534.21
R409 vss.n4890 vss.n4889 1534.21
R410 vss.n20222 vss.n20221 1505.26
R411 vss.n20221 vss.n20220 1505.26
R412 vss.n20100 vss.n19189 1505.26
R413 vss.n20091 vss.n19189 1505.26
R414 vss.n19975 vss.n19974 1505.26
R415 vss.n19974 vss.n19973 1505.26
R416 vss.n19844 vss.n19402 1505.26
R417 vss.n19728 vss.n19727 1505.26
R418 vss.n19727 vss.n19726 1505.26
R419 vss.n20356 vss.n20355 1505.26
R420 vss.n20355 vss.n20354 1505.26
R421 vss.n18954 vss.n17682 1505.26
R422 vss.n18945 vss.n17682 1505.26
R423 vss.n18829 vss.n18828 1505.26
R424 vss.n18828 vss.n18827 1505.26
R425 vss.n17901 vss.n17889 1505.26
R426 vss.n18704 vss.n17901 1505.26
R427 vss.n18588 vss.n18587 1505.26
R428 vss.n18587 vss.n18586 1505.26
R429 vss.n18114 vss.n18102 1505.26
R430 vss.n18463 vss.n18114 1505.26
R431 vss.n18347 vss.n18346 1505.26
R432 vss.n18346 vss.n18345 1505.26
R433 vss.n6832 vss.n6831 1505.26
R434 vss.n6831 vss.n6830 1505.26
R435 vss.n6710 vss.n5799 1505.26
R436 vss.n6701 vss.n5799 1505.26
R437 vss.n6585 vss.n6584 1505.26
R438 vss.n6584 vss.n6583 1505.26
R439 vss.n6454 vss.n6012 1505.26
R440 vss.n6338 vss.n6337 1505.26
R441 vss.n6337 vss.n6336 1505.26
R442 vss.n6966 vss.n6965 1505.26
R443 vss.n6965 vss.n6964 1505.26
R444 vss.n5564 vss.n4292 1505.26
R445 vss.n5555 vss.n4292 1505.26
R446 vss.n5439 vss.n5438 1505.26
R447 vss.n5438 vss.n5437 1505.26
R448 vss.n4511 vss.n4499 1505.26
R449 vss.n5314 vss.n4511 1505.26
R450 vss.n5198 vss.n5197 1505.26
R451 vss.n5197 vss.n5196 1505.26
R452 vss.n4724 vss.n4712 1505.26
R453 vss.n5073 vss.n4724 1505.26
R454 vss.n4957 vss.n4956 1505.26
R455 vss.n4956 vss.n4955 1505.26
R456 vss.n19402 ldomc_0.otaldom_0.nmoslm_0.vss 1418.42
R457 vss.n6012 bandgapmd_0.otam_1.nmoslm_0.vss 1418.42
R458 vss.n9201 vss.n9160 1049.71
R459 vss.n9198 vss.t328 1049.49
R460 vss.n9202 vss.n9201 1049.22
R461 vss.n18690 ldomc_0.otaldom_0.nmosrm_0.vss 897.368
R462 vss.n5300 vss 897.368
R463 vss.n13107 vss.n13106 883.464
R464 vss.n10683 vss.n10682 883.464
R465 vss.n14085 vss.n14084 883.464
R466 vss.n11845 vss.n11844 883.464
R467 vss.n10186 vss.n10185 676.517
R468 ldomc_0.otaldom_0.nmosrm_0.vss vss.n17914 636.842
R469 vss vss.n4524 636.842
R470 vss.n20412 vss.n17547 627.409
R471 vss.n7022 vss.n4157 627.409
R472 vss.n20408 vss.n20407 587.338
R473 vss.n7018 vss.n7017 587.338
R474 vss.n20319 vss.n20318 585.902
R475 vss.n6929 vss.n6928 585.902
R476 vss.n20309 vss.n20308 585.432
R477 vss.n6919 vss.n6918 585.432
R478 vss.n18275 vss.n18274 585
R479 vss.n18279 vss.n18275 585
R480 vss.n18209 vss.n18206 585
R481 vss.n18206 vss.n18205 585
R482 vss.n18198 vss.n18194 585
R483 vss.n18369 vss.n18194 585
R484 vss.n18383 vss.n18382 585
R485 vss.n18382 vss.n18381 585
R486 vss.n18174 vss.n18173 585
R487 vss.n18175 vss.n18174 585
R488 vss.n18104 vss.n18100 585
R489 vss.n18474 vss.n18100 585
R490 vss.n18488 vss.n18487 585
R491 vss.n18487 vss.n18486 585
R492 vss.n18077 vss.n18074 585
R493 vss.n18074 vss.n18073 585
R494 vss.n18066 vss.n18060 585
R495 vss.n18520 vss.n18060 585
R496 vss.n17996 vss.n17993 585
R497 vss.n17993 vss.n17992 585
R498 vss.n17985 vss.n17981 585
R499 vss.n18610 vss.n17981 585
R500 vss.n18624 vss.n18623 585
R501 vss.n18623 vss.n18622 585
R502 vss.n17961 vss.n17960 585
R503 vss.n17962 vss.n17961 585
R504 vss.n17891 vss.n17887 585
R505 vss.n18715 vss.n17887 585
R506 vss.n18729 vss.n18728 585
R507 vss.n18728 vss.n18727 585
R508 vss.n17864 vss.n17861 585
R509 vss.n17861 vss.n17860 585
R510 vss.n17853 vss.n17847 585
R511 vss.n18761 vss.n17847 585
R512 vss.n17783 vss.n17780 585
R513 vss.n17780 vss.n17779 585
R514 vss.n17772 vss.n17768 585
R515 vss.n18851 vss.n17768 585
R516 vss.n18865 vss.n18864 585
R517 vss.n18864 vss.n18863 585
R518 vss.n17748 vss.n17747 585
R519 vss.n17749 vss.n17748 585
R520 vss.n18958 vss.n18957 585
R521 vss.n18957 vss.n18956 585
R522 vss.n17667 vss.n17664 585
R523 vss.n17664 vss.n17663 585
R524 vss.n17655 vss.n17652 585
R525 vss.n18990 vss.n17652 585
R526 vss.n19002 vss.n17639 585
R527 vss.n17639 vss.n17638 585
R528 vss.n19028 vss.n19027 585
R529 vss.n19029 vss.n19028 585
R530 vss.n19026 vss.n17628 585
R531 vss.n17628 vss.n17627 585
R532 vss.n19016 vss.n19015 585
R533 vss.n19017 vss.n19016 585
R534 vss.n17633 vss.n17632 585
R535 vss.n19018 vss.n17633 585
R536 vss.n19013 vss.n19012 585
R537 vss.n19012 vss.n19011 585
R538 vss.n17637 vss.n17636 585
R539 vss.n19010 vss.n17637 585
R540 vss.n19001 vss.n19000 585
R541 vss.n19000 vss.n18999 585
R542 vss.n18996 vss.n18995 585
R543 vss.n18997 vss.n18996 585
R544 vss.n18994 vss.n17645 585
R545 vss.n17645 vss.n17644 585
R546 vss.n18988 vss.n18987 585
R547 vss.n18989 vss.n18988 585
R548 vss.n18981 vss.n18980 585
R549 vss.n18980 vss.n18979 585
R550 vss.n17662 vss.n17661 585
R551 vss.n18978 vss.n17662 585
R552 vss.n17670 vss.n17668 585
R553 vss.n17672 vss.n17670 585
R554 vss.n17675 vss.n17671 585
R555 vss.n18967 vss.n17671 585
R556 vss.n18965 vss.n18964 585
R557 vss.n18966 vss.n18965 585
R558 vss.n17681 vss.n17680 585
R559 vss.n18955 vss.n17681 585
R560 vss.n17688 vss.n17687 585
R561 vss.n18944 vss.n17688 585
R562 vss.n18942 vss.n18941 585
R563 vss.n18943 vss.n18942 585
R564 vss.n17696 vss.n17693 585
R565 vss.n17701 vss.n17696 585
R566 vss.n17699 vss.n17698 585
R567 vss.n17700 vss.n17699 585
R568 vss.n17697 vss.n17694 585
R569 vss.n18930 vss.n17697 585
R570 vss.n18928 vss.n18927 585
R571 vss.n18929 vss.n18928 585
R572 vss.n17707 vss.n17706 585
R573 vss.n18918 vss.n17707 585
R574 vss.n18921 vss.n18920 585
R575 vss.n18920 vss.n18919 585
R576 vss.n17712 vss.n17709 585
R577 vss.n17709 vss.n17708 585
R578 vss.n17718 vss.n17715 585
R579 vss.n17720 vss.n17718 585
R580 vss.n18905 vss.n18904 585
R581 vss.n18906 vss.n18905 585
R582 vss.n17719 vss.n17716 585
R583 vss.n18907 vss.n17719 585
R584 vss.n18898 vss.n18897 585
R585 vss.n18897 vss.n18896 585
R586 vss.n17726 vss.n17725 585
R587 vss.n18895 vss.n17726 585
R588 vss.n17736 vss.n17734 585
R589 vss.n17738 vss.n17736 585
R590 vss.n17731 vss.n17728 585
R591 vss.n17728 vss.n17727 585
R592 vss.n17737 vss.n17735 585
R593 vss.n18886 vss.n17737 585
R594 vss.n18884 vss.n18883 585
R595 vss.n18885 vss.n18884 585
R596 vss.n17745 vss.n17743 585
R597 vss.n17750 vss.n17745 585
R598 vss.n17753 vss.n17746 585
R599 vss.n18874 vss.n17746 585
R600 vss.n18872 vss.n18871 585
R601 vss.n18873 vss.n18872 585
R602 vss.n17759 vss.n17758 585
R603 vss.n18862 vss.n17759 585
R604 vss.n17764 vss.n17761 585
R605 vss.n17761 vss.n17760 585
R606 vss.n17767 vss.n17765 585
R607 vss.n17769 vss.n17767 585
R608 vss.n18849 vss.n18848 585
R609 vss.n18850 vss.n18849 585
R610 vss.n18842 vss.n18841 585
R611 vss.n18841 vss.n18840 585
R612 vss.n17778 vss.n17777 585
R613 vss.n18839 vss.n17778 585
R614 vss.n17786 vss.n17784 585
R615 vss.n17788 vss.n17786 585
R616 vss.n17793 vss.n17790 585
R617 vss.n17790 vss.n17789 585
R618 vss.n17799 vss.n17796 585
R619 vss.n17801 vss.n17799 585
R620 vss.n18815 vss.n18814 585
R621 vss.n18816 vss.n18815 585
R622 vss.n17800 vss.n17797 585
R623 vss.n18817 vss.n17800 585
R624 vss.n18808 vss.n18807 585
R625 vss.n18807 vss.n18806 585
R626 vss.n17807 vss.n17806 585
R627 vss.n18805 vss.n17807 585
R628 vss.n17818 vss.n17815 585
R629 vss.n17820 vss.n17818 585
R630 vss.n17812 vss.n17809 585
R631 vss.n17809 vss.n17808 585
R632 vss.n17819 vss.n17816 585
R633 vss.n18794 vss.n17819 585
R634 vss.n18792 vss.n18791 585
R635 vss.n18793 vss.n18792 585
R636 vss.n17826 vss.n17825 585
R637 vss.n18782 vss.n17826 585
R638 vss.n18785 vss.n18784 585
R639 vss.n18784 vss.n18783 585
R640 vss.n17831 vss.n17828 585
R641 vss.n17828 vss.n17827 585
R642 vss.n17837 vss.n17834 585
R643 vss.n17839 vss.n17837 585
R644 vss.n18769 vss.n18768 585
R645 vss.n18770 vss.n18769 585
R646 vss.n17838 vss.n17835 585
R647 vss.n18771 vss.n17838 585
R648 vss.n17848 vss.n17842 585
R649 vss.n17849 vss.n17848 585
R650 vss.n17846 vss.n17844 585
R651 vss.n17850 vss.n17846 585
R652 vss.n18759 vss.n18758 585
R653 vss.n18760 vss.n18759 585
R654 vss.n18752 vss.n18751 585
R655 vss.n18751 vss.n18750 585
R656 vss.n17859 vss.n17858 585
R657 vss.n18749 vss.n17859 585
R658 vss.n17867 vss.n17865 585
R659 vss.n17869 vss.n17867 585
R660 vss.n17872 vss.n17868 585
R661 vss.n18738 vss.n17868 585
R662 vss.n18736 vss.n18735 585
R663 vss.n18737 vss.n18736 585
R664 vss.n17878 vss.n17877 585
R665 vss.n18726 vss.n17878 585
R666 vss.n17883 vss.n17880 585
R667 vss.n17880 vss.n17879 585
R668 vss.n17886 vss.n17884 585
R669 vss.n17888 vss.n17886 585
R670 vss.n18713 vss.n18712 585
R671 vss.n18714 vss.n18713 585
R672 vss.n17900 vss.n17897 585
R673 vss.n18703 vss.n17900 585
R674 vss.n18701 vss.n18700 585
R675 vss.n18702 vss.n18701 585
R676 vss.n17909 vss.n17906 585
R677 vss.n17914 vss.n17909 585
R678 vss.n17912 vss.n17911 585
R679 vss.n17913 vss.n17912 585
R680 vss.n17910 vss.n17907 585
R681 vss.n18689 vss.n17910 585
R682 vss.n18687 vss.n18686 585
R683 vss.n18688 vss.n18687 585
R684 vss.n17920 vss.n17919 585
R685 vss.n18677 vss.n17920 585
R686 vss.n18680 vss.n18679 585
R687 vss.n18679 vss.n18678 585
R688 vss.n17925 vss.n17922 585
R689 vss.n17922 vss.n17921 585
R690 vss.n17931 vss.n17928 585
R691 vss.n17933 vss.n17931 585
R692 vss.n18664 vss.n18663 585
R693 vss.n18665 vss.n18664 585
R694 vss.n17932 vss.n17929 585
R695 vss.n18666 vss.n17932 585
R696 vss.n18657 vss.n18656 585
R697 vss.n18656 vss.n18655 585
R698 vss.n17939 vss.n17938 585
R699 vss.n18654 vss.n17939 585
R700 vss.n17949 vss.n17947 585
R701 vss.n17951 vss.n17949 585
R702 vss.n17944 vss.n17941 585
R703 vss.n17941 vss.n17940 585
R704 vss.n17950 vss.n17948 585
R705 vss.n18645 vss.n17950 585
R706 vss.n18643 vss.n18642 585
R707 vss.n18644 vss.n18643 585
R708 vss.n17958 vss.n17956 585
R709 vss.n17963 vss.n17958 585
R710 vss.n17966 vss.n17959 585
R711 vss.n18633 vss.n17959 585
R712 vss.n18631 vss.n18630 585
R713 vss.n18632 vss.n18631 585
R714 vss.n17972 vss.n17971 585
R715 vss.n18621 vss.n17972 585
R716 vss.n17977 vss.n17974 585
R717 vss.n17974 vss.n17973 585
R718 vss.n17980 vss.n17978 585
R719 vss.n17982 vss.n17980 585
R720 vss.n18608 vss.n18607 585
R721 vss.n18609 vss.n18608 585
R722 vss.n18601 vss.n18600 585
R723 vss.n18600 vss.n18599 585
R724 vss.n17991 vss.n17990 585
R725 vss.n18598 vss.n17991 585
R726 vss.n17999 vss.n17997 585
R727 vss.n18001 vss.n17999 585
R728 vss.n18006 vss.n18003 585
R729 vss.n18003 vss.n18002 585
R730 vss.n18012 vss.n18009 585
R731 vss.n18014 vss.n18012 585
R732 vss.n18574 vss.n18573 585
R733 vss.n18575 vss.n18574 585
R734 vss.n18013 vss.n18010 585
R735 vss.n18576 vss.n18013 585
R736 vss.n18567 vss.n18566 585
R737 vss.n18566 vss.n18565 585
R738 vss.n18020 vss.n18019 585
R739 vss.n18564 vss.n18020 585
R740 vss.n18031 vss.n18028 585
R741 vss.n18033 vss.n18031 585
R742 vss.n18025 vss.n18022 585
R743 vss.n18022 vss.n18021 585
R744 vss.n18032 vss.n18029 585
R745 vss.n18553 vss.n18032 585
R746 vss.n18551 vss.n18550 585
R747 vss.n18552 vss.n18551 585
R748 vss.n18039 vss.n18038 585
R749 vss.n18541 vss.n18039 585
R750 vss.n18544 vss.n18543 585
R751 vss.n18543 vss.n18542 585
R752 vss.n18044 vss.n18041 585
R753 vss.n18041 vss.n18040 585
R754 vss.n18050 vss.n18047 585
R755 vss.n18052 vss.n18050 585
R756 vss.n18528 vss.n18527 585
R757 vss.n18529 vss.n18528 585
R758 vss.n18051 vss.n18048 585
R759 vss.n18530 vss.n18051 585
R760 vss.n18061 vss.n18055 585
R761 vss.n18062 vss.n18061 585
R762 vss.n18059 vss.n18057 585
R763 vss.n18063 vss.n18059 585
R764 vss.n18518 vss.n18517 585
R765 vss.n18519 vss.n18518 585
R766 vss.n18511 vss.n18510 585
R767 vss.n18510 vss.n18509 585
R768 vss.n18072 vss.n18071 585
R769 vss.n18508 vss.n18072 585
R770 vss.n18080 vss.n18078 585
R771 vss.n18082 vss.n18080 585
R772 vss.n18085 vss.n18081 585
R773 vss.n18497 vss.n18081 585
R774 vss.n18495 vss.n18494 585
R775 vss.n18496 vss.n18495 585
R776 vss.n18091 vss.n18090 585
R777 vss.n18485 vss.n18091 585
R778 vss.n18096 vss.n18093 585
R779 vss.n18093 vss.n18092 585
R780 vss.n18099 vss.n18097 585
R781 vss.n18101 vss.n18099 585
R782 vss.n18472 vss.n18471 585
R783 vss.n18473 vss.n18472 585
R784 vss.n18113 vss.n18110 585
R785 vss.n18462 vss.n18113 585
R786 vss.n18460 vss.n18459 585
R787 vss.n18461 vss.n18460 585
R788 vss.n18122 vss.n18119 585
R789 vss.n18127 vss.n18122 585
R790 vss.n18125 vss.n18124 585
R791 vss.n18126 vss.n18125 585
R792 vss.n18123 vss.n18120 585
R793 vss.n18448 vss.n18123 585
R794 vss.n18446 vss.n18445 585
R795 vss.n18447 vss.n18446 585
R796 vss.n18133 vss.n18132 585
R797 vss.n18436 vss.n18133 585
R798 vss.n18439 vss.n18438 585
R799 vss.n18438 vss.n18437 585
R800 vss.n18138 vss.n18135 585
R801 vss.n18135 vss.n18134 585
R802 vss.n18144 vss.n18141 585
R803 vss.n18146 vss.n18144 585
R804 vss.n18423 vss.n18422 585
R805 vss.n18424 vss.n18423 585
R806 vss.n18145 vss.n18142 585
R807 vss.n18425 vss.n18145 585
R808 vss.n18416 vss.n18415 585
R809 vss.n18415 vss.n18414 585
R810 vss.n18152 vss.n18151 585
R811 vss.n18413 vss.n18152 585
R812 vss.n18162 vss.n18160 585
R813 vss.n18164 vss.n18162 585
R814 vss.n18157 vss.n18154 585
R815 vss.n18154 vss.n18153 585
R816 vss.n18163 vss.n18161 585
R817 vss.n18404 vss.n18163 585
R818 vss.n18402 vss.n18401 585
R819 vss.n18403 vss.n18402 585
R820 vss.n18171 vss.n18169 585
R821 vss.n18176 vss.n18171 585
R822 vss.n18179 vss.n18172 585
R823 vss.n18392 vss.n18172 585
R824 vss.n18390 vss.n18389 585
R825 vss.n18391 vss.n18390 585
R826 vss.n18185 vss.n18184 585
R827 vss.n18380 vss.n18185 585
R828 vss.n18190 vss.n18187 585
R829 vss.n18187 vss.n18186 585
R830 vss.n18193 vss.n18191 585
R831 vss.n18195 vss.n18193 585
R832 vss.n18367 vss.n18366 585
R833 vss.n18368 vss.n18367 585
R834 vss.n18360 vss.n18359 585
R835 vss.n18359 vss.n18358 585
R836 vss.n18204 vss.n18203 585
R837 vss.n18357 vss.n18204 585
R838 vss.n18212 vss.n18210 585
R839 vss.n18214 vss.n18212 585
R840 vss.n18219 vss.n18216 585
R841 vss.n18216 vss.n18215 585
R842 vss.n18225 vss.n18222 585
R843 vss.n18227 vss.n18225 585
R844 vss.n18333 vss.n18332 585
R845 vss.n18334 vss.n18333 585
R846 vss.n18226 vss.n18223 585
R847 vss.n18335 vss.n18226 585
R848 vss.n18326 vss.n18325 585
R849 vss.n18325 vss.n18324 585
R850 vss.n18233 vss.n18232 585
R851 vss.n18323 vss.n18233 585
R852 vss.n18244 vss.n18241 585
R853 vss.n18246 vss.n18244 585
R854 vss.n18238 vss.n18235 585
R855 vss.n18235 vss.n18234 585
R856 vss.n18245 vss.n18242 585
R857 vss.n18312 vss.n18245 585
R858 vss.n18310 vss.n18309 585
R859 vss.n18311 vss.n18310 585
R860 vss.n18252 vss.n18251 585
R861 vss.n18300 vss.n18252 585
R862 vss.n18303 vss.n18302 585
R863 vss.n18302 vss.n18301 585
R864 vss.n18257 vss.n18254 585
R865 vss.n18254 vss.n18253 585
R866 vss.n18263 vss.n18260 585
R867 vss.n18265 vss.n18263 585
R868 vss.n18287 vss.n18286 585
R869 vss.n18288 vss.n18287 585
R870 vss.n18264 vss.n18261 585
R871 vss.n18289 vss.n18264 585
R872 vss.n18276 vss.n18268 585
R873 vss.n18277 vss.n18276 585
R874 vss.n18272 vss.n18270 585
R875 vss.n18278 vss.n18272 585
R876 vss.n17625 vss.n17624 585
R877 vss.n19603 vss.n19591 585
R878 vss.n19603 vss.n19596 585
R879 vss.n17592 vss.n17587 585
R880 vss.n17594 vss.n17592 585
R881 vss.n20352 vss.n17595 585
R882 vss.n20347 vss.n20346 585
R883 vss.n20341 vss.n17598 585
R884 vss.n20336 vss.n20335 585
R885 vss.n20330 vss.n20329 585
R886 vss.n20325 vss.n17603 585
R887 vss.n20321 vss.n20320 585
R888 vss.n17614 vss.n17611 585
R889 vss.n20302 vss.n17615 585
R890 vss.n20324 vss.n17575 585
R891 vss.n20324 vss.n20323 585
R892 vss.n20328 vss.n17602 585
R893 vss.n20334 vss.n20333 585
R894 vss.n19611 vss.n19610 585
R895 vss.n19610 vss.n19609 585
R896 vss.n20350 vss.n20349 585
R897 vss.n20344 vss.n17597 585
R898 vss.n20340 vss.n20339 585
R899 vss.n19633 vss.n19632 585
R900 vss.n19632 vss.n19631 585
R901 vss.n19648 vss.n19647 585
R902 vss.n19649 vss.n19648 585
R903 vss.n19665 vss.n19664 585
R904 vss.n19664 vss.n19663 585
R905 vss.n19741 vss.n19740 585
R906 vss.n19740 vss.n19739 585
R907 vss.n19478 vss.n19475 585
R908 vss.n19475 vss.n19474 585
R909 vss.n19467 vss.n19460 585
R910 vss.n19773 vss.n19460 585
R911 vss.n19451 vss.n19449 585
R912 vss.n19785 vss.n19451 585
R913 vss.n19389 vss.n19385 585
R914 vss.n19866 vss.n19385 585
R915 vss.n19880 vss.n19879 585
R916 vss.n19879 vss.n19878 585
R917 vss.n19895 vss.n19894 585
R918 vss.n19896 vss.n19895 585
R919 vss.n19912 vss.n19911 585
R920 vss.n19911 vss.n19910 585
R921 vss.n19988 vss.n19987 585
R922 vss.n19987 vss.n19986 585
R923 vss.n19271 vss.n19268 585
R924 vss.n19268 vss.n19267 585
R925 vss.n19260 vss.n19253 585
R926 vss.n20020 vss.n19253 585
R927 vss.n19244 vss.n19242 585
R928 vss.n20032 vss.n19244 585
R929 vss.n19182 vss.n19178 585
R930 vss.n20113 vss.n19178 585
R931 vss.n20127 vss.n20126 585
R932 vss.n20126 vss.n20125 585
R933 vss.n20142 vss.n20141 585
R934 vss.n20143 vss.n20142 585
R935 vss.n20159 vss.n20158 585
R936 vss.n20158 vss.n20157 585
R937 vss.n20235 vss.n20234 585
R938 vss.n20234 vss.n20233 585
R939 vss.n19064 vss.n19061 585
R940 vss.n19061 vss.n19060 585
R941 vss.n19052 vss.n19049 585
R942 vss.n20267 vss.n19049 585
R943 vss.n20279 vss.n19037 585
R944 vss.n19037 vss.n19036 585
R945 vss.n20293 vss.n20292 585
R946 vss.n20294 vss.n20293 585
R947 vss.n17621 vss.n17617 585
R948 vss.n20286 vss.n20285 585
R949 vss.n20285 vss.n20284 585
R950 vss.n19035 vss.n19034 585
R951 vss.n20283 vss.n19035 585
R952 vss.n20278 vss.n20277 585
R953 vss.n20277 vss.n20276 585
R954 vss.n20273 vss.n20272 585
R955 vss.n20274 vss.n20273 585
R956 vss.n20271 vss.n19041 585
R957 vss.n19041 vss.n19040 585
R958 vss.n20265 vss.n20264 585
R959 vss.n20266 vss.n20265 585
R960 vss.n20258 vss.n20257 585
R961 vss.n20257 vss.n20256 585
R962 vss.n19059 vss.n19058 585
R963 vss.n20255 vss.n19059 585
R964 vss.n19067 vss.n19065 585
R965 vss.n19069 vss.n19067 585
R966 vss.n19072 vss.n19068 585
R967 vss.n20244 vss.n19068 585
R968 vss.n20242 vss.n20241 585
R969 vss.n20243 vss.n20242 585
R970 vss.n19078 vss.n19077 585
R971 vss.n20232 vss.n19078 585
R972 vss.n19083 vss.n19080 585
R973 vss.n19080 vss.n19079 585
R974 vss.n19086 vss.n19084 585
R975 vss.n19088 vss.n19086 585
R976 vss.n19099 vss.n19096 585
R977 vss.n19101 vss.n19099 585
R978 vss.n19093 vss.n19090 585
R979 vss.n19090 vss.n19089 585
R980 vss.n19100 vss.n19097 585
R981 vss.n20210 vss.n19100 585
R982 vss.n20208 vss.n20207 585
R983 vss.n20209 vss.n20208 585
R984 vss.n19107 vss.n19106 585
R985 vss.n20198 vss.n19107 585
R986 vss.n20201 vss.n20200 585
R987 vss.n20200 vss.n20199 585
R988 vss.n19112 vss.n19109 585
R989 vss.n19109 vss.n19108 585
R990 vss.n19118 vss.n19115 585
R991 vss.n19120 vss.n19118 585
R992 vss.n20185 vss.n20184 585
R993 vss.n20186 vss.n20185 585
R994 vss.n19119 vss.n19116 585
R995 vss.n20187 vss.n19119 585
R996 vss.n20178 vss.n20177 585
R997 vss.n20177 vss.n20176 585
R998 vss.n19126 vss.n19125 585
R999 vss.n20175 vss.n19126 585
R1000 vss.n19137 vss.n19134 585
R1001 vss.n19139 vss.n19137 585
R1002 vss.n19131 vss.n19128 585
R1003 vss.n19128 vss.n19127 585
R1004 vss.n19138 vss.n19135 585
R1005 vss.n20164 vss.n19138 585
R1006 vss.n20162 vss.n20161 585
R1007 vss.n20163 vss.n20162 585
R1008 vss.n19144 vss.n19143 585
R1009 vss.n20156 vss.n19144 585
R1010 vss.n20148 vss.n19146 585
R1011 vss.n19146 vss.n19145 585
R1012 vss.n20147 vss.n20146 585
R1013 vss.n20146 vss.n20145 585
R1014 vss.n20140 vss.n19152 585
R1015 vss.n19152 vss.n19151 585
R1016 vss.n19162 vss.n19159 585
R1017 vss.n20136 vss.n19159 585
R1018 vss.n20134 vss.n20133 585
R1019 vss.n20135 vss.n20134 585
R1020 vss.n19169 vss.n19168 585
R1021 vss.n20124 vss.n19169 585
R1022 vss.n19174 vss.n19171 585
R1023 vss.n19171 vss.n19170 585
R1024 vss.n19177 vss.n19175 585
R1025 vss.n19179 vss.n19177 585
R1026 vss.n20111 vss.n20110 585
R1027 vss.n20112 vss.n20111 585
R1028 vss.n20104 vss.n20103 585
R1029 vss.n20103 vss.n20102 585
R1030 vss.n19188 vss.n19187 585
R1031 vss.n20101 vss.n19188 585
R1032 vss.n20088 vss.n20087 585
R1033 vss.n20089 vss.n20088 585
R1034 vss.n19195 vss.n19194 585
R1035 vss.n20090 vss.n19195 585
R1036 vss.n19206 vss.n19205 585
R1037 vss.n19207 vss.n19206 585
R1038 vss.n19203 vss.n19200 585
R1039 vss.n19208 vss.n19203 585
R1040 vss.n20074 vss.n20073 585
R1041 vss.n20075 vss.n20074 585
R1042 vss.n19204 vss.n19201 585
R1043 vss.n20076 vss.n19204 585
R1044 vss.n20067 vss.n20066 585
R1045 vss.n20066 vss.n20065 585
R1046 vss.n19214 vss.n19213 585
R1047 vss.n20064 vss.n19214 585
R1048 vss.n19225 vss.n19222 585
R1049 vss.n19227 vss.n19225 585
R1050 vss.n19219 vss.n19216 585
R1051 vss.n19216 vss.n19215 585
R1052 vss.n19226 vss.n19223 585
R1053 vss.n20053 vss.n19226 585
R1054 vss.n20051 vss.n20050 585
R1055 vss.n20052 vss.n20051 585
R1056 vss.n19233 vss.n19232 585
R1057 vss.n20041 vss.n19233 585
R1058 vss.n20044 vss.n20043 585
R1059 vss.n20043 vss.n20042 585
R1060 vss.n19238 vss.n19235 585
R1061 vss.n19235 vss.n19234 585
R1062 vss.n19243 vss.n19241 585
R1063 vss.n19245 vss.n19243 585
R1064 vss.n20030 vss.n20029 585
R1065 vss.n20031 vss.n20030 585
R1066 vss.n19255 vss.n19254 585
R1067 vss.n19256 vss.n19255 585
R1068 vss.n19252 vss.n19250 585
R1069 vss.n19257 vss.n19252 585
R1070 vss.n20018 vss.n20017 585
R1071 vss.n20019 vss.n20018 585
R1072 vss.n20011 vss.n20010 585
R1073 vss.n20010 vss.n20009 585
R1074 vss.n19266 vss.n19265 585
R1075 vss.n20008 vss.n19266 585
R1076 vss.n19274 vss.n19272 585
R1077 vss.n19276 vss.n19274 585
R1078 vss.n19279 vss.n19275 585
R1079 vss.n19997 vss.n19275 585
R1080 vss.n19995 vss.n19994 585
R1081 vss.n19996 vss.n19995 585
R1082 vss.n19285 vss.n19284 585
R1083 vss.n19985 vss.n19285 585
R1084 vss.n19290 vss.n19287 585
R1085 vss.n19287 vss.n19286 585
R1086 vss.n19293 vss.n19291 585
R1087 vss.n19295 vss.n19293 585
R1088 vss.n19306 vss.n19303 585
R1089 vss.n19308 vss.n19306 585
R1090 vss.n19300 vss.n19297 585
R1091 vss.n19297 vss.n19296 585
R1092 vss.n19307 vss.n19304 585
R1093 vss.n19963 vss.n19307 585
R1094 vss.n19961 vss.n19960 585
R1095 vss.n19962 vss.n19961 585
R1096 vss.n19314 vss.n19313 585
R1097 vss.n19951 vss.n19314 585
R1098 vss.n19954 vss.n19953 585
R1099 vss.n19953 vss.n19952 585
R1100 vss.n19319 vss.n19316 585
R1101 vss.n19316 vss.n19315 585
R1102 vss.n19325 vss.n19322 585
R1103 vss.n19327 vss.n19325 585
R1104 vss.n19938 vss.n19937 585
R1105 vss.n19939 vss.n19938 585
R1106 vss.n19326 vss.n19323 585
R1107 vss.n19940 vss.n19326 585
R1108 vss.n19931 vss.n19930 585
R1109 vss.n19930 vss.n19929 585
R1110 vss.n19333 vss.n19332 585
R1111 vss.n19928 vss.n19333 585
R1112 vss.n19344 vss.n19341 585
R1113 vss.n19346 vss.n19344 585
R1114 vss.n19338 vss.n19335 585
R1115 vss.n19335 vss.n19334 585
R1116 vss.n19345 vss.n19342 585
R1117 vss.n19917 vss.n19345 585
R1118 vss.n19915 vss.n19914 585
R1119 vss.n19916 vss.n19915 585
R1120 vss.n19351 vss.n19350 585
R1121 vss.n19909 vss.n19351 585
R1122 vss.n19901 vss.n19353 585
R1123 vss.n19353 vss.n19352 585
R1124 vss.n19900 vss.n19899 585
R1125 vss.n19899 vss.n19898 585
R1126 vss.n19893 vss.n19359 585
R1127 vss.n19359 vss.n19358 585
R1128 vss.n19369 vss.n19366 585
R1129 vss.n19889 vss.n19366 585
R1130 vss.n19887 vss.n19886 585
R1131 vss.n19888 vss.n19887 585
R1132 vss.n19376 vss.n19375 585
R1133 vss.n19877 vss.n19376 585
R1134 vss.n19381 vss.n19378 585
R1135 vss.n19378 vss.n19377 585
R1136 vss.n19384 vss.n19382 585
R1137 vss.n19386 vss.n19384 585
R1138 vss.n19864 vss.n19863 585
R1139 vss.n19865 vss.n19864 585
R1140 vss.n19857 vss.n19856 585
R1141 vss.n19856 vss.n19855 585
R1142 vss.n19395 vss.n19394 585
R1143 vss.n19854 vss.n19395 585
R1144 vss.n19841 vss.n19840 585
R1145 vss.n19842 vss.n19841 585
R1146 vss.n19401 vss.n19400 585
R1147 vss.n19843 vss.n19401 585
R1148 vss.n19413 vss.n19412 585
R1149 vss.n19414 vss.n19413 585
R1150 vss.n19410 vss.n19407 585
R1151 vss.n19415 vss.n19410 585
R1152 vss.n19827 vss.n19826 585
R1153 vss.n19828 vss.n19827 585
R1154 vss.n19411 vss.n19408 585
R1155 vss.n19829 vss.n19411 585
R1156 vss.n19820 vss.n19819 585
R1157 vss.n19819 vss.n19818 585
R1158 vss.n19421 vss.n19420 585
R1159 vss.n19817 vss.n19421 585
R1160 vss.n19432 vss.n19429 585
R1161 vss.n19434 vss.n19432 585
R1162 vss.n19426 vss.n19423 585
R1163 vss.n19423 vss.n19422 585
R1164 vss.n19433 vss.n19430 585
R1165 vss.n19806 vss.n19433 585
R1166 vss.n19804 vss.n19803 585
R1167 vss.n19805 vss.n19804 585
R1168 vss.n19440 vss.n19439 585
R1169 vss.n19794 vss.n19440 585
R1170 vss.n19797 vss.n19796 585
R1171 vss.n19796 vss.n19795 585
R1172 vss.n19445 vss.n19442 585
R1173 vss.n19442 vss.n19441 585
R1174 vss.n19450 vss.n19448 585
R1175 vss.n19452 vss.n19450 585
R1176 vss.n19783 vss.n19782 585
R1177 vss.n19784 vss.n19783 585
R1178 vss.n19462 vss.n19461 585
R1179 vss.n19463 vss.n19462 585
R1180 vss.n19459 vss.n19457 585
R1181 vss.n19464 vss.n19459 585
R1182 vss.n19771 vss.n19770 585
R1183 vss.n19772 vss.n19771 585
R1184 vss.n19764 vss.n19763 585
R1185 vss.n19763 vss.n19762 585
R1186 vss.n19473 vss.n19472 585
R1187 vss.n19761 vss.n19473 585
R1188 vss.n19481 vss.n19479 585
R1189 vss.n19483 vss.n19481 585
R1190 vss.n19486 vss.n19482 585
R1191 vss.n19750 vss.n19482 585
R1192 vss.n19748 vss.n19747 585
R1193 vss.n19749 vss.n19748 585
R1194 vss.n19492 vss.n19491 585
R1195 vss.n19738 vss.n19492 585
R1196 vss.n19497 vss.n19494 585
R1197 vss.n19494 vss.n19493 585
R1198 vss.n19500 vss.n19498 585
R1199 vss.n19502 vss.n19500 585
R1200 vss.n19513 vss.n19510 585
R1201 vss.n19515 vss.n19513 585
R1202 vss.n19507 vss.n19504 585
R1203 vss.n19504 vss.n19503 585
R1204 vss.n19514 vss.n19511 585
R1205 vss.n19716 vss.n19514 585
R1206 vss.n19714 vss.n19713 585
R1207 vss.n19715 vss.n19714 585
R1208 vss.n19521 vss.n19520 585
R1209 vss.n19704 vss.n19521 585
R1210 vss.n19707 vss.n19706 585
R1211 vss.n19706 vss.n19705 585
R1212 vss.n19526 vss.n19523 585
R1213 vss.n19523 vss.n19522 585
R1214 vss.n19532 vss.n19529 585
R1215 vss.n19534 vss.n19532 585
R1216 vss.n19691 vss.n19690 585
R1217 vss.n19692 vss.n19691 585
R1218 vss.n19533 vss.n19530 585
R1219 vss.n19693 vss.n19533 585
R1220 vss.n19684 vss.n19683 585
R1221 vss.n19683 vss.n19682 585
R1222 vss.n19540 vss.n19539 585
R1223 vss.n19681 vss.n19540 585
R1224 vss.n19551 vss.n19548 585
R1225 vss.n19553 vss.n19551 585
R1226 vss.n19545 vss.n19542 585
R1227 vss.n19542 vss.n19541 585
R1228 vss.n19552 vss.n19549 585
R1229 vss.n19670 vss.n19552 585
R1230 vss.n19668 vss.n19667 585
R1231 vss.n19669 vss.n19668 585
R1232 vss.n19558 vss.n19557 585
R1233 vss.n19662 vss.n19558 585
R1234 vss.n19654 vss.n19560 585
R1235 vss.n19560 vss.n19559 585
R1236 vss.n19653 vss.n19652 585
R1237 vss.n19652 vss.n19651 585
R1238 vss.n19646 vss.n19566 585
R1239 vss.n19566 vss.n19565 585
R1240 vss.n19576 vss.n19573 585
R1241 vss.n19642 vss.n19573 585
R1242 vss.n19640 vss.n19639 585
R1243 vss.n19641 vss.n19640 585
R1244 vss.n19583 vss.n19582 585
R1245 vss.n19630 vss.n19583 585
R1246 vss.n19597 vss.n19585 585
R1247 vss.n19585 vss.n19584 585
R1248 vss.n19599 vss.n19598 585
R1249 vss.n19600 vss.n19599 585
R1250 vss.n19606 vss.n19605 585
R1251 vss.n19607 vss.n19606 585
R1252 vss.n20299 vss.n17616 585
R1253 vss.n20298 vss.n20297 585
R1254 vss.n20310 vss.n20309 585
R1255 vss.n20314 vss.n20313 585
R1256 vss.n20313 vss.n20312 585
R1257 vss.n20319 vss.n17606 585
R1258 vss.n20410 vss.n17547 585
R1259 vss.n12555 vss.n12554 585
R1260 vss.n12548 vss.n12547 585
R1261 vss.n11177 vss.n11176 585
R1262 vss.n10999 vss.n10998 585
R1263 vss.n10979 vss.n10978 585
R1264 vss.n10969 vss.n10968 585
R1265 vss.n12017 vss.n12016 585
R1266 vss.n12040 vss.n12039 585
R1267 vss.n12168 vss.n12167 585
R1268 vss.n12116 vss.n12115 585
R1269 vss.n12118 vss.n12117 585
R1270 vss.n12128 vss.n12127 585
R1271 vss.n12126 vss.n12125 585
R1272 vss.n12140 vss.n12139 585
R1273 vss.n12142 vss.n12141 585
R1274 vss.n12182 vss.n12181 585
R1275 vss.n12196 vss.n12195 585
R1276 vss.n12223 vss.n12222 585
R1277 vss.n12067 vss.n12066 585
R1278 vss.n12050 vss.n12049 585
R1279 vss.n10796 vss.n10795 585
R1280 vss.n12000 vss.n11999 585
R1281 vss.n10852 vss.n10851 585
R1282 vss.n11972 vss.n11971 585
R1283 vss.n10878 vss.n10877 585
R1284 vss.n10876 vss.n10875 585
R1285 vss.n11974 vss.n11973 585
R1286 vss.n11986 vss.n11985 585
R1287 vss.n11944 vss.n11943 585
R1288 vss.n11946 vss.n11945 585
R1289 vss.n11920 vss.n11919 585
R1290 vss.n11918 vss.n11917 585
R1291 vss.n11320 vss.n11319 585
R1292 vss.n11295 vss.n11294 585
R1293 vss.n11279 vss.n11278 585
R1294 vss.n11253 vss.n11252 585
R1295 vss.n10959 vss.n10958 585
R1296 vss.n11193 vss.n11192 585
R1297 vss.n11156 vss.n11155 585
R1298 vss.n14369 vss.n14368 585
R1299 vss.n14308 vss.n14307 585
R1300 vss.n13876 vss.n13875 585
R1301 vss.n13849 vss.n13848 585
R1302 vss.n11660 vss.n11659 585
R1303 vss.n11821 vss.n11820 585
R1304 vss.n11780 vss.n11779 585
R1305 vss.n11716 vss.n11715 585
R1306 vss.n11080 vss.n11079 585
R1307 vss.n11090 vss.n11089 585
R1308 vss.n11070 vss.n11069 585
R1309 vss.n11060 vss.n11059 585
R1310 vss.n11114 vss.n11113 585
R1311 vss.n11124 vss.n11123 585
R1312 vss.n11743 vss.n11742 585
R1313 vss.n11796 vss.n11795 585
R1314 vss.n11671 vss.n11670 585
R1315 vss.n11673 vss.n11672 585
R1316 vss.n11662 vss.n11661 585
R1317 vss.n11633 vss.n11632 585
R1318 vss.n11635 vss.n11634 585
R1319 vss.n11624 vss.n11623 585
R1320 vss.n11622 vss.n11621 585
R1321 vss.n11608 vss.n11607 585
R1322 vss.n14007 vss.n14006 585
R1323 vss.n13986 vss.n13985 585
R1324 vss.n14048 vss.n14047 585
R1325 vss.n14070 vss.n14069 585
R1326 vss.n13822 vss.n13821 585
R1327 vss.n13832 vss.n13831 585
R1328 vss.n13910 vss.n13909 585
R1329 vss.n14294 vss.n14293 585
R1330 vss.n14334 vss.n14333 585
R1331 vss.n14336 vss.n14335 585
R1332 vss.n14371 vss.n14370 585
R1333 vss.n14415 vss.n14414 585
R1334 vss.n14417 vss.n14416 585
R1335 vss.n14257 vss.n14256 585
R1336 vss.n14812 vss.n14811 585
R1337 vss.n14784 vss.n14783 585
R1338 vss.n14737 vss.n14736 585
R1339 vss.n13363 vss.n13362 585
R1340 vss.n13383 vss.n13382 585
R1341 vss.n14678 vss.n14677 585
R1342 vss.n13528 vss.n13527 585
R1343 vss.n14611 vss.n14610 585
R1344 vss.n14551 vss.n14550 585
R1345 vss.n14519 vss.n14518 585
R1346 vss.n14465 vss.n14464 585
R1347 vss.n14195 vss.n14194 585
R1348 vss.n14205 vss.n14204 585
R1349 vss.n14247 vss.n14246 585
R1350 vss.n14237 vss.n14236 585
R1351 vss.n14217 vss.n14216 585
R1352 vss.n14227 vss.n14226 585
R1353 vss.n14185 vss.n14184 585
R1354 vss.n14503 vss.n14502 585
R1355 vss.n14536 vss.n14535 585
R1356 vss.n14553 vss.n14552 585
R1357 vss.n14591 vss.n14590 585
R1358 vss.n14593 vss.n14592 585
R1359 vss.n13541 vss.n13540 585
R1360 vss.n13539 vss.n13538 585
R1361 vss.n14613 vss.n14612 585
R1362 vss.n14625 vss.n14624 585
R1363 vss.n13511 vss.n13510 585
R1364 vss.n14692 vss.n14691 585
R1365 vss.n13347 vss.n13346 585
R1366 vss.n14770 vss.n14769 585
R1367 vss.n14798 vss.n14797 585
R1368 vss.n14814 vss.n14813 585
R1369 vss.n13254 vss.n13253 585
R1370 vss.n13256 vss.n13255 585
R1371 vss.n13272 vss.n13271 585
R1372 vss.n13270 vss.n13269 585
R1373 vss.n12886 vss.n12885 585
R1374 vss.n14831 vss.n14830 585
R1375 vss.n14833 vss.n14832 585
R1376 vss.n14861 vss.n14860 585
R1377 vss.n14859 vss.n14858 585
R1378 vss.n14902 vss.n14901 585
R1379 vss.n14904 vss.n14903 585
R1380 vss.n14889 vss.n14888 585
R1381 vss.n14874 vss.n14873 585
R1382 vss.n12837 vss.n12836 585
R1383 vss.n12852 vss.n12851 585
R1384 vss.n12867 vss.n12866 585
R1385 vss.n12888 vss.n12887 585
R1386 vss.n12917 vss.n12916 585
R1387 vss.n12910 vss.n12909 585
R1388 vss.n12811 vss.n12810 585
R1389 vss.n12804 vss.n12803 585
R1390 vss.n15052 vss.n15051 585
R1391 vss.n15045 vss.n15044 585
R1392 vss.n15050 vss.n15049 585
R1393 vss.n12477 vss.n12476 585
R1394 vss.n10484 vss.n10483 585
R1395 vss.n10486 vss.n10485 585
R1396 vss.n10516 vss.n10515 585
R1397 vss.n10514 vss.n10513 585
R1398 vss.n10544 vss.n10543 585
R1399 vss.n10546 vss.n10545 585
R1400 vss.n12701 vss.n12700 585
R1401 vss.n12685 vss.n12684 585
R1402 vss.n12668 vss.n12667 585
R1403 vss.n12652 vss.n12651 585
R1404 vss.n12462 vss.n12461 585
R1405 vss.n12479 vss.n12478 585
R1406 vss.n12504 vss.n12503 585
R1407 vss.n12497 vss.n12496 585
R1408 vss.n4885 vss.n4884 585
R1409 vss.n4889 vss.n4885 585
R1410 vss.n4819 vss.n4816 585
R1411 vss.n4816 vss.n4815 585
R1412 vss.n4808 vss.n4804 585
R1413 vss.n4979 vss.n4804 585
R1414 vss.n4993 vss.n4992 585
R1415 vss.n4992 vss.n4991 585
R1416 vss.n4784 vss.n4783 585
R1417 vss.n4785 vss.n4784 585
R1418 vss.n4714 vss.n4710 585
R1419 vss.n5084 vss.n4710 585
R1420 vss.n5098 vss.n5097 585
R1421 vss.n5097 vss.n5096 585
R1422 vss.n4687 vss.n4684 585
R1423 vss.n4684 vss.n4683 585
R1424 vss.n4676 vss.n4670 585
R1425 vss.n5130 vss.n4670 585
R1426 vss.n4606 vss.n4603 585
R1427 vss.n4603 vss.n4602 585
R1428 vss.n4595 vss.n4591 585
R1429 vss.n5220 vss.n4591 585
R1430 vss.n5234 vss.n5233 585
R1431 vss.n5233 vss.n5232 585
R1432 vss.n4571 vss.n4570 585
R1433 vss.n4572 vss.n4571 585
R1434 vss.n4501 vss.n4497 585
R1435 vss.n5325 vss.n4497 585
R1436 vss.n5339 vss.n5338 585
R1437 vss.n5338 vss.n5337 585
R1438 vss.n4474 vss.n4471 585
R1439 vss.n4471 vss.n4470 585
R1440 vss.n4463 vss.n4457 585
R1441 vss.n5371 vss.n4457 585
R1442 vss.n4393 vss.n4390 585
R1443 vss.n4390 vss.n4389 585
R1444 vss.n4382 vss.n4378 585
R1445 vss.n5461 vss.n4378 585
R1446 vss.n5475 vss.n5474 585
R1447 vss.n5474 vss.n5473 585
R1448 vss.n4358 vss.n4357 585
R1449 vss.n4359 vss.n4358 585
R1450 vss.n5568 vss.n5567 585
R1451 vss.n5567 vss.n5566 585
R1452 vss.n4277 vss.n4274 585
R1453 vss.n4274 vss.n4273 585
R1454 vss.n4265 vss.n4262 585
R1455 vss.n5600 vss.n4262 585
R1456 vss.n5612 vss.n4249 585
R1457 vss.n4249 vss.n4248 585
R1458 vss.n5638 vss.n5637 585
R1459 vss.n5639 vss.n5638 585
R1460 vss.n5636 vss.n4238 585
R1461 vss.n4238 vss.n4237 585
R1462 vss.n5626 vss.n5625 585
R1463 vss.n5627 vss.n5626 585
R1464 vss.n4243 vss.n4242 585
R1465 vss.n5628 vss.n4243 585
R1466 vss.n5623 vss.n5622 585
R1467 vss.n5622 vss.n5621 585
R1468 vss.n4247 vss.n4246 585
R1469 vss.n5620 vss.n4247 585
R1470 vss.n5611 vss.n5610 585
R1471 vss.n5610 vss.n5609 585
R1472 vss.n5606 vss.n5605 585
R1473 vss.n5607 vss.n5606 585
R1474 vss.n5604 vss.n4255 585
R1475 vss.n4255 vss.n4254 585
R1476 vss.n5598 vss.n5597 585
R1477 vss.n5599 vss.n5598 585
R1478 vss.n5591 vss.n5590 585
R1479 vss.n5590 vss.n5589 585
R1480 vss.n4272 vss.n4271 585
R1481 vss.n5588 vss.n4272 585
R1482 vss.n4280 vss.n4278 585
R1483 vss.n4282 vss.n4280 585
R1484 vss.n4285 vss.n4281 585
R1485 vss.n5577 vss.n4281 585
R1486 vss.n5575 vss.n5574 585
R1487 vss.n5576 vss.n5575 585
R1488 vss.n4291 vss.n4290 585
R1489 vss.n5565 vss.n4291 585
R1490 vss.n4298 vss.n4297 585
R1491 vss.n5554 vss.n4298 585
R1492 vss.n5552 vss.n5551 585
R1493 vss.n5553 vss.n5552 585
R1494 vss.n4306 vss.n4303 585
R1495 vss.n4311 vss.n4306 585
R1496 vss.n4309 vss.n4308 585
R1497 vss.n4310 vss.n4309 585
R1498 vss.n4307 vss.n4304 585
R1499 vss.n5540 vss.n4307 585
R1500 vss.n5538 vss.n5537 585
R1501 vss.n5539 vss.n5538 585
R1502 vss.n4317 vss.n4316 585
R1503 vss.n5528 vss.n4317 585
R1504 vss.n5531 vss.n5530 585
R1505 vss.n5530 vss.n5529 585
R1506 vss.n4322 vss.n4319 585
R1507 vss.n4319 vss.n4318 585
R1508 vss.n4328 vss.n4325 585
R1509 vss.n4330 vss.n4328 585
R1510 vss.n5515 vss.n5514 585
R1511 vss.n5516 vss.n5515 585
R1512 vss.n4329 vss.n4326 585
R1513 vss.n5517 vss.n4329 585
R1514 vss.n5508 vss.n5507 585
R1515 vss.n5507 vss.n5506 585
R1516 vss.n4336 vss.n4335 585
R1517 vss.n5505 vss.n4336 585
R1518 vss.n4346 vss.n4344 585
R1519 vss.n4348 vss.n4346 585
R1520 vss.n4341 vss.n4338 585
R1521 vss.n4338 vss.n4337 585
R1522 vss.n4347 vss.n4345 585
R1523 vss.n5496 vss.n4347 585
R1524 vss.n5494 vss.n5493 585
R1525 vss.n5495 vss.n5494 585
R1526 vss.n4355 vss.n4353 585
R1527 vss.n4360 vss.n4355 585
R1528 vss.n4363 vss.n4356 585
R1529 vss.n5484 vss.n4356 585
R1530 vss.n5482 vss.n5481 585
R1531 vss.n5483 vss.n5482 585
R1532 vss.n4369 vss.n4368 585
R1533 vss.n5472 vss.n4369 585
R1534 vss.n4374 vss.n4371 585
R1535 vss.n4371 vss.n4370 585
R1536 vss.n4377 vss.n4375 585
R1537 vss.n4379 vss.n4377 585
R1538 vss.n5459 vss.n5458 585
R1539 vss.n5460 vss.n5459 585
R1540 vss.n5452 vss.n5451 585
R1541 vss.n5451 vss.n5450 585
R1542 vss.n4388 vss.n4387 585
R1543 vss.n5449 vss.n4388 585
R1544 vss.n4396 vss.n4394 585
R1545 vss.n4398 vss.n4396 585
R1546 vss.n4403 vss.n4400 585
R1547 vss.n4400 vss.n4399 585
R1548 vss.n4409 vss.n4406 585
R1549 vss.n4411 vss.n4409 585
R1550 vss.n5425 vss.n5424 585
R1551 vss.n5426 vss.n5425 585
R1552 vss.n4410 vss.n4407 585
R1553 vss.n5427 vss.n4410 585
R1554 vss.n5418 vss.n5417 585
R1555 vss.n5417 vss.n5416 585
R1556 vss.n4417 vss.n4416 585
R1557 vss.n5415 vss.n4417 585
R1558 vss.n4428 vss.n4425 585
R1559 vss.n4430 vss.n4428 585
R1560 vss.n4422 vss.n4419 585
R1561 vss.n4419 vss.n4418 585
R1562 vss.n4429 vss.n4426 585
R1563 vss.n5404 vss.n4429 585
R1564 vss.n5402 vss.n5401 585
R1565 vss.n5403 vss.n5402 585
R1566 vss.n4436 vss.n4435 585
R1567 vss.n5392 vss.n4436 585
R1568 vss.n5395 vss.n5394 585
R1569 vss.n5394 vss.n5393 585
R1570 vss.n4441 vss.n4438 585
R1571 vss.n4438 vss.n4437 585
R1572 vss.n4447 vss.n4444 585
R1573 vss.n4449 vss.n4447 585
R1574 vss.n5379 vss.n5378 585
R1575 vss.n5380 vss.n5379 585
R1576 vss.n4448 vss.n4445 585
R1577 vss.n5381 vss.n4448 585
R1578 vss.n4458 vss.n4452 585
R1579 vss.n4459 vss.n4458 585
R1580 vss.n4456 vss.n4454 585
R1581 vss.n4460 vss.n4456 585
R1582 vss.n5369 vss.n5368 585
R1583 vss.n5370 vss.n5369 585
R1584 vss.n5362 vss.n5361 585
R1585 vss.n5361 vss.n5360 585
R1586 vss.n4469 vss.n4468 585
R1587 vss.n5359 vss.n4469 585
R1588 vss.n4477 vss.n4475 585
R1589 vss.n4479 vss.n4477 585
R1590 vss.n4482 vss.n4478 585
R1591 vss.n5348 vss.n4478 585
R1592 vss.n5346 vss.n5345 585
R1593 vss.n5347 vss.n5346 585
R1594 vss.n4488 vss.n4487 585
R1595 vss.n5336 vss.n4488 585
R1596 vss.n4493 vss.n4490 585
R1597 vss.n4490 vss.n4489 585
R1598 vss.n4496 vss.n4494 585
R1599 vss.n4498 vss.n4496 585
R1600 vss.n5323 vss.n5322 585
R1601 vss.n5324 vss.n5323 585
R1602 vss.n4510 vss.n4507 585
R1603 vss.n5313 vss.n4510 585
R1604 vss.n5311 vss.n5310 585
R1605 vss.n5312 vss.n5311 585
R1606 vss.n4519 vss.n4516 585
R1607 vss.n4524 vss.n4519 585
R1608 vss.n4522 vss.n4521 585
R1609 vss.n4523 vss.n4522 585
R1610 vss.n4520 vss.n4517 585
R1611 vss.n5299 vss.n4520 585
R1612 vss.n5297 vss.n5296 585
R1613 vss.n5298 vss.n5297 585
R1614 vss.n4530 vss.n4529 585
R1615 vss.n5287 vss.n4530 585
R1616 vss.n5290 vss.n5289 585
R1617 vss.n5289 vss.n5288 585
R1618 vss.n4535 vss.n4532 585
R1619 vss.n4532 vss.n4531 585
R1620 vss.n4541 vss.n4538 585
R1621 vss.n4543 vss.n4541 585
R1622 vss.n5274 vss.n5273 585
R1623 vss.n5275 vss.n5274 585
R1624 vss.n4542 vss.n4539 585
R1625 vss.n5276 vss.n4542 585
R1626 vss.n5267 vss.n5266 585
R1627 vss.n5266 vss.n5265 585
R1628 vss.n4549 vss.n4548 585
R1629 vss.n5264 vss.n4549 585
R1630 vss.n4559 vss.n4557 585
R1631 vss.n4561 vss.n4559 585
R1632 vss.n4554 vss.n4551 585
R1633 vss.n4551 vss.n4550 585
R1634 vss.n4560 vss.n4558 585
R1635 vss.n5255 vss.n4560 585
R1636 vss.n5253 vss.n5252 585
R1637 vss.n5254 vss.n5253 585
R1638 vss.n4568 vss.n4566 585
R1639 vss.n4573 vss.n4568 585
R1640 vss.n4576 vss.n4569 585
R1641 vss.n5243 vss.n4569 585
R1642 vss.n5241 vss.n5240 585
R1643 vss.n5242 vss.n5241 585
R1644 vss.n4582 vss.n4581 585
R1645 vss.n5231 vss.n4582 585
R1646 vss.n4587 vss.n4584 585
R1647 vss.n4584 vss.n4583 585
R1648 vss.n4590 vss.n4588 585
R1649 vss.n4592 vss.n4590 585
R1650 vss.n5218 vss.n5217 585
R1651 vss.n5219 vss.n5218 585
R1652 vss.n5211 vss.n5210 585
R1653 vss.n5210 vss.n5209 585
R1654 vss.n4601 vss.n4600 585
R1655 vss.n5208 vss.n4601 585
R1656 vss.n4609 vss.n4607 585
R1657 vss.n4611 vss.n4609 585
R1658 vss.n4616 vss.n4613 585
R1659 vss.n4613 vss.n4612 585
R1660 vss.n4622 vss.n4619 585
R1661 vss.n4624 vss.n4622 585
R1662 vss.n5184 vss.n5183 585
R1663 vss.n5185 vss.n5184 585
R1664 vss.n4623 vss.n4620 585
R1665 vss.n5186 vss.n4623 585
R1666 vss.n5177 vss.n5176 585
R1667 vss.n5176 vss.n5175 585
R1668 vss.n4630 vss.n4629 585
R1669 vss.n5174 vss.n4630 585
R1670 vss.n4641 vss.n4638 585
R1671 vss.n4643 vss.n4641 585
R1672 vss.n4635 vss.n4632 585
R1673 vss.n4632 vss.n4631 585
R1674 vss.n4642 vss.n4639 585
R1675 vss.n5163 vss.n4642 585
R1676 vss.n5161 vss.n5160 585
R1677 vss.n5162 vss.n5161 585
R1678 vss.n4649 vss.n4648 585
R1679 vss.n5151 vss.n4649 585
R1680 vss.n5154 vss.n5153 585
R1681 vss.n5153 vss.n5152 585
R1682 vss.n4654 vss.n4651 585
R1683 vss.n4651 vss.n4650 585
R1684 vss.n4660 vss.n4657 585
R1685 vss.n4662 vss.n4660 585
R1686 vss.n5138 vss.n5137 585
R1687 vss.n5139 vss.n5138 585
R1688 vss.n4661 vss.n4658 585
R1689 vss.n5140 vss.n4661 585
R1690 vss.n4671 vss.n4665 585
R1691 vss.n4672 vss.n4671 585
R1692 vss.n4669 vss.n4667 585
R1693 vss.n4673 vss.n4669 585
R1694 vss.n5128 vss.n5127 585
R1695 vss.n5129 vss.n5128 585
R1696 vss.n5121 vss.n5120 585
R1697 vss.n5120 vss.n5119 585
R1698 vss.n4682 vss.n4681 585
R1699 vss.n5118 vss.n4682 585
R1700 vss.n4690 vss.n4688 585
R1701 vss.n4692 vss.n4690 585
R1702 vss.n4695 vss.n4691 585
R1703 vss.n5107 vss.n4691 585
R1704 vss.n5105 vss.n5104 585
R1705 vss.n5106 vss.n5105 585
R1706 vss.n4701 vss.n4700 585
R1707 vss.n5095 vss.n4701 585
R1708 vss.n4706 vss.n4703 585
R1709 vss.n4703 vss.n4702 585
R1710 vss.n4709 vss.n4707 585
R1711 vss.n4711 vss.n4709 585
R1712 vss.n5082 vss.n5081 585
R1713 vss.n5083 vss.n5082 585
R1714 vss.n4723 vss.n4720 585
R1715 vss.n5072 vss.n4723 585
R1716 vss.n5070 vss.n5069 585
R1717 vss.n5071 vss.n5070 585
R1718 vss.n4732 vss.n4729 585
R1719 vss.n4737 vss.n4732 585
R1720 vss.n4735 vss.n4734 585
R1721 vss.n4736 vss.n4735 585
R1722 vss.n4733 vss.n4730 585
R1723 vss.n5058 vss.n4733 585
R1724 vss.n5056 vss.n5055 585
R1725 vss.n5057 vss.n5056 585
R1726 vss.n4743 vss.n4742 585
R1727 vss.n5046 vss.n4743 585
R1728 vss.n5049 vss.n5048 585
R1729 vss.n5048 vss.n5047 585
R1730 vss.n4748 vss.n4745 585
R1731 vss.n4745 vss.n4744 585
R1732 vss.n4754 vss.n4751 585
R1733 vss.n4756 vss.n4754 585
R1734 vss.n5033 vss.n5032 585
R1735 vss.n5034 vss.n5033 585
R1736 vss.n4755 vss.n4752 585
R1737 vss.n5035 vss.n4755 585
R1738 vss.n5026 vss.n5025 585
R1739 vss.n5025 vss.n5024 585
R1740 vss.n4762 vss.n4761 585
R1741 vss.n5023 vss.n4762 585
R1742 vss.n4772 vss.n4770 585
R1743 vss.n4774 vss.n4772 585
R1744 vss.n4767 vss.n4764 585
R1745 vss.n4764 vss.n4763 585
R1746 vss.n4773 vss.n4771 585
R1747 vss.n5014 vss.n4773 585
R1748 vss.n5012 vss.n5011 585
R1749 vss.n5013 vss.n5012 585
R1750 vss.n4781 vss.n4779 585
R1751 vss.n4786 vss.n4781 585
R1752 vss.n4789 vss.n4782 585
R1753 vss.n5002 vss.n4782 585
R1754 vss.n5000 vss.n4999 585
R1755 vss.n5001 vss.n5000 585
R1756 vss.n4795 vss.n4794 585
R1757 vss.n4990 vss.n4795 585
R1758 vss.n4800 vss.n4797 585
R1759 vss.n4797 vss.n4796 585
R1760 vss.n4803 vss.n4801 585
R1761 vss.n4805 vss.n4803 585
R1762 vss.n4977 vss.n4976 585
R1763 vss.n4978 vss.n4977 585
R1764 vss.n4970 vss.n4969 585
R1765 vss.n4969 vss.n4968 585
R1766 vss.n4814 vss.n4813 585
R1767 vss.n4967 vss.n4814 585
R1768 vss.n4822 vss.n4820 585
R1769 vss.n4824 vss.n4822 585
R1770 vss.n4829 vss.n4826 585
R1771 vss.n4826 vss.n4825 585
R1772 vss.n4835 vss.n4832 585
R1773 vss.n4837 vss.n4835 585
R1774 vss.n4943 vss.n4942 585
R1775 vss.n4944 vss.n4943 585
R1776 vss.n4836 vss.n4833 585
R1777 vss.n4945 vss.n4836 585
R1778 vss.n4936 vss.n4935 585
R1779 vss.n4935 vss.n4934 585
R1780 vss.n4843 vss.n4842 585
R1781 vss.n4933 vss.n4843 585
R1782 vss.n4854 vss.n4851 585
R1783 vss.n4856 vss.n4854 585
R1784 vss.n4848 vss.n4845 585
R1785 vss.n4845 vss.n4844 585
R1786 vss.n4855 vss.n4852 585
R1787 vss.n4922 vss.n4855 585
R1788 vss.n4920 vss.n4919 585
R1789 vss.n4921 vss.n4920 585
R1790 vss.n4862 vss.n4861 585
R1791 vss.n4910 vss.n4862 585
R1792 vss.n4913 vss.n4912 585
R1793 vss.n4912 vss.n4911 585
R1794 vss.n4867 vss.n4864 585
R1795 vss.n4864 vss.n4863 585
R1796 vss.n4873 vss.n4870 585
R1797 vss.n4875 vss.n4873 585
R1798 vss.n4897 vss.n4896 585
R1799 vss.n4898 vss.n4897 585
R1800 vss.n4874 vss.n4871 585
R1801 vss.n4899 vss.n4874 585
R1802 vss.n4886 vss.n4878 585
R1803 vss.n4887 vss.n4886 585
R1804 vss.n4882 vss.n4880 585
R1805 vss.n4888 vss.n4882 585
R1806 vss.n4235 vss.n4234 585
R1807 vss.n6213 vss.n6201 585
R1808 vss.n6213 vss.n6206 585
R1809 vss.n4202 vss.n4197 585
R1810 vss.n4204 vss.n4202 585
R1811 vss.n6962 vss.n4205 585
R1812 vss.n6957 vss.n6956 585
R1813 vss.n6951 vss.n4208 585
R1814 vss.n6946 vss.n6945 585
R1815 vss.n6940 vss.n6939 585
R1816 vss.n6935 vss.n4213 585
R1817 vss.n6931 vss.n6930 585
R1818 vss.n4224 vss.n4221 585
R1819 vss.n6912 vss.n4225 585
R1820 vss.n6934 vss.n4185 585
R1821 vss.n6934 vss.n6933 585
R1822 vss.n6938 vss.n4212 585
R1823 vss.n6944 vss.n6943 585
R1824 vss.n6221 vss.n6220 585
R1825 vss.n6220 vss.n6219 585
R1826 vss.n6960 vss.n6959 585
R1827 vss.n6954 vss.n4207 585
R1828 vss.n6950 vss.n6949 585
R1829 vss.n6243 vss.n6242 585
R1830 vss.n6242 vss.n6241 585
R1831 vss.n6258 vss.n6257 585
R1832 vss.n6259 vss.n6258 585
R1833 vss.n6275 vss.n6274 585
R1834 vss.n6274 vss.n6273 585
R1835 vss.n6351 vss.n6350 585
R1836 vss.n6350 vss.n6349 585
R1837 vss.n6088 vss.n6085 585
R1838 vss.n6085 vss.n6084 585
R1839 vss.n6077 vss.n6070 585
R1840 vss.n6383 vss.n6070 585
R1841 vss.n6061 vss.n6059 585
R1842 vss.n6395 vss.n6061 585
R1843 vss.n5999 vss.n5995 585
R1844 vss.n6476 vss.n5995 585
R1845 vss.n6490 vss.n6489 585
R1846 vss.n6489 vss.n6488 585
R1847 vss.n6505 vss.n6504 585
R1848 vss.n6506 vss.n6505 585
R1849 vss.n6522 vss.n6521 585
R1850 vss.n6521 vss.n6520 585
R1851 vss.n6598 vss.n6597 585
R1852 vss.n6597 vss.n6596 585
R1853 vss.n5881 vss.n5878 585
R1854 vss.n5878 vss.n5877 585
R1855 vss.n5870 vss.n5863 585
R1856 vss.n6630 vss.n5863 585
R1857 vss.n5854 vss.n5852 585
R1858 vss.n6642 vss.n5854 585
R1859 vss.n5792 vss.n5788 585
R1860 vss.n6723 vss.n5788 585
R1861 vss.n6737 vss.n6736 585
R1862 vss.n6736 vss.n6735 585
R1863 vss.n6752 vss.n6751 585
R1864 vss.n6753 vss.n6752 585
R1865 vss.n6769 vss.n6768 585
R1866 vss.n6768 vss.n6767 585
R1867 vss.n6845 vss.n6844 585
R1868 vss.n6844 vss.n6843 585
R1869 vss.n5674 vss.n5671 585
R1870 vss.n5671 vss.n5670 585
R1871 vss.n5662 vss.n5659 585
R1872 vss.n6877 vss.n5659 585
R1873 vss.n6889 vss.n5647 585
R1874 vss.n5647 vss.n5646 585
R1875 vss.n6903 vss.n6902 585
R1876 vss.n6904 vss.n6903 585
R1877 vss.n4231 vss.n4227 585
R1878 vss.n6896 vss.n6895 585
R1879 vss.n6895 vss.n6894 585
R1880 vss.n5645 vss.n5644 585
R1881 vss.n6893 vss.n5645 585
R1882 vss.n6888 vss.n6887 585
R1883 vss.n6887 vss.n6886 585
R1884 vss.n6883 vss.n6882 585
R1885 vss.n6884 vss.n6883 585
R1886 vss.n6881 vss.n5651 585
R1887 vss.n5651 vss.n5650 585
R1888 vss.n6875 vss.n6874 585
R1889 vss.n6876 vss.n6875 585
R1890 vss.n6868 vss.n6867 585
R1891 vss.n6867 vss.n6866 585
R1892 vss.n5669 vss.n5668 585
R1893 vss.n6865 vss.n5669 585
R1894 vss.n5677 vss.n5675 585
R1895 vss.n5679 vss.n5677 585
R1896 vss.n5682 vss.n5678 585
R1897 vss.n6854 vss.n5678 585
R1898 vss.n6852 vss.n6851 585
R1899 vss.n6853 vss.n6852 585
R1900 vss.n5688 vss.n5687 585
R1901 vss.n6842 vss.n5688 585
R1902 vss.n5693 vss.n5690 585
R1903 vss.n5690 vss.n5689 585
R1904 vss.n5696 vss.n5694 585
R1905 vss.n5698 vss.n5696 585
R1906 vss.n5709 vss.n5706 585
R1907 vss.n5711 vss.n5709 585
R1908 vss.n5703 vss.n5700 585
R1909 vss.n5700 vss.n5699 585
R1910 vss.n5710 vss.n5707 585
R1911 vss.n6820 vss.n5710 585
R1912 vss.n6818 vss.n6817 585
R1913 vss.n6819 vss.n6818 585
R1914 vss.n5717 vss.n5716 585
R1915 vss.n6808 vss.n5717 585
R1916 vss.n6811 vss.n6810 585
R1917 vss.n6810 vss.n6809 585
R1918 vss.n5722 vss.n5719 585
R1919 vss.n5719 vss.n5718 585
R1920 vss.n5728 vss.n5725 585
R1921 vss.n5730 vss.n5728 585
R1922 vss.n6795 vss.n6794 585
R1923 vss.n6796 vss.n6795 585
R1924 vss.n5729 vss.n5726 585
R1925 vss.n6797 vss.n5729 585
R1926 vss.n6788 vss.n6787 585
R1927 vss.n6787 vss.n6786 585
R1928 vss.n5736 vss.n5735 585
R1929 vss.n6785 vss.n5736 585
R1930 vss.n5747 vss.n5744 585
R1931 vss.n5749 vss.n5747 585
R1932 vss.n5741 vss.n5738 585
R1933 vss.n5738 vss.n5737 585
R1934 vss.n5748 vss.n5745 585
R1935 vss.n6774 vss.n5748 585
R1936 vss.n6772 vss.n6771 585
R1937 vss.n6773 vss.n6772 585
R1938 vss.n5754 vss.n5753 585
R1939 vss.n6766 vss.n5754 585
R1940 vss.n6758 vss.n5756 585
R1941 vss.n5756 vss.n5755 585
R1942 vss.n6757 vss.n6756 585
R1943 vss.n6756 vss.n6755 585
R1944 vss.n6750 vss.n5762 585
R1945 vss.n5762 vss.n5761 585
R1946 vss.n5772 vss.n5769 585
R1947 vss.n6746 vss.n5769 585
R1948 vss.n6744 vss.n6743 585
R1949 vss.n6745 vss.n6744 585
R1950 vss.n5779 vss.n5778 585
R1951 vss.n6734 vss.n5779 585
R1952 vss.n5784 vss.n5781 585
R1953 vss.n5781 vss.n5780 585
R1954 vss.n5787 vss.n5785 585
R1955 vss.n5789 vss.n5787 585
R1956 vss.n6721 vss.n6720 585
R1957 vss.n6722 vss.n6721 585
R1958 vss.n6714 vss.n6713 585
R1959 vss.n6713 vss.n6712 585
R1960 vss.n5798 vss.n5797 585
R1961 vss.n6711 vss.n5798 585
R1962 vss.n6698 vss.n6697 585
R1963 vss.n6699 vss.n6698 585
R1964 vss.n5805 vss.n5804 585
R1965 vss.n6700 vss.n5805 585
R1966 vss.n5816 vss.n5815 585
R1967 vss.n5817 vss.n5816 585
R1968 vss.n5813 vss.n5810 585
R1969 vss.n5818 vss.n5813 585
R1970 vss.n6684 vss.n6683 585
R1971 vss.n6685 vss.n6684 585
R1972 vss.n5814 vss.n5811 585
R1973 vss.n6686 vss.n5814 585
R1974 vss.n6677 vss.n6676 585
R1975 vss.n6676 vss.n6675 585
R1976 vss.n5824 vss.n5823 585
R1977 vss.n6674 vss.n5824 585
R1978 vss.n5835 vss.n5832 585
R1979 vss.n5837 vss.n5835 585
R1980 vss.n5829 vss.n5826 585
R1981 vss.n5826 vss.n5825 585
R1982 vss.n5836 vss.n5833 585
R1983 vss.n6663 vss.n5836 585
R1984 vss.n6661 vss.n6660 585
R1985 vss.n6662 vss.n6661 585
R1986 vss.n5843 vss.n5842 585
R1987 vss.n6651 vss.n5843 585
R1988 vss.n6654 vss.n6653 585
R1989 vss.n6653 vss.n6652 585
R1990 vss.n5848 vss.n5845 585
R1991 vss.n5845 vss.n5844 585
R1992 vss.n5853 vss.n5851 585
R1993 vss.n5855 vss.n5853 585
R1994 vss.n6640 vss.n6639 585
R1995 vss.n6641 vss.n6640 585
R1996 vss.n5865 vss.n5864 585
R1997 vss.n5866 vss.n5865 585
R1998 vss.n5862 vss.n5860 585
R1999 vss.n5867 vss.n5862 585
R2000 vss.n6628 vss.n6627 585
R2001 vss.n6629 vss.n6628 585
R2002 vss.n6621 vss.n6620 585
R2003 vss.n6620 vss.n6619 585
R2004 vss.n5876 vss.n5875 585
R2005 vss.n6618 vss.n5876 585
R2006 vss.n5884 vss.n5882 585
R2007 vss.n5886 vss.n5884 585
R2008 vss.n5889 vss.n5885 585
R2009 vss.n6607 vss.n5885 585
R2010 vss.n6605 vss.n6604 585
R2011 vss.n6606 vss.n6605 585
R2012 vss.n5895 vss.n5894 585
R2013 vss.n6595 vss.n5895 585
R2014 vss.n5900 vss.n5897 585
R2015 vss.n5897 vss.n5896 585
R2016 vss.n5903 vss.n5901 585
R2017 vss.n5905 vss.n5903 585
R2018 vss.n5916 vss.n5913 585
R2019 vss.n5918 vss.n5916 585
R2020 vss.n5910 vss.n5907 585
R2021 vss.n5907 vss.n5906 585
R2022 vss.n5917 vss.n5914 585
R2023 vss.n6573 vss.n5917 585
R2024 vss.n6571 vss.n6570 585
R2025 vss.n6572 vss.n6571 585
R2026 vss.n5924 vss.n5923 585
R2027 vss.n6561 vss.n5924 585
R2028 vss.n6564 vss.n6563 585
R2029 vss.n6563 vss.n6562 585
R2030 vss.n5929 vss.n5926 585
R2031 vss.n5926 vss.n5925 585
R2032 vss.n5935 vss.n5932 585
R2033 vss.n5937 vss.n5935 585
R2034 vss.n6548 vss.n6547 585
R2035 vss.n6549 vss.n6548 585
R2036 vss.n5936 vss.n5933 585
R2037 vss.n6550 vss.n5936 585
R2038 vss.n6541 vss.n6540 585
R2039 vss.n6540 vss.n6539 585
R2040 vss.n5943 vss.n5942 585
R2041 vss.n6538 vss.n5943 585
R2042 vss.n5954 vss.n5951 585
R2043 vss.n5956 vss.n5954 585
R2044 vss.n5948 vss.n5945 585
R2045 vss.n5945 vss.n5944 585
R2046 vss.n5955 vss.n5952 585
R2047 vss.n6527 vss.n5955 585
R2048 vss.n6525 vss.n6524 585
R2049 vss.n6526 vss.n6525 585
R2050 vss.n5961 vss.n5960 585
R2051 vss.n6519 vss.n5961 585
R2052 vss.n6511 vss.n5963 585
R2053 vss.n5963 vss.n5962 585
R2054 vss.n6510 vss.n6509 585
R2055 vss.n6509 vss.n6508 585
R2056 vss.n6503 vss.n5969 585
R2057 vss.n5969 vss.n5968 585
R2058 vss.n5979 vss.n5976 585
R2059 vss.n6499 vss.n5976 585
R2060 vss.n6497 vss.n6496 585
R2061 vss.n6498 vss.n6497 585
R2062 vss.n5986 vss.n5985 585
R2063 vss.n6487 vss.n5986 585
R2064 vss.n5991 vss.n5988 585
R2065 vss.n5988 vss.n5987 585
R2066 vss.n5994 vss.n5992 585
R2067 vss.n5996 vss.n5994 585
R2068 vss.n6474 vss.n6473 585
R2069 vss.n6475 vss.n6474 585
R2070 vss.n6467 vss.n6466 585
R2071 vss.n6466 vss.n6465 585
R2072 vss.n6005 vss.n6004 585
R2073 vss.n6464 vss.n6005 585
R2074 vss.n6451 vss.n6450 585
R2075 vss.n6452 vss.n6451 585
R2076 vss.n6011 vss.n6010 585
R2077 vss.n6453 vss.n6011 585
R2078 vss.n6023 vss.n6022 585
R2079 vss.n6024 vss.n6023 585
R2080 vss.n6020 vss.n6017 585
R2081 vss.n6025 vss.n6020 585
R2082 vss.n6437 vss.n6436 585
R2083 vss.n6438 vss.n6437 585
R2084 vss.n6021 vss.n6018 585
R2085 vss.n6439 vss.n6021 585
R2086 vss.n6430 vss.n6429 585
R2087 vss.n6429 vss.n6428 585
R2088 vss.n6031 vss.n6030 585
R2089 vss.n6427 vss.n6031 585
R2090 vss.n6042 vss.n6039 585
R2091 vss.n6044 vss.n6042 585
R2092 vss.n6036 vss.n6033 585
R2093 vss.n6033 vss.n6032 585
R2094 vss.n6043 vss.n6040 585
R2095 vss.n6416 vss.n6043 585
R2096 vss.n6414 vss.n6413 585
R2097 vss.n6415 vss.n6414 585
R2098 vss.n6050 vss.n6049 585
R2099 vss.n6404 vss.n6050 585
R2100 vss.n6407 vss.n6406 585
R2101 vss.n6406 vss.n6405 585
R2102 vss.n6055 vss.n6052 585
R2103 vss.n6052 vss.n6051 585
R2104 vss.n6060 vss.n6058 585
R2105 vss.n6062 vss.n6060 585
R2106 vss.n6393 vss.n6392 585
R2107 vss.n6394 vss.n6393 585
R2108 vss.n6072 vss.n6071 585
R2109 vss.n6073 vss.n6072 585
R2110 vss.n6069 vss.n6067 585
R2111 vss.n6074 vss.n6069 585
R2112 vss.n6381 vss.n6380 585
R2113 vss.n6382 vss.n6381 585
R2114 vss.n6374 vss.n6373 585
R2115 vss.n6373 vss.n6372 585
R2116 vss.n6083 vss.n6082 585
R2117 vss.n6371 vss.n6083 585
R2118 vss.n6091 vss.n6089 585
R2119 vss.n6093 vss.n6091 585
R2120 vss.n6096 vss.n6092 585
R2121 vss.n6360 vss.n6092 585
R2122 vss.n6358 vss.n6357 585
R2123 vss.n6359 vss.n6358 585
R2124 vss.n6102 vss.n6101 585
R2125 vss.n6348 vss.n6102 585
R2126 vss.n6107 vss.n6104 585
R2127 vss.n6104 vss.n6103 585
R2128 vss.n6110 vss.n6108 585
R2129 vss.n6112 vss.n6110 585
R2130 vss.n6123 vss.n6120 585
R2131 vss.n6125 vss.n6123 585
R2132 vss.n6117 vss.n6114 585
R2133 vss.n6114 vss.n6113 585
R2134 vss.n6124 vss.n6121 585
R2135 vss.n6326 vss.n6124 585
R2136 vss.n6324 vss.n6323 585
R2137 vss.n6325 vss.n6324 585
R2138 vss.n6131 vss.n6130 585
R2139 vss.n6314 vss.n6131 585
R2140 vss.n6317 vss.n6316 585
R2141 vss.n6316 vss.n6315 585
R2142 vss.n6136 vss.n6133 585
R2143 vss.n6133 vss.n6132 585
R2144 vss.n6142 vss.n6139 585
R2145 vss.n6144 vss.n6142 585
R2146 vss.n6301 vss.n6300 585
R2147 vss.n6302 vss.n6301 585
R2148 vss.n6143 vss.n6140 585
R2149 vss.n6303 vss.n6143 585
R2150 vss.n6294 vss.n6293 585
R2151 vss.n6293 vss.n6292 585
R2152 vss.n6150 vss.n6149 585
R2153 vss.n6291 vss.n6150 585
R2154 vss.n6161 vss.n6158 585
R2155 vss.n6163 vss.n6161 585
R2156 vss.n6155 vss.n6152 585
R2157 vss.n6152 vss.n6151 585
R2158 vss.n6162 vss.n6159 585
R2159 vss.n6280 vss.n6162 585
R2160 vss.n6278 vss.n6277 585
R2161 vss.n6279 vss.n6278 585
R2162 vss.n6168 vss.n6167 585
R2163 vss.n6272 vss.n6168 585
R2164 vss.n6264 vss.n6170 585
R2165 vss.n6170 vss.n6169 585
R2166 vss.n6263 vss.n6262 585
R2167 vss.n6262 vss.n6261 585
R2168 vss.n6256 vss.n6176 585
R2169 vss.n6176 vss.n6175 585
R2170 vss.n6186 vss.n6183 585
R2171 vss.n6252 vss.n6183 585
R2172 vss.n6250 vss.n6249 585
R2173 vss.n6251 vss.n6250 585
R2174 vss.n6193 vss.n6192 585
R2175 vss.n6240 vss.n6193 585
R2176 vss.n6207 vss.n6195 585
R2177 vss.n6195 vss.n6194 585
R2178 vss.n6209 vss.n6208 585
R2179 vss.n6210 vss.n6209 585
R2180 vss.n6216 vss.n6215 585
R2181 vss.n6217 vss.n6216 585
R2182 vss.n6909 vss.n4226 585
R2183 vss.n6908 vss.n6907 585
R2184 vss.n6920 vss.n6919 585
R2185 vss.n6924 vss.n6923 585
R2186 vss.n6923 vss.n6922 585
R2187 vss.n6929 vss.n4216 585
R2188 vss.n7020 vss.n4157 585
R2189 vss.n12171 vss.n12170 562.79
R2190 vss.n11989 vss.n11988 562.79
R2191 vss.n11323 vss.n11322 562.79
R2192 vss.n14311 vss.n14310 562.79
R2193 vss.n11611 vss.n11610 562.79
R2194 vss.n11824 vss.n11823 562.79
R2195 vss.n14801 vss.n14800 562.79
R2196 vss.n14628 vss.n14627 562.79
R2197 vss.n14539 vss.n14538 562.79
R2198 vss.n14260 vss.n14259 562.79
R2199 vss.n14892 vss.n14891 562.79
R2200 vss.n15054 vss.n15053 562.79
R2201 vss.n12704 vss.n12703 562.79
R2202 vss.n16898 vss.n16897 492.105
R2203 vss.n17134 vss.n17133 492.105
R2204 vss.n15943 vss.n15942 492.105
R2205 vss.n16179 vss.n16178 492.105
R2206 vss.n15419 vss.n15418 492.105
R2207 vss.n15655 vss.n15654 492.105
R2208 vss.n16366 vss.n16365 492.105
R2209 vss.n16602 vss.n16601 492.105
R2210 vss.n20222 vss.n19088 463.157
R2211 vss.n20220 vss.n19089 463.157
R2212 vss.n20101 vss.n20100 463.157
R2213 vss.n20091 vss.n20090 463.157
R2214 vss.n19975 vss.n19295 463.157
R2215 vss.n19973 vss.n19296 463.157
R2216 vss.n19854 vss.n19853 463.157
R2217 vss.n19844 vss.n19843 463.157
R2218 vss.n19728 vss.n19502 463.157
R2219 vss.n19726 vss.n19503 463.157
R2220 vss.n20356 vss.n17594 463.157
R2221 vss.n20354 vss.n17595 463.157
R2222 vss.n18955 vss.n18954 463.157
R2223 vss.n18945 vss.n18944 463.157
R2224 vss.n18829 vss.n17788 463.157
R2225 vss.n18827 vss.n17789 463.157
R2226 vss.n18714 vss.n17889 463.157
R2227 vss.n18704 vss.n18703 463.157
R2228 vss.n18588 vss.n18001 463.157
R2229 vss.n18586 vss.n18002 463.157
R2230 vss.n18473 vss.n18102 463.157
R2231 vss.n18463 vss.n18462 463.157
R2232 vss.n18347 vss.n18214 463.157
R2233 vss.n18345 vss.n18215 463.157
R2234 vss.n6832 vss.n5698 463.157
R2235 vss.n6830 vss.n5699 463.157
R2236 vss.n6711 vss.n6710 463.157
R2237 vss.n6701 vss.n6700 463.157
R2238 vss.n6585 vss.n5905 463.157
R2239 vss.n6583 vss.n5906 463.157
R2240 vss.n6464 vss.n6463 463.157
R2241 vss.n6454 vss.n6453 463.157
R2242 vss.n6338 vss.n6112 463.157
R2243 vss.n6336 vss.n6113 463.157
R2244 vss.n6966 vss.n4204 463.157
R2245 vss.n6964 vss.n4205 463.157
R2246 vss.n5565 vss.n5564 463.157
R2247 vss.n5555 vss.n5554 463.157
R2248 vss.n5439 vss.n4398 463.157
R2249 vss.n5437 vss.n4399 463.157
R2250 vss.n5324 vss.n4499 463.157
R2251 vss.n5314 vss.n5313 463.157
R2252 vss.n5198 vss.n4611 463.157
R2253 vss.n5196 vss.n4612 463.157
R2254 vss.n5083 vss.n4712 463.157
R2255 vss.n5073 vss.n5072 463.157
R2256 vss.n4957 vss.n4824 463.157
R2257 vss.n4955 vss.n4825 463.157
R2258 vss.n16775 vss.n16774 463.157
R2259 vss.n16793 vss.n16792 463.157
R2260 vss.n17007 vss.n17006 463.157
R2261 vss.n17024 vss.n17023 463.157
R2262 vss.n17243 vss.n17242 463.157
R2263 vss.n17262 vss.n17261 463.157
R2264 vss.n15236 vss.n15235 463.157
R2265 vss.n15319 vss.n15318 463.157
R2266 vss.n15527 vss.n15526 463.157
R2267 vss.n15544 vss.n15543 463.157
R2268 vss.n15763 vss.n15762 463.157
R2269 vss.n15778 vss.n15777 463.157
R2270 vss.n16474 vss.n16473 463.157
R2271 vss.n16491 vss.n16490 463.157
R2272 vss.n12185 vss.n12184 460.465
R2273 vss.n10855 vss.n10854 460.465
R2274 vss.n11298 vss.n11297 460.465
R2275 vss.n11159 vss.n11158 460.465
R2276 vss.n14297 vss.n14296 460.465
R2277 vss.n14010 vss.n14009 460.465
R2278 vss.n11799 vss.n11798 460.465
R2279 vss.n11083 vss.n11082 460.465
R2280 vss.n14787 vss.n14786 460.465
R2281 vss.n13531 vss.n13530 460.465
R2282 vss.n14522 vss.n14521 460.465
R2283 vss.n14240 vss.n14239 460.465
R2284 vss.n14877 vss.n14876 460.465
R2285 vss.n12807 vss.n12806 460.465
R2286 vss.n12688 vss.n12687 460.465
R2287 vss.n12551 vss.n12550 460.465
R2288 vss.n17337 vss.n17336 457.142
R2289 vss.n17348 vss.n17347 457.142
R2290 vss.n17359 vss.n17358 457.142
R2291 vss.n17370 vss.n17369 457.142
R2292 vss.n17381 vss.n17380 457.142
R2293 vss.n17392 vss.n17391 457.142
R2294 vss.n17414 vss.n17413 457.142
R2295 vss.n17425 vss.n17424 457.142
R2296 vss.n17436 vss.n17435 457.142
R2297 vss.n17447 vss.n17446 457.142
R2298 vss.n17458 vss.n17457 457.142
R2299 vss.n17469 vss.n17468 457.142
R2300 vss.n17480 vss.n17479 457.142
R2301 vss.n3495 vss.n3494 457.142
R2302 vss.n3506 vss.n3505 457.142
R2303 vss.n3517 vss.n3516 457.142
R2304 vss.n3528 vss.n3527 457.142
R2305 vss.n3539 vss.n3538 457.142
R2306 vss.n3550 vss.n3549 457.142
R2307 vss.n4024 vss.n4023 457.142
R2308 vss.n4035 vss.n4034 457.142
R2309 vss.n4046 vss.n4045 457.142
R2310 vss.n4057 vss.n4056 457.142
R2311 vss.n4068 vss.n4067 457.142
R2312 vss.n4079 vss.n4078 457.142
R2313 vss.n4090 vss.n4089 457.142
R2314 vss.n20284 vss.n20283 434.21
R2315 vss.n20276 vss.n19036 434.21
R2316 vss.n20164 vss.n20163 434.21
R2317 vss.n20157 vss.n20156 434.21
R2318 vss.n19245 vss.n19234 434.21
R2319 vss.n20032 vss.n20031 434.21
R2320 vss.n19917 vss.n19916 434.21
R2321 vss.n19910 vss.n19909 434.21
R2322 vss.n19452 vss.n19441 434.21
R2323 vss.n19785 vss.n19784 434.21
R2324 vss.n19670 vss.n19669 434.21
R2325 vss.n19663 vss.n19662 434.21
R2326 vss.n20312 vss.n17614 434.21
R2327 vss.n20310 vss.n17615 434.21
R2328 vss.n19018 vss.n19017 434.21
R2329 vss.n19011 vss.n19010 434.21
R2330 vss.n17738 vss.n17727 434.21
R2331 vss.n18886 vss.n18885 434.21
R2332 vss.n18771 vss.n18770 434.21
R2333 vss.n17850 vss.n17849 434.21
R2334 vss.n17951 vss.n17940 434.21
R2335 vss.n18645 vss.n18644 434.21
R2336 vss.n18530 vss.n18529 434.21
R2337 vss.n18063 vss.n18062 434.21
R2338 vss.n18164 vss.n18153 434.21
R2339 vss.n18404 vss.n18403 434.21
R2340 vss.n18289 vss.n18288 434.21
R2341 vss.n18278 vss.n18277 434.21
R2342 vss.n6894 vss.n6893 434.21
R2343 vss.n6886 vss.n5646 434.21
R2344 vss.n6774 vss.n6773 434.21
R2345 vss.n6767 vss.n6766 434.21
R2346 vss.n5855 vss.n5844 434.21
R2347 vss.n6642 vss.n6641 434.21
R2348 vss.n6527 vss.n6526 434.21
R2349 vss.n6520 vss.n6519 434.21
R2350 vss.n6062 vss.n6051 434.21
R2351 vss.n6395 vss.n6394 434.21
R2352 vss.n6280 vss.n6279 434.21
R2353 vss.n6273 vss.n6272 434.21
R2354 vss.n6922 vss.n4224 434.21
R2355 vss.n6920 vss.n4225 434.21
R2356 vss.n5628 vss.n5627 434.21
R2357 vss.n5621 vss.n5620 434.21
R2358 vss.n4348 vss.n4337 434.21
R2359 vss.n5496 vss.n5495 434.21
R2360 vss.n5381 vss.n5380 434.21
R2361 vss.n4460 vss.n4459 434.21
R2362 vss.n4561 vss.n4550 434.21
R2363 vss.n5255 vss.n5254 434.21
R2364 vss.n5140 vss.n5139 434.21
R2365 vss.n4673 vss.n4672 434.21
R2366 vss.n4774 vss.n4763 434.21
R2367 vss.n5014 vss.n5013 434.21
R2368 vss.n4899 vss.n4898 434.21
R2369 vss.n4888 vss.n4887 434.21
R2370 vss.n16885 vss.n16884 434.21
R2371 vss.n16908 vss.n16907 434.21
R2372 vss.n17121 vss.n17120 434.21
R2373 vss.n17144 vss.n17143 434.21
R2374 vss.n15931 vss.n15930 434.21
R2375 vss.n15955 vss.n15954 434.21
R2376 vss.n16167 vss.n16166 434.21
R2377 vss.n16191 vss.n16190 434.21
R2378 vss.n16247 vss.n16246 434.21
R2379 vss.n15407 vss.n15406 434.21
R2380 vss.n15428 vss.n15427 434.21
R2381 vss.n15643 vss.n15642 434.21
R2382 vss.n15664 vss.n15663 434.21
R2383 vss.n16354 vss.n16353 434.21
R2384 vss.n16375 vss.n16374 434.21
R2385 vss.n16590 vss.n16589 434.21
R2386 vss.n16611 vss.n16610 434.21
R2387 vss.n16670 vss.n16669 434.21
R2388 vss.n14275 vss.n14274 431.372
R2389 vss.n11040 vss.n11039 431.372
R2390 vss.n12526 vss.n12525 431.372
R2391 vss.n13226 vss.n13225 431.372
R2392 vss.n20232 vss.n20231 405.263
R2393 vss.n20211 vss.n20210 405.263
R2394 vss.n20112 vss.n19180 405.263
R2395 vss.n19207 vss.n19196 405.263
R2396 vss.n19985 vss.n19984 405.263
R2397 vss.n19964 vss.n19963 405.263
R2398 vss.n19865 vss.n19387 405.263
R2399 vss.n19414 vss.n19403 405.263
R2400 vss.n19738 vss.n19737 405.263
R2401 vss.n19717 vss.n19716 405.263
R2402 vss.n19608 vss.n19607 405.263
R2403 vss.n20348 vss.n20347 405.263
R2404 vss.n18966 vss.n17673 405.263
R2405 vss.n17700 vss.n17689 405.263
R2406 vss.n18839 vss.n18838 405.263
R2407 vss.n18818 vss.n18817 405.263
R2408 vss.n18716 vss.n17888 405.263
R2409 vss.n17913 vss.n17902 405.263
R2410 vss.n18598 vss.n18597 405.263
R2411 vss.n18577 vss.n18576 405.263
R2412 vss.n18475 vss.n18101 405.263
R2413 vss.n18126 vss.n18115 405.263
R2414 vss.n18357 vss.n18356 405.263
R2415 vss.n18336 vss.n18335 405.263
R2416 vss.n6842 vss.n6841 405.263
R2417 vss.n6821 vss.n6820 405.263
R2418 vss.n6722 vss.n5790 405.263
R2419 vss.n5817 vss.n5806 405.263
R2420 vss.n6595 vss.n6594 405.263
R2421 vss.n6574 vss.n6573 405.263
R2422 vss.n6475 vss.n5997 405.263
R2423 vss.n6024 vss.n6013 405.263
R2424 vss.n6348 vss.n6347 405.263
R2425 vss.n6327 vss.n6326 405.263
R2426 vss.n6218 vss.n6217 405.263
R2427 vss.n6958 vss.n6957 405.263
R2428 vss.n5576 vss.n4283 405.263
R2429 vss.n4310 vss.n4299 405.263
R2430 vss.n5449 vss.n5448 405.263
R2431 vss.n5428 vss.n5427 405.263
R2432 vss.n5326 vss.n4498 405.263
R2433 vss.n4523 vss.n4512 405.263
R2434 vss.n5208 vss.n5207 405.263
R2435 vss.n5187 vss.n5186 405.263
R2436 vss.n5085 vss.n4711 405.263
R2437 vss.n4736 vss.n4725 405.263
R2438 vss.n4967 vss.n4966 405.263
R2439 vss.n4946 vss.n4945 405.263
R2440 vss.n16763 vss.n16762 405.263
R2441 vss.n16804 vss.n16803 405.263
R2442 vss.n16993 vss.n16992 405.263
R2443 vss.n17038 vss.n17037 405.263
R2444 vss.n17229 vss.n17228 405.263
R2445 vss.n17293 vss.n17292 405.263
R2446 vss.n15246 vss.n15245 405.263
R2447 vss.n15224 vss.n15223 405.263
R2448 vss.n15513 vss.n15512 405.263
R2449 vss.n15560 vss.n15559 405.263
R2450 vss.n15749 vss.n15748 405.263
R2451 vss.n15790 vss.n15789 405.263
R2452 vss.n16460 vss.n16459 405.263
R2453 vss.n16507 vss.n16506 405.263
R2454 vss.n22599 vss.n22598 400
R2455 vss.n22580 vss.n22579 400
R2456 vss.n22391 vss.n22390 400
R2457 vss.n22372 vss.n22371 400
R2458 vss.n22183 vss.n22182 400
R2459 vss.n22164 vss.n22163 400
R2460 vss.n21527 vss.n21526 400
R2461 vss.n21508 vss.n21507 400
R2462 vss.n21319 vss.n21318 400
R2463 vss.n21300 vss.n21299 400
R2464 vss.n21111 vss.n21110 400
R2465 vss.n21092 vss.n21091 400
R2466 vss.n20903 vss.n20902 400
R2467 vss.n8762 vss.n8761 400
R2468 vss.n8743 vss.n8742 400
R2469 vss.n8554 vss.n8553 400
R2470 vss.n8535 vss.n8534 400
R2471 vss.n8346 vss.n8345 400
R2472 vss.n8327 vss.n8326 400
R2473 vss.n8138 vss.n8137 400
R2474 vss.n8119 vss.n8118 400
R2475 vss.n7930 vss.n7929 400
R2476 vss.n7911 vss.n7910 400
R2477 vss.n7721 vss.n7720 400
R2478 vss.n7702 vss.n7701 400
R2479 vss.n7513 vss.n7512 400
R2480 vss.n9653 vss.n9651 394
R2481 vss.n10218 vss.n10216 394
R2482 vss.n1 vss.n20294 339.711
R2483 vss.n20274 vss.n19040 376.315
R2484 vss.n19139 vss.n19127 376.315
R2485 vss.n20145 vss.n19145 376.315
R2486 vss.n20042 vss.n20041 376.315
R2487 vss.n19257 vss.n19256 376.315
R2488 vss.n19346 vss.n19334 376.315
R2489 vss.n19898 vss.n19352 376.315
R2490 vss.n19795 vss.n19794 376.315
R2491 vss.n19464 vss.n19463 376.315
R2492 vss.n19553 vss.n19541 376.315
R2493 vss.n19651 vss.n19559 376.315
R2494 vss.n20321 vss.n17606 376.315
R2495 vss.n20299 vss.n20298 376.315
R2496 vss.n19029 vss.n17627 376.315
R2497 vss.n18999 vss.n17638 376.315
R2498 vss.n18896 vss.n18895 376.315
R2499 vss.n17750 vss.n17749 376.315
R2500 vss.n17839 vss.n17827 376.315
R2501 vss.n18761 vss.n18760 376.315
R2502 vss.n18655 vss.n18654 376.315
R2503 vss.n17963 vss.n17962 376.315
R2504 vss.n18052 vss.n18040 376.315
R2505 vss.n18520 vss.n18519 376.315
R2506 vss.n18414 vss.n18413 376.315
R2507 vss.n18176 vss.n18175 376.315
R2508 vss.n18265 vss.n18253 376.315
R2509 vss.n18279 vss.n3 339.711
R2510 vss.n5 vss.n6904 339.711
R2511 vss.n6884 vss.n5650 376.315
R2512 vss.n5749 vss.n5737 376.315
R2513 vss.n6755 vss.n5755 376.315
R2514 vss.n6652 vss.n6651 376.315
R2515 vss.n5867 vss.n5866 376.315
R2516 vss.n5956 vss.n5944 376.315
R2517 vss.n6508 vss.n5962 376.315
R2518 vss.n6405 vss.n6404 376.315
R2519 vss.n6074 vss.n6073 376.315
R2520 vss.n6163 vss.n6151 376.315
R2521 vss.n6261 vss.n6169 376.315
R2522 vss.n6931 vss.n4216 376.315
R2523 vss.n6909 vss.n6908 376.315
R2524 vss.n5639 vss.n4237 376.315
R2525 vss.n5609 vss.n4248 376.315
R2526 vss.n5506 vss.n5505 376.315
R2527 vss.n4360 vss.n4359 376.315
R2528 vss.n4449 vss.n4437 376.315
R2529 vss.n5371 vss.n5370 376.315
R2530 vss.n5265 vss.n5264 376.315
R2531 vss.n4573 vss.n4572 376.315
R2532 vss.n4662 vss.n4650 376.315
R2533 vss.n5130 vss.n5129 376.315
R2534 vss.n5024 vss.n5023 376.315
R2535 vss.n4786 vss.n4785 376.315
R2536 vss.n4875 vss.n4863 376.315
R2537 vss.n4889 vss.n7 339.711
R2538 vss.n16692 vss.n16691 376.315
R2539 vss.n16871 vss.n16870 376.315
R2540 vss.n16922 vss.n16921 376.315
R2541 vss.n17107 vss.n17106 376.315
R2542 vss.n17158 vss.n17157 376.315
R2543 vss.n17269 vss.n17268 376.315
R2544 vss.n15917 vss.n15916 376.315
R2545 vss.n15969 vss.n15968 376.315
R2546 vss.n16153 vss.n16152 376.315
R2547 vss.n16205 vss.n16204 376.315
R2548 vss.n16278 vss.n16277 376.315
R2549 vss.n15393 vss.n15392 376.315
R2550 vss.n15442 vss.n15441 376.315
R2551 vss.n15629 vss.n15628 376.315
R2552 vss.n15678 vss.n15677 376.315
R2553 vss.n15857 vss.n15856 376.315
R2554 vss.n16340 vss.n16339 376.315
R2555 vss.n16389 vss.n16388 376.315
R2556 vss.n16576 vss.n16575 376.315
R2557 vss.n16625 vss.n16624 376.315
R2558 vss.n14357 vss.n14356 373.856
R2559 vss.n13863 vss.n13862 373.856
R2560 vss.n14491 vss.n14490 373.856
R2561 vss.n14398 vss.n14397 373.856
R2562 vss.n13978 vss.n13977 373.856
R2563 vss.n11573 vss.n11572 373.856
R2564 vss.n11760 vss.n11759 373.856
R2565 vss.n11050 vss.n11049 373.856
R2566 vss.n12425 vss.n12424 373.856
R2567 vss.n12598 vss.n12597 373.856
R2568 vss.n12583 vss.n12582 373.856
R2569 vss.n12079 vss.n12078 373.856
R2570 vss.n14661 vss.n14660 373.856
R2571 vss.n13580 vss.n13579 373.856
R2572 vss.n15015 vss.n15014 373.856
R2573 vss.n10506 vss.n10505 373.856
R2574 vss.n13298 vss.n13297 373.856
R2575 vss.n13339 vss.n13338 373.856
R2576 vss.n13240 vss.n13239 373.856
R2577 vss.n14961 vss.n14960 373.856
R2578 vss.n10824 vss.n10823 373.856
R2579 vss.n10898 vss.n10897 373.856
R2580 vss.n10951 vss.n10950 373.856
R2581 vss.n11011 vss.n11010 373.856
R2582 vss.n20531 vss.n20530 367.823
R2583 vss.n20558 vss.n20553 367.823
R2584 vss.n20760 vss.n20759 367.823
R2585 vss.n20780 vss.n20775 367.823
R2586 vss.n7141 vss.n7140 367.823
R2587 vss.n7168 vss.n7163 367.823
R2588 vss.n7370 vss.n7369 367.823
R2589 vss.n7390 vss.n7385 367.823
R2590 vss.n1757 vss.n1756 367.823
R2591 vss.n1777 vss.n1772 367.823
R2592 vss.n1988 vss.n1987 367.823
R2593 vss.n2017 vss.n2010 367.823
R2594 vss.n2233 vss.n2232 367.823
R2595 vss.n2261 vss.n2254 367.823
R2596 vss.n2477 vss.n2476 367.823
R2597 vss.n2505 vss.n2498 367.823
R2598 vss.n2722 vss.n2721 367.823
R2599 vss.n2750 vss.n2743 367.823
R2600 vss.n2960 vss.n2959 367.823
R2601 vss.n2988 vss.n2981 367.823
R2602 vss.n3204 vss.n3203 367.823
R2603 vss.n3233 vss.n3226 367.823
R2604 vss.n15206 vss.n15205 367.823
R2605 vss.n15186 vss.n15181 367.823
R2606 vss.n218 vss.n217 367.823
R2607 vss.n238 vss.n233 367.823
R2608 vss.n449 vss.n448 367.823
R2609 vss.n478 vss.n471 367.823
R2610 vss.n694 vss.n693 367.823
R2611 vss.n722 vss.n715 367.823
R2612 vss.n938 vss.n937 367.823
R2613 vss.n966 vss.n959 367.823
R2614 vss.n1183 vss.n1182 367.823
R2615 vss.n1211 vss.n1204 367.823
R2616 vss.n23306 vss.n23305 367.823
R2617 vss.n23278 vss.n23271 367.823
R2618 vss.n23062 vss.n23061 367.823
R2619 vss.n23033 vss.n23026 367.823
R2620 vss.n1399 vss.n1398 367.823
R2621 vss.n22820 vss.n22815 367.823
R2622 vss.n12199 vss.n12198 358.139
R2623 vss.n12003 vss.n12002 358.139
R2624 vss.n11282 vss.n11281 358.139
R2625 vss.n11180 vss.n11179 358.139
R2626 vss.n13879 vss.n13878 358.139
R2627 vss.n13989 vss.n13988 358.139
R2628 vss.n11783 vss.n11782 358.139
R2629 vss.n11093 vss.n11092 358.139
R2630 vss.n14773 vss.n14772 358.139
R2631 vss.n13514 vss.n13513 358.139
R2632 vss.n14506 vss.n14505 358.139
R2633 vss.n14220 vss.n14219 358.139
R2634 vss.n12840 vss.n12839 358.139
R2635 vss.n12813 vss.n12812 358.139
R2636 vss.n12671 vss.n12670 358.139
R2637 vss.n12557 vss.n12556 358.139
R2638 vss.n20243 vss.n19070 347.368
R2639 vss.n20199 vss.n19102 347.368
R2640 vss.n20114 vss.n19179 347.368
R2641 vss.n20077 vss.n20076 347.368
R2642 vss.n19996 vss.n19277 347.368
R2643 vss.n19952 vss.n19309 347.368
R2644 vss.n19867 vss.n19386 347.368
R2645 vss.n19830 vss.n19829 347.368
R2646 vss.n19749 vss.n19484 347.368
R2647 vss.n19705 vss.n19516 347.368
R2648 vss.n19601 vss.n19600 347.368
R2649 vss.n20342 vss.n20341 347.368
R2650 vss.n18968 vss.n17672 347.368
R2651 vss.n18931 vss.n18930 347.368
R2652 vss.n18850 vss.n17770 347.368
R2653 vss.n18806 vss.n17802 347.368
R2654 vss.n18726 vss.n18725 347.368
R2655 vss.n18690 vss.n18689 347.368
R2656 vss.n18609 vss.n17983 347.368
R2657 vss.n18565 vss.n18015 347.368
R2658 vss.n18485 vss.n18484 347.368
R2659 vss.n18449 vss.n18448 347.368
R2660 vss.n18368 vss.n18196 347.368
R2661 vss.n18324 vss.n18228 347.368
R2662 vss.n6853 vss.n5680 347.368
R2663 vss.n6809 vss.n5712 347.368
R2664 vss.n6724 vss.n5789 347.368
R2665 vss.n6687 vss.n6686 347.368
R2666 vss.n6606 vss.n5887 347.368
R2667 vss.n6562 vss.n5919 347.368
R2668 vss.n6477 vss.n5996 347.368
R2669 vss.n6440 vss.n6439 347.368
R2670 vss.n6359 vss.n6094 347.368
R2671 vss.n6315 vss.n6126 347.368
R2672 vss.n6211 vss.n6210 347.368
R2673 vss.n6952 vss.n6951 347.368
R2674 vss.n5578 vss.n4282 347.368
R2675 vss.n5541 vss.n5540 347.368
R2676 vss.n5460 vss.n4380 347.368
R2677 vss.n5416 vss.n4412 347.368
R2678 vss.n5336 vss.n5335 347.368
R2679 vss.n5300 vss.n5299 347.368
R2680 vss.n5219 vss.n4593 347.368
R2681 vss.n5175 vss.n4625 347.368
R2682 vss.n5095 vss.n5094 347.368
R2683 vss.n5059 vss.n5058 347.368
R2684 vss.n4978 vss.n4806 347.368
R2685 vss.n4934 vss.n4838 347.368
R2686 vss.n16749 vss.n16748 347.368
R2687 vss.n16818 vss.n16817 347.368
R2688 vss.n16979 vss.n16978 347.368
R2689 vss.n17052 vss.n17051 347.368
R2690 vss.n17215 vss.n17214 347.368
R2691 vss.n17303 vss.n17302 347.368
R2692 vss.n15298 vss.n15297 347.368
R2693 vss.n15337 vss.n15336 347.368
R2694 vss.n15499 vss.n15498 347.368
R2695 vss.n15574 vss.n15573 347.368
R2696 vss.n15735 vss.n15734 347.368
R2697 vss.n15802 vss.n15801 347.368
R2698 vss.n16446 vss.n16445 347.368
R2699 vss.n16521 vss.n16520 347.368
R2700 vss.n22613 vss.n22612 342.857
R2701 vss.n22566 vss.n22565 342.857
R2702 vss.n22405 vss.n22404 342.857
R2703 vss.n22358 vss.n22357 342.857
R2704 vss.n22197 vss.n22196 342.857
R2705 vss.n22150 vss.n22149 342.857
R2706 vss.n21541 vss.n21540 342.857
R2707 vss.n21494 vss.n21493 342.857
R2708 vss.n21333 vss.n21332 342.857
R2709 vss.n21286 vss.n21285 342.857
R2710 vss.n21125 vss.n21124 342.857
R2711 vss.n21078 vss.n21077 342.857
R2712 vss.n20917 vss.n20916 342.857
R2713 vss.n8776 vss.n8775 342.857
R2714 vss.n8729 vss.n8728 342.857
R2715 vss.n8568 vss.n8567 342.857
R2716 vss.n8521 vss.n8520 342.857
R2717 vss.n8360 vss.n8359 342.857
R2718 vss.n8313 vss.n8312 342.857
R2719 vss.n8152 vss.n8151 342.857
R2720 vss.n8105 vss.n8104 342.857
R2721 vss.n7944 vss.n7943 342.857
R2722 vss.n7897 vss.n7896 342.857
R2723 vss.n7735 vss.n7734 342.857
R2724 vss.n7688 vss.n7687 342.857
R2725 vss.n7527 vss.n7526 342.857
R2726 vss.n20267 vss.n20266 318.421
R2727 vss.n20176 vss.n20175 318.421
R2728 vss.n20143 vss.n19151 318.421
R2729 vss.n20053 vss.n20052 318.421
R2730 vss.n20020 vss.n20019 318.421
R2731 vss.n19929 vss.n19928 318.421
R2732 vss.n19896 vss.n19358 318.421
R2733 vss.n19806 vss.n19805 318.421
R2734 vss.n19773 vss.n19772 318.421
R2735 vss.n19682 vss.n19681 318.421
R2736 vss.n19649 vss.n19565 318.421
R2737 vss.n20323 vss.n17603 318.421
R2738 vss.n18997 vss.n17644 318.421
R2739 vss.n18907 vss.n18906 318.421
R2740 vss.n18874 vss.n18873 318.421
R2741 vss.n18783 vss.n18782 318.421
R2742 vss.n18750 vss.n18749 318.421
R2743 vss.n18666 vss.n18665 318.421
R2744 vss.n18633 vss.n18632 318.421
R2745 vss.n18542 vss.n18541 318.421
R2746 vss.n18509 vss.n18508 318.421
R2747 vss.n18425 vss.n18424 318.421
R2748 vss.n18392 vss.n18391 318.421
R2749 vss.n18301 vss.n18300 318.421
R2750 vss.n6877 vss.n6876 318.421
R2751 vss.n6786 vss.n6785 318.421
R2752 vss.n6753 vss.n5761 318.421
R2753 vss.n6663 vss.n6662 318.421
R2754 vss.n6630 vss.n6629 318.421
R2755 vss.n6539 vss.n6538 318.421
R2756 vss.n6506 vss.n5968 318.421
R2757 vss.n6416 vss.n6415 318.421
R2758 vss.n6383 vss.n6382 318.421
R2759 vss.n6292 vss.n6291 318.421
R2760 vss.n6259 vss.n6175 318.421
R2761 vss.n6933 vss.n4213 318.421
R2762 vss.n5607 vss.n4254 318.421
R2763 vss.n5517 vss.n5516 318.421
R2764 vss.n5484 vss.n5483 318.421
R2765 vss.n5393 vss.n5392 318.421
R2766 vss.n5360 vss.n5359 318.421
R2767 vss.n5276 vss.n5275 318.421
R2768 vss.n5243 vss.n5242 318.421
R2769 vss.n5152 vss.n5151 318.421
R2770 vss.n5119 vss.n5118 318.421
R2771 vss.n5035 vss.n5034 318.421
R2772 vss.n5002 vss.n5001 318.421
R2773 vss.n4911 vss.n4910 318.421
R2774 vss.n16706 vss.n16705 318.421
R2775 vss.n16857 vss.n16856 318.421
R2776 vss.n16936 vss.n16935 318.421
R2777 vss.n17093 vss.n17092 318.421
R2778 vss.n17172 vss.n17171 318.421
R2779 vss.n17310 vss.n17309 318.421
R2780 vss.n15903 vss.n15902 318.421
R2781 vss.n15983 vss.n15982 318.421
R2782 vss.n16139 vss.n16138 318.421
R2783 vss.n16219 vss.n16218 318.421
R2784 vss.n15255 vss.n15254 318.421
R2785 vss.n15379 vss.n15378 318.421
R2786 vss.n15456 vss.n15455 318.421
R2787 vss.n15615 vss.n15614 318.421
R2788 vss.n15692 vss.n15691 318.421
R2789 vss.n15843 vss.n15842 318.421
R2790 vss.n16326 vss.n16325 318.421
R2791 vss.n16403 vss.n16402 318.421
R2792 vss.n16562 vss.n16561 318.421
R2793 vss.n16639 vss.n16638 318.421
R2794 vss.n14325 vss.n14324 316.339
R2795 vss.n13898 vss.n13897 316.339
R2796 vss.n14456 vss.n14455 316.339
R2797 vss.n14426 vss.n14425 316.339
R2798 vss.n13999 vss.n13998 316.339
R2799 vss.n11591 vss.n11590 316.339
R2800 vss.n11734 vss.n11733 316.339
R2801 vss.n11142 vss.n11141 316.339
R2802 vss.n12453 vss.n12452 316.339
R2803 vss.n12615 vss.n12614 316.339
R2804 vss.n12154 vss.n12153 316.339
R2805 vss.n12211 vss.n12210 316.339
R2806 vss.n14638 vss.n14637 316.339
R2807 vss.n13560 vss.n13559 316.339
R2808 vss.n15031 vss.n15030 316.339
R2809 vss.n10476 vss.n10475 316.339
R2810 vss.n13314 vss.n13313 316.339
R2811 vss.n14751 vss.n14750 316.339
R2812 vss.n14918 vss.n14917 316.339
R2813 vss.n14946 vss.n14945 316.339
R2814 vss.n10844 vss.n10843 316.339
R2815 vss.n10888 vss.n10887 316.339
R2816 vss.n11244 vss.n11243 316.339
R2817 vss.n11209 vss.n11208 316.339
R2818 vss.n12920 vss.n12917 307.088
R2819 vss.n12814 vss.n12811 307.088
R2820 vss.n15055 vss.n15052 307.088
R2821 vss.n12507 vss.n12504 307.088
R2822 vss.n12558 vss.n12555 307.088
R2823 vss.n22732 vss.n22731 292.5
R2824 vss.n22718 vss.n22717 292.5
R2825 vss.n22702 vss.n22701 292.5
R2826 vss.n22704 vss.n22703 292.5
R2827 vss.n22681 vss.n22680 292.5
R2828 vss.n22685 vss.n22684 292.5
R2829 vss.n22669 vss.n22668 292.5
R2830 vss.n22655 vss.n22654 292.5
R2831 vss.n22524 vss.n22523 292.5
R2832 vss.n22510 vss.n22509 292.5
R2833 vss.n22494 vss.n22493 292.5
R2834 vss.n22496 vss.n22495 292.5
R2835 vss.n22473 vss.n22472 292.5
R2836 vss.n22477 vss.n22476 292.5
R2837 vss.n22461 vss.n22460 292.5
R2838 vss.n22447 vss.n22446 292.5
R2839 vss.n22316 vss.n22315 292.5
R2840 vss.n22302 vss.n22301 292.5
R2841 vss.n22286 vss.n22285 292.5
R2842 vss.n22288 vss.n22287 292.5
R2843 vss.n22265 vss.n22264 292.5
R2844 vss.n22269 vss.n22268 292.5
R2845 vss.n22253 vss.n22252 292.5
R2846 vss.n22239 vss.n22238 292.5
R2847 vss.n22108 vss.n22107 292.5
R2848 vss.n22094 vss.n22093 292.5
R2849 vss.n22076 vss.n22075 292.5
R2850 vss.n22078 vss.n22077 292.5
R2851 vss.n21595 vss.n21594 292.5
R2852 vss.n21599 vss.n21598 292.5
R2853 vss.n21585 vss.n21584 292.5
R2854 vss.n17404 vss.n17403 292.5
R2855 vss.n21452 vss.n21451 292.5
R2856 vss.n21438 vss.n21437 292.5
R2857 vss.n21422 vss.n21421 292.5
R2858 vss.n21424 vss.n21423 292.5
R2859 vss.n21401 vss.n21400 292.5
R2860 vss.n21405 vss.n21404 292.5
R2861 vss.n21389 vss.n21388 292.5
R2862 vss.n21375 vss.n21374 292.5
R2863 vss.n21244 vss.n21243 292.5
R2864 vss.n21230 vss.n21229 292.5
R2865 vss.n21214 vss.n21213 292.5
R2866 vss.n21216 vss.n21215 292.5
R2867 vss.n21193 vss.n21192 292.5
R2868 vss.n21197 vss.n21196 292.5
R2869 vss.n21181 vss.n21180 292.5
R2870 vss.n21167 vss.n21166 292.5
R2871 vss.n21036 vss.n21035 292.5
R2872 vss.n21022 vss.n21021 292.5
R2873 vss.n21006 vss.n21005 292.5
R2874 vss.n21008 vss.n21007 292.5
R2875 vss.n20985 vss.n20984 292.5
R2876 vss.n20989 vss.n20988 292.5
R2877 vss.n20973 vss.n20972 292.5
R2878 vss.n20959 vss.n20958 292.5
R2879 vss.n20439 vss.n20438 292.5
R2880 vss.n20435 vss.n20434 292.5
R2881 vss.n20433 vss.n20432 292.5
R2882 vss.n20430 vss.n20429 292.5
R2883 vss.n20441 vss.n20440 292.5
R2884 vss.n20450 vss.n20449 292.5
R2885 vss.n20466 vss.n20465 292.5
R2886 vss.n20481 vss.n20480 292.5
R2887 vss.n20496 vss.n20495 292.5
R2888 vss.n20512 vss.n20511 292.5
R2889 vss.n20529 vss.n20528 292.5
R2890 vss.n20557 vss.n20556 292.5
R2891 vss.n20572 vss.n20571 292.5
R2892 vss.n20587 vss.n20586 292.5
R2893 vss.n20602 vss.n20601 292.5
R2894 vss.n20617 vss.n20616 292.5
R2895 vss.n20632 vss.n20631 292.5
R2896 vss.n20647 vss.n20646 292.5
R2897 vss.n17523 vss.n17522 292.5
R2898 vss.n17524 vss.n17523 292.5
R2899 vss.n17511 vss.n17510 292.5
R2900 vss.n20665 vss.n20664 292.5
R2901 vss.n20680 vss.n20679 292.5
R2902 vss.n20695 vss.n20694 292.5
R2903 vss.n20710 vss.n20709 292.5
R2904 vss.n20725 vss.n20724 292.5
R2905 vss.n20740 vss.n20739 292.5
R2906 vss.n20758 vss.n20757 292.5
R2907 vss.n20779 vss.n20778 292.5
R2908 vss.n20794 vss.n20793 292.5
R2909 vss.n20810 vss.n20809 292.5
R2910 vss.n20825 vss.n20824 292.5
R2911 vss.n20840 vss.n20839 292.5
R2912 vss.n20856 vss.n20855 292.5
R2913 vss.n20879 vss.n20878 292.5
R2914 vss.n20881 vss.n20880 292.5
R2915 vss.n20884 vss.n20883 292.5
R2916 vss.n20886 vss.n20885 292.5
R2917 vss.n20890 vss.n20889 292.5
R2918 vss.n17684 vss.n17683 292.5
R2919 vss.n17683 vss.n17682 292.5
R2920 vss.n17791 vss.n17787 292.5
R2921 vss.n18828 vss.n17787 292.5
R2922 vss.n17899 vss.n17898 292.5
R2923 vss.n17901 vss.n17899 292.5
R2924 vss.n18004 vss.n18000 292.5
R2925 vss.n18587 vss.n18000 292.5
R2926 vss.n18112 vss.n18111 292.5
R2927 vss.n18114 vss.n18112 292.5
R2928 vss.n18217 vss.n18213 292.5
R2929 vss.n18346 vss.n18213 292.5
R2930 vss.n17593 vss.n17582 292.5
R2931 vss.n20355 vss.n17593 292.5
R2932 vss.n19091 vss.n19087 292.5
R2933 vss.n20221 vss.n19087 292.5
R2934 vss.n19191 vss.n19190 292.5
R2935 vss.n19190 vss.n19189 292.5
R2936 vss.n19298 vss.n19294 292.5
R2937 vss.n19974 vss.n19294 292.5
R2938 vss.n19397 vss.n19396 292.5
R2939 vss.n19402 vss.n19396 292.5
R2940 vss.n19505 vss.n19501 292.5
R2941 vss.n19727 vss.n19501 292.5
R2942 vss.n9239 vss.n9205 292.5
R2943 vss.n9205 vss.n9204 292.5
R2944 vss.n9242 vss.n9241 292.5
R2945 vss.n9241 vss.n9240 292.5
R2946 vss.n9245 vss.n9244 292.5
R2947 vss.n9244 vss.n9243 292.5
R2948 vss.n9248 vss.n9247 292.5
R2949 vss.n9247 vss.n9246 292.5
R2950 vss.n9251 vss.n9250 292.5
R2951 vss.n9250 vss.n9249 292.5
R2952 vss.n9254 vss.n9253 292.5
R2953 vss.n9253 vss.n9252 292.5
R2954 vss.n9257 vss.n9256 292.5
R2955 vss.n9256 vss.n9255 292.5
R2956 vss.n9260 vss.n9259 292.5
R2957 vss.n9259 vss.n9258 292.5
R2958 vss.n9263 vss.n9262 292.5
R2959 vss.n9262 vss.n9261 292.5
R2960 vss.n9266 vss.n9265 292.5
R2961 vss.n9265 vss.n9264 292.5
R2962 vss.n9269 vss.n9268 292.5
R2963 vss.n9268 vss.n9267 292.5
R2964 vss.n9272 vss.n9271 292.5
R2965 vss.n9271 vss.n9270 292.5
R2966 vss.n9275 vss.n9274 292.5
R2967 vss.n9274 vss.n9273 292.5
R2968 vss.n9278 vss.n9277 292.5
R2969 vss.n9277 vss.n9276 292.5
R2970 vss.n9281 vss.n9280 292.5
R2971 vss.n9280 vss.n9279 292.5
R2972 vss.n9284 vss.n9283 292.5
R2973 vss.n9283 vss.n9282 292.5
R2974 vss.n9287 vss.n9286 292.5
R2975 vss.n9286 vss.n9285 292.5
R2976 vss.n9290 vss.n9289 292.5
R2977 vss.n9289 vss.n9288 292.5
R2978 vss.n9293 vss.n9292 292.5
R2979 vss.n9292 vss.n9291 292.5
R2980 vss.n9296 vss.n9295 292.5
R2981 vss.n9295 vss.n9294 292.5
R2982 vss.n9299 vss.n9298 292.5
R2983 vss.n9298 vss.n9297 292.5
R2984 vss.n9302 vss.n9301 292.5
R2985 vss.n9301 vss.n9300 292.5
R2986 vss.n9305 vss.n9304 292.5
R2987 vss.n9304 vss.n9303 292.5
R2988 vss.n9308 vss.n9307 292.5
R2989 vss.n9307 vss.n9306 292.5
R2990 vss.n9311 vss.n9310 292.5
R2991 vss.n9310 vss.n9309 292.5
R2992 vss.n9314 vss.n9313 292.5
R2993 vss.n9313 vss.n9312 292.5
R2994 vss.n9317 vss.n9316 292.5
R2995 vss.n9316 vss.n9315 292.5
R2996 vss.n9320 vss.n9319 292.5
R2997 vss.n9319 vss.n9318 292.5
R2998 vss.n9323 vss.n9322 292.5
R2999 vss.n9322 vss.n9321 292.5
R3000 vss.n9326 vss.n9325 292.5
R3001 vss.n9325 vss.n9324 292.5
R3002 vss.n9329 vss.n9328 292.5
R3003 vss.n9328 vss.n9327 292.5
R3004 vss.n9332 vss.n9331 292.5
R3005 vss.n9331 vss.n9330 292.5
R3006 vss.n9335 vss.n9334 292.5
R3007 vss.n9334 vss.n9333 292.5
R3008 vss.n9338 vss.n9337 292.5
R3009 vss.n9337 vss.n9336 292.5
R3010 vss.n9341 vss.n9340 292.5
R3011 vss.n9340 vss.n9339 292.5
R3012 vss.n9344 vss.n9343 292.5
R3013 vss.n9343 vss.n9342 292.5
R3014 vss.n9347 vss.n9346 292.5
R3015 vss.n9346 vss.n9345 292.5
R3016 vss.n9350 vss.n9349 292.5
R3017 vss.n9349 vss.n9348 292.5
R3018 vss.n9353 vss.n9352 292.5
R3019 vss.n9352 vss.n9351 292.5
R3020 vss.n9356 vss.n9355 292.5
R3021 vss.n9355 vss.n9354 292.5
R3022 vss.n9359 vss.n9358 292.5
R3023 vss.n9358 vss.n9357 292.5
R3024 vss.n9362 vss.n9361 292.5
R3025 vss.n9361 vss.n9360 292.5
R3026 vss.n9365 vss.n9364 292.5
R3027 vss.n9364 vss.n9363 292.5
R3028 vss.n9368 vss.n9367 292.5
R3029 vss.n9367 vss.n9366 292.5
R3030 vss.n9371 vss.n9370 292.5
R3031 vss.n9370 vss.n9369 292.5
R3032 vss.n9374 vss.n9373 292.5
R3033 vss.n9373 vss.n9372 292.5
R3034 vss.n9377 vss.n9376 292.5
R3035 vss.n9376 vss.n9375 292.5
R3036 vss.n9380 vss.n9379 292.5
R3037 vss.n9379 vss.n9378 292.5
R3038 vss.n9383 vss.n9382 292.5
R3039 vss.n9382 vss.n9381 292.5
R3040 vss.n9386 vss.n9385 292.5
R3041 vss.n9385 vss.n9384 292.5
R3042 vss.n9389 vss.n9388 292.5
R3043 vss.n9388 vss.n9387 292.5
R3044 vss.n9392 vss.n9391 292.5
R3045 vss.n9391 vss.n9390 292.5
R3046 vss.n9395 vss.n9394 292.5
R3047 vss.n9394 vss.n9393 292.5
R3048 vss.n9398 vss.n9397 292.5
R3049 vss.n9397 vss.n9396 292.5
R3050 vss.n9401 vss.n9400 292.5
R3051 vss.n9400 vss.n9399 292.5
R3052 vss.n9404 vss.n9403 292.5
R3053 vss.n9403 vss.n9402 292.5
R3054 vss.n9407 vss.n9406 292.5
R3055 vss.n9406 vss.n9405 292.5
R3056 vss.n9410 vss.n9409 292.5
R3057 vss.n9409 vss.n9408 292.5
R3058 vss.n9413 vss.n9412 292.5
R3059 vss.n9412 vss.n9411 292.5
R3060 vss.n9416 vss.n9415 292.5
R3061 vss.n9415 vss.n9414 292.5
R3062 vss.n9419 vss.n9418 292.5
R3063 vss.n9418 vss.n9417 292.5
R3064 vss.n9422 vss.n9421 292.5
R3065 vss.n9421 vss.n9420 292.5
R3066 vss.n9425 vss.n9424 292.5
R3067 vss.n9424 vss.n9423 292.5
R3068 vss.n9428 vss.n9427 292.5
R3069 vss.n9427 vss.n9426 292.5
R3070 vss.n9431 vss.n9430 292.5
R3071 vss.n9430 vss.n9429 292.5
R3072 vss.n9434 vss.n9433 292.5
R3073 vss.n9433 vss.n9432 292.5
R3074 vss.n9437 vss.n9436 292.5
R3075 vss.n9436 vss.n9435 292.5
R3076 vss.n9440 vss.n9439 292.5
R3077 vss.n9439 vss.n9438 292.5
R3078 vss.n9443 vss.n9442 292.5
R3079 vss.n9442 vss.n9441 292.5
R3080 vss.n9446 vss.n9445 292.5
R3081 vss.n9445 vss.n9444 292.5
R3082 vss.n9449 vss.n9448 292.5
R3083 vss.n9448 vss.n9447 292.5
R3084 vss.n9452 vss.n9451 292.5
R3085 vss.n9451 vss.n9450 292.5
R3086 vss.n9455 vss.n9454 292.5
R3087 vss.n9454 vss.n9453 292.5
R3088 vss.n9458 vss.n9457 292.5
R3089 vss.n9457 vss.n9456 292.5
R3090 vss.n9461 vss.n9460 292.5
R3091 vss.n9460 vss.n9459 292.5
R3092 vss.n9464 vss.n9463 292.5
R3093 vss.n9463 vss.n9462 292.5
R3094 vss.n9467 vss.n9466 292.5
R3095 vss.n9466 vss.n9465 292.5
R3096 vss.n9470 vss.n9469 292.5
R3097 vss.n9469 vss.n9468 292.5
R3098 vss.n9473 vss.n9472 292.5
R3099 vss.n9472 vss.n9471 292.5
R3100 vss.n9476 vss.n9475 292.5
R3101 vss.n9475 vss.n9474 292.5
R3102 vss.n9479 vss.n9478 292.5
R3103 vss.n9478 vss.n9477 292.5
R3104 vss.n9482 vss.n9481 292.5
R3105 vss.n9481 vss.n9480 292.5
R3106 vss.n9485 vss.n9484 292.5
R3107 vss.n9484 vss.n9483 292.5
R3108 vss.n9488 vss.n9487 292.5
R3109 vss.n9487 vss.n9486 292.5
R3110 vss.n9491 vss.n9490 292.5
R3111 vss.n9490 vss.n9489 292.5
R3112 vss.n9494 vss.n9493 292.5
R3113 vss.n9493 vss.n9492 292.5
R3114 vss.n9497 vss.n9496 292.5
R3115 vss.n9496 vss.n9495 292.5
R3116 vss.n9500 vss.n9499 292.5
R3117 vss.n9499 vss.n9498 292.5
R3118 vss.n9503 vss.n9502 292.5
R3119 vss.n9502 vss.n9501 292.5
R3120 vss.n9506 vss.n9505 292.5
R3121 vss.n9505 vss.n9504 292.5
R3122 vss.n9509 vss.n9508 292.5
R3123 vss.n9508 vss.n9507 292.5
R3124 vss.n9512 vss.n9511 292.5
R3125 vss.n9511 vss.n9510 292.5
R3126 vss.n9515 vss.n9514 292.5
R3127 vss.n9514 vss.n9513 292.5
R3128 vss.n9518 vss.n9517 292.5
R3129 vss.n9517 vss.n9516 292.5
R3130 vss.n9521 vss.n9520 292.5
R3131 vss.n9520 vss.n9519 292.5
R3132 vss.n9524 vss.n9523 292.5
R3133 vss.n9523 vss.n9522 292.5
R3134 vss.n9527 vss.n9526 292.5
R3135 vss.n9526 vss.n9525 292.5
R3136 vss.n9530 vss.n9529 292.5
R3137 vss.n9529 vss.n9528 292.5
R3138 vss.n9533 vss.n9532 292.5
R3139 vss.n9532 vss.n9531 292.5
R3140 vss.n9536 vss.n9535 292.5
R3141 vss.n9535 vss.n9534 292.5
R3142 vss.n9539 vss.n9538 292.5
R3143 vss.n9538 vss.n9537 292.5
R3144 vss.n9542 vss.n9541 292.5
R3145 vss.n9541 vss.n9540 292.5
R3146 vss.n9545 vss.n9544 292.5
R3147 vss.n9544 vss.n9543 292.5
R3148 vss.n9548 vss.n9547 292.5
R3149 vss.n9547 vss.n9546 292.5
R3150 vss.n9551 vss.n9550 292.5
R3151 vss.n9550 vss.n9549 292.5
R3152 vss.n9554 vss.n9553 292.5
R3153 vss.n9553 vss.n9552 292.5
R3154 vss.n9557 vss.n9556 292.5
R3155 vss.n9556 vss.n9555 292.5
R3156 vss.n9560 vss.n9559 292.5
R3157 vss.n9559 vss.n9558 292.5
R3158 vss.n9563 vss.n9562 292.5
R3159 vss.n9562 vss.n9561 292.5
R3160 vss.n9566 vss.n9565 292.5
R3161 vss.n9565 vss.n9564 292.5
R3162 vss.n9569 vss.n9568 292.5
R3163 vss.n9568 vss.n9567 292.5
R3164 vss.n9572 vss.n9571 292.5
R3165 vss.n9571 vss.n9570 292.5
R3166 vss.n9575 vss.n9574 292.5
R3167 vss.n9574 vss.n9573 292.5
R3168 vss.n9578 vss.n9577 292.5
R3169 vss.n9577 vss.n9576 292.5
R3170 vss.n9581 vss.n9580 292.5
R3171 vss.n9580 vss.n9579 292.5
R3172 vss.n9584 vss.n9583 292.5
R3173 vss.n9583 vss.n9582 292.5
R3174 vss.n9587 vss.n9586 292.5
R3175 vss.n9586 vss.n9585 292.5
R3176 vss.n9590 vss.n9589 292.5
R3177 vss.n9589 vss.n9588 292.5
R3178 vss.n9593 vss.n9592 292.5
R3179 vss.n9592 vss.n9591 292.5
R3180 vss.n9596 vss.n9595 292.5
R3181 vss.n9595 vss.n9594 292.5
R3182 vss.n9599 vss.n9598 292.5
R3183 vss.n9598 vss.n9597 292.5
R3184 vss.n9602 vss.n9601 292.5
R3185 vss.n9601 vss.n9600 292.5
R3186 vss.n9605 vss.n9604 292.5
R3187 vss.n9604 vss.n9603 292.5
R3188 vss.n9608 vss.n9607 292.5
R3189 vss.n9607 vss.n9606 292.5
R3190 vss.n9611 vss.n9610 292.5
R3191 vss.n9610 vss.n9609 292.5
R3192 vss.n9614 vss.n9613 292.5
R3193 vss.n9613 vss.n9612 292.5
R3194 vss.n9617 vss.n9616 292.5
R3195 vss.n9616 vss.n9615 292.5
R3196 vss.n9620 vss.n9619 292.5
R3197 vss.n9619 vss.n9618 292.5
R3198 vss.n9623 vss.n9622 292.5
R3199 vss.n9622 vss.n9621 292.5
R3200 vss.n9626 vss.n9625 292.5
R3201 vss.n9625 vss.n9624 292.5
R3202 vss.n9629 vss.n9628 292.5
R3203 vss.n9628 vss.n9627 292.5
R3204 vss.n9632 vss.n9631 292.5
R3205 vss.n9631 vss.n9630 292.5
R3206 vss.n9635 vss.n9634 292.5
R3207 vss.n9634 vss.n9633 292.5
R3208 vss.n9779 vss.n9778 292.5
R3209 vss.n9778 vss.n9777 292.5
R3210 vss.n9776 vss.n9775 292.5
R3211 vss.n9775 vss.n9774 292.5
R3212 vss.n9773 vss.n9772 292.5
R3213 vss.n9772 vss.n9771 292.5
R3214 vss.n9770 vss.n9769 292.5
R3215 vss.n9769 vss.n9768 292.5
R3216 vss.n9767 vss.n9766 292.5
R3217 vss.n9766 vss.n9765 292.5
R3218 vss.n9764 vss.n9763 292.5
R3219 vss.n9763 vss.n9762 292.5
R3220 vss.n9761 vss.n9760 292.5
R3221 vss.n9760 vss.n9759 292.5
R3222 vss.n9758 vss.n9757 292.5
R3223 vss.n9757 vss.n9756 292.5
R3224 vss.n9755 vss.n9754 292.5
R3225 vss.n9754 vss.n9753 292.5
R3226 vss.n9752 vss.n9751 292.5
R3227 vss.n9751 vss.n9750 292.5
R3228 vss.n9749 vss.n9748 292.5
R3229 vss.n9748 vss.n9747 292.5
R3230 vss.n9208 vss.n9207 292.5
R3231 vss.n9207 vss.n9206 292.5
R3232 vss.n9211 vss.n9210 292.5
R3233 vss.n9210 vss.n9209 292.5
R3234 vss.n9214 vss.n9213 292.5
R3235 vss.n9213 vss.n9212 292.5
R3236 vss.n9217 vss.n9216 292.5
R3237 vss.n9216 vss.n9215 292.5
R3238 vss.n9220 vss.n9219 292.5
R3239 vss.n9219 vss.n9218 292.5
R3240 vss.n9223 vss.n9222 292.5
R3241 vss.n9222 vss.n9221 292.5
R3242 vss.n9226 vss.n9225 292.5
R3243 vss.n9225 vss.n9224 292.5
R3244 vss.n9229 vss.n9228 292.5
R3245 vss.n9228 vss.n9227 292.5
R3246 vss.n9232 vss.n9231 292.5
R3247 vss.n9231 vss.n9230 292.5
R3248 vss.n9235 vss.n9234 292.5
R3249 vss.n9234 vss.n9233 292.5
R3250 vss.n9238 vss.n9237 292.5
R3251 vss.n9237 vss.n9236 292.5
R3252 vss.n10175 vss.n10174 292.5
R3253 vss.n10174 vss.n10173 292.5
R3254 vss.n10172 vss.n10171 292.5
R3255 vss.n10171 vss.n10170 292.5
R3256 vss.n10169 vss.n10168 292.5
R3257 vss.n10168 vss.n10167 292.5
R3258 vss.n10166 vss.n10165 292.5
R3259 vss.n10165 vss.n10164 292.5
R3260 vss.n10163 vss.n10162 292.5
R3261 vss.n10162 vss.n10161 292.5
R3262 vss.n10160 vss.n10159 292.5
R3263 vss.n10159 vss.n10158 292.5
R3264 vss.n10157 vss.n10156 292.5
R3265 vss.n10156 vss.n10155 292.5
R3266 vss.n10154 vss.n10153 292.5
R3267 vss.n10153 vss.n10152 292.5
R3268 vss.n10151 vss.n10150 292.5
R3269 vss.n10150 vss.n10149 292.5
R3270 vss.n10148 vss.n10147 292.5
R3271 vss.n10147 vss.n10146 292.5
R3272 vss.n10145 vss.n10144 292.5
R3273 vss.n10144 vss.n10143 292.5
R3274 vss.n10142 vss.n10141 292.5
R3275 vss.n10141 vss.n10140 292.5
R3276 vss.n10139 vss.n10138 292.5
R3277 vss.n10138 vss.n10137 292.5
R3278 vss.n10136 vss.n10135 292.5
R3279 vss.n10135 vss.n10134 292.5
R3280 vss.n10133 vss.n10132 292.5
R3281 vss.n10132 vss.n10131 292.5
R3282 vss.n10130 vss.n10129 292.5
R3283 vss.n10129 vss.n10128 292.5
R3284 vss.n10127 vss.n10126 292.5
R3285 vss.n10126 vss.n10125 292.5
R3286 vss.n10124 vss.n10123 292.5
R3287 vss.n10123 vss.n10122 292.5
R3288 vss.n10121 vss.n10120 292.5
R3289 vss.n10120 vss.n10119 292.5
R3290 vss.n10118 vss.n10117 292.5
R3291 vss.n10117 vss.n10116 292.5
R3292 vss.n10115 vss.n10114 292.5
R3293 vss.n10114 vss.n10113 292.5
R3294 vss.n10112 vss.n10111 292.5
R3295 vss.n10111 vss.n10110 292.5
R3296 vss.n10109 vss.n10108 292.5
R3297 vss.n10108 vss.n10107 292.5
R3298 vss.n10106 vss.n10105 292.5
R3299 vss.n10105 vss.n10104 292.5
R3300 vss.n10103 vss.n10102 292.5
R3301 vss.n10102 vss.n10101 292.5
R3302 vss.n10100 vss.n10099 292.5
R3303 vss.n10099 vss.n10098 292.5
R3304 vss.n10097 vss.n10096 292.5
R3305 vss.n10096 vss.n10095 292.5
R3306 vss.n10094 vss.n10093 292.5
R3307 vss.n10093 vss.n10092 292.5
R3308 vss.n10091 vss.n10090 292.5
R3309 vss.n10090 vss.n10089 292.5
R3310 vss.n10088 vss.n10087 292.5
R3311 vss.n10087 vss.n10086 292.5
R3312 vss.n10085 vss.n10084 292.5
R3313 vss.n10084 vss.n10083 292.5
R3314 vss.n10082 vss.n10081 292.5
R3315 vss.n10081 vss.n10080 292.5
R3316 vss.n10079 vss.n10078 292.5
R3317 vss.n10078 vss.n10077 292.5
R3318 vss.n10076 vss.n10075 292.5
R3319 vss.n10075 vss.n10074 292.5
R3320 vss.n10073 vss.n10072 292.5
R3321 vss.n10072 vss.n10071 292.5
R3322 vss.n10070 vss.n10069 292.5
R3323 vss.n10069 vss.n10068 292.5
R3324 vss.n10067 vss.n10066 292.5
R3325 vss.n10066 vss.n10065 292.5
R3326 vss.n10064 vss.n10063 292.5
R3327 vss.n10063 vss.n10062 292.5
R3328 vss.n10061 vss.n10060 292.5
R3329 vss.n10060 vss.n10059 292.5
R3330 vss.n10058 vss.n10057 292.5
R3331 vss.n10057 vss.n10056 292.5
R3332 vss.n10055 vss.n10054 292.5
R3333 vss.n10054 vss.n10053 292.5
R3334 vss.n10052 vss.n10051 292.5
R3335 vss.n10051 vss.n10050 292.5
R3336 vss.n10049 vss.n10048 292.5
R3337 vss.n10048 vss.n10047 292.5
R3338 vss.n10046 vss.n10045 292.5
R3339 vss.n10045 vss.n10044 292.5
R3340 vss.n10043 vss.n10042 292.5
R3341 vss.n10042 vss.n10041 292.5
R3342 vss.n10040 vss.n10039 292.5
R3343 vss.n10039 vss.n10038 292.5
R3344 vss.n10037 vss.n10036 292.5
R3345 vss.n10036 vss.n10035 292.5
R3346 vss.n10034 vss.n10033 292.5
R3347 vss.n10033 vss.n10032 292.5
R3348 vss.n10031 vss.n10030 292.5
R3349 vss.n10030 vss.n10029 292.5
R3350 vss.n10028 vss.n10027 292.5
R3351 vss.n10027 vss.n10026 292.5
R3352 vss.n10025 vss.n10024 292.5
R3353 vss.n10024 vss.n10023 292.5
R3354 vss.n10022 vss.n10021 292.5
R3355 vss.n10021 vss.n10020 292.5
R3356 vss.n10019 vss.n10018 292.5
R3357 vss.n10018 vss.n10017 292.5
R3358 vss.n10016 vss.n10015 292.5
R3359 vss.n10015 vss.n10014 292.5
R3360 vss.n10013 vss.n10012 292.5
R3361 vss.n10012 vss.n10011 292.5
R3362 vss.n10010 vss.n10009 292.5
R3363 vss.n10009 vss.n10008 292.5
R3364 vss.n10007 vss.n10006 292.5
R3365 vss.n10006 vss.n10005 292.5
R3366 vss.n10004 vss.n10003 292.5
R3367 vss.n10003 vss.n10002 292.5
R3368 vss.n10001 vss.n10000 292.5
R3369 vss.n10000 vss.n9999 292.5
R3370 vss.n9998 vss.n9997 292.5
R3371 vss.n9997 vss.n9996 292.5
R3372 vss.n9995 vss.n9994 292.5
R3373 vss.n9994 vss.n9993 292.5
R3374 vss.n9992 vss.n9991 292.5
R3375 vss.n9991 vss.n9990 292.5
R3376 vss.n9989 vss.n9988 292.5
R3377 vss.n9988 vss.n9987 292.5
R3378 vss.n9986 vss.n9985 292.5
R3379 vss.n9985 vss.n9984 292.5
R3380 vss.n9983 vss.n9982 292.5
R3381 vss.n9982 vss.n9981 292.5
R3382 vss.n9980 vss.n9979 292.5
R3383 vss.n9979 vss.n9978 292.5
R3384 vss.n9977 vss.n9976 292.5
R3385 vss.n9976 vss.n9975 292.5
R3386 vss.n9974 vss.n9973 292.5
R3387 vss.n9973 vss.n9972 292.5
R3388 vss.n9971 vss.n9970 292.5
R3389 vss.n9970 vss.n9969 292.5
R3390 vss.n9968 vss.n9967 292.5
R3391 vss.n9967 vss.n9966 292.5
R3392 vss.n9965 vss.n9964 292.5
R3393 vss.n9964 vss.n9963 292.5
R3394 vss.n9962 vss.n9961 292.5
R3395 vss.n9961 vss.n9960 292.5
R3396 vss.n9959 vss.n9958 292.5
R3397 vss.n9958 vss.n9957 292.5
R3398 vss.n9956 vss.n9955 292.5
R3399 vss.n9955 vss.n9954 292.5
R3400 vss.n9953 vss.n9952 292.5
R3401 vss.n9952 vss.n9951 292.5
R3402 vss.n9950 vss.n9949 292.5
R3403 vss.n9949 vss.n9948 292.5
R3404 vss.n9947 vss.n9946 292.5
R3405 vss.n9946 vss.n9945 292.5
R3406 vss.n9944 vss.n9943 292.5
R3407 vss.n9943 vss.n9942 292.5
R3408 vss.n9941 vss.n9940 292.5
R3409 vss.n9940 vss.n9939 292.5
R3410 vss.n9938 vss.n9937 292.5
R3411 vss.n9937 vss.n9936 292.5
R3412 vss.n9935 vss.n9934 292.5
R3413 vss.n9934 vss.n9933 292.5
R3414 vss.n9932 vss.n9931 292.5
R3415 vss.n9931 vss.n9930 292.5
R3416 vss.n9929 vss.n9928 292.5
R3417 vss.n9928 vss.n9927 292.5
R3418 vss.n9926 vss.n9925 292.5
R3419 vss.n9925 vss.n9924 292.5
R3420 vss.n9923 vss.n9922 292.5
R3421 vss.n9922 vss.n9921 292.5
R3422 vss.n9920 vss.n9919 292.5
R3423 vss.n9919 vss.n9918 292.5
R3424 vss.n9917 vss.n9916 292.5
R3425 vss.n9916 vss.n9915 292.5
R3426 vss.n9914 vss.n9913 292.5
R3427 vss.n9913 vss.n9912 292.5
R3428 vss.n9911 vss.n9910 292.5
R3429 vss.n9910 vss.n9909 292.5
R3430 vss.n9908 vss.n9907 292.5
R3431 vss.n9907 vss.n9906 292.5
R3432 vss.n9905 vss.n9904 292.5
R3433 vss.n9904 vss.n9903 292.5
R3434 vss.n9902 vss.n9901 292.5
R3435 vss.n9901 vss.n9900 292.5
R3436 vss.n9899 vss.n9898 292.5
R3437 vss.n9898 vss.n9897 292.5
R3438 vss.n9896 vss.n9895 292.5
R3439 vss.n9895 vss.n9894 292.5
R3440 vss.n9893 vss.n9892 292.5
R3441 vss.n9892 vss.n9891 292.5
R3442 vss.n9890 vss.n9889 292.5
R3443 vss.n9889 vss.n9888 292.5
R3444 vss.n9887 vss.n9886 292.5
R3445 vss.n9886 vss.n9885 292.5
R3446 vss.n9884 vss.n9883 292.5
R3447 vss.n9883 vss.n9882 292.5
R3448 vss.n9881 vss.n9880 292.5
R3449 vss.n9880 vss.n9879 292.5
R3450 vss.n9878 vss.n9877 292.5
R3451 vss.n9877 vss.n9876 292.5
R3452 vss.n9875 vss.n9874 292.5
R3453 vss.n9874 vss.n9873 292.5
R3454 vss.n9872 vss.n9871 292.5
R3455 vss.n9871 vss.n9870 292.5
R3456 vss.n9869 vss.n9868 292.5
R3457 vss.n9868 vss.n9867 292.5
R3458 vss.n9866 vss.n9865 292.5
R3459 vss.n9865 vss.n9864 292.5
R3460 vss.n9863 vss.n9862 292.5
R3461 vss.n9862 vss.n9861 292.5
R3462 vss.n9860 vss.n9859 292.5
R3463 vss.n9859 vss.n9858 292.5
R3464 vss.n9857 vss.n9856 292.5
R3465 vss.n9856 vss.n9855 292.5
R3466 vss.n9854 vss.n9853 292.5
R3467 vss.n9853 vss.n9852 292.5
R3468 vss.n9851 vss.n9850 292.5
R3469 vss.n9850 vss.n9849 292.5
R3470 vss.n9848 vss.n9847 292.5
R3471 vss.n9847 vss.n9846 292.5
R3472 vss.n9845 vss.n9844 292.5
R3473 vss.n9844 vss.n9843 292.5
R3474 vss.n9842 vss.n9841 292.5
R3475 vss.n9841 vss.n9840 292.5
R3476 vss.n9839 vss.n9838 292.5
R3477 vss.n9838 vss.n9837 292.5
R3478 vss.n9836 vss.n9835 292.5
R3479 vss.n9835 vss.n9834 292.5
R3480 vss.n9833 vss.n9832 292.5
R3481 vss.n9832 vss.n9831 292.5
R3482 vss.n9830 vss.n9829 292.5
R3483 vss.n9829 vss.n9828 292.5
R3484 vss.n9827 vss.n9826 292.5
R3485 vss.n9826 vss.n9825 292.5
R3486 vss.n9824 vss.n9823 292.5
R3487 vss.n9823 vss.n9822 292.5
R3488 vss.n9821 vss.n9820 292.5
R3489 vss.n9820 vss.n9819 292.5
R3490 vss.n9818 vss.n9817 292.5
R3491 vss.n9817 vss.n9816 292.5
R3492 vss.n9815 vss.n9814 292.5
R3493 vss.n9814 vss.n9813 292.5
R3494 vss.n9812 vss.n9811 292.5
R3495 vss.n9811 vss.n9810 292.5
R3496 vss.n9809 vss.n9808 292.5
R3497 vss.n9808 vss.n9807 292.5
R3498 vss.n9806 vss.n9805 292.5
R3499 vss.n9805 vss.n9804 292.5
R3500 vss.n9803 vss.n9802 292.5
R3501 vss.n9802 vss.n9801 292.5
R3502 vss.n9800 vss.n9799 292.5
R3503 vss.n9799 vss.n9798 292.5
R3504 vss.n9797 vss.n9796 292.5
R3505 vss.n9796 vss.n9795 292.5
R3506 vss.n9794 vss.n9793 292.5
R3507 vss.n9793 vss.n9792 292.5
R3508 vss.n9791 vss.n9790 292.5
R3509 vss.n9790 vss.n9789 292.5
R3510 vss.n9788 vss.n9787 292.5
R3511 vss.n9787 vss.n9786 292.5
R3512 vss.n9785 vss.n9784 292.5
R3513 vss.n9784 vss.n9783 292.5
R3514 vss.n9782 vss.n9781 292.5
R3515 vss.n9781 vss.n9780 292.5
R3516 vss.n10178 vss.n10177 292.5
R3517 vss.n10177 vss.n10176 292.5
R3518 vss.n12112 vss.n12111 292.5
R3519 vss.n12111 vss.n12110 292.5
R3520 vss.n12134 vss.n12133 292.5
R3521 vss.n12133 vss.n12132 292.5
R3522 vss.n10906 vss.n10905 292.5
R3523 vss.n10905 vss.n10904 292.5
R3524 vss.n10909 vss.n10908 292.5
R3525 vss.n10908 vss.n10907 292.5
R3526 vss.n11583 vss.n11582 292.5
R3527 vss.n11582 vss.n11581 292.5
R3528 vss.n11580 vss.n11579 292.5
R3529 vss.n11579 vss.n11578 292.5
R3530 vss.n14383 vss.n14382 292.5
R3531 vss.n14382 vss.n14381 292.5
R3532 vss.n14380 vss.n14379 292.5
R3533 vss.n14379 vss.n14378 292.5
R3534 vss.n13590 vss.n13589 292.5
R3535 vss.n13589 vss.n13588 292.5
R3536 vss.n13587 vss.n13586 292.5
R3537 vss.n13586 vss.n13585 292.5
R3538 vss.n13262 vss.n13261 292.5
R3539 vss.n13261 vss.n13260 292.5
R3540 vss.n13266 vss.n13265 292.5
R3541 vss.n13265 vss.n13264 292.5
R3542 vss.n14845 vss.n14844 292.5
R3543 vss.n14844 vss.n14843 292.5
R3544 vss.n14848 vss.n14847 292.5
R3545 vss.n14847 vss.n14846 292.5
R3546 vss.n12722 vss.n12721 292.5
R3547 vss.n12721 vss.n12720 292.5
R3548 vss.n12725 vss.n12724 292.5
R3549 vss.n12724 vss.n12723 292.5
R3550 vss.n7049 vss.n7048 292.5
R3551 vss.n7045 vss.n7044 292.5
R3552 vss.n7043 vss.n7042 292.5
R3553 vss.n7040 vss.n7039 292.5
R3554 vss.n7051 vss.n7050 292.5
R3555 vss.n7060 vss.n7059 292.5
R3556 vss.n7076 vss.n7075 292.5
R3557 vss.n7091 vss.n7090 292.5
R3558 vss.n7106 vss.n7105 292.5
R3559 vss.n7122 vss.n7121 292.5
R3560 vss.n7139 vss.n7138 292.5
R3561 vss.n7167 vss.n7166 292.5
R3562 vss.n7182 vss.n7181 292.5
R3563 vss.n7197 vss.n7196 292.5
R3564 vss.n7212 vss.n7211 292.5
R3565 vss.n7227 vss.n7226 292.5
R3566 vss.n7242 vss.n7241 292.5
R3567 vss.n7257 vss.n7256 292.5
R3568 vss.n4133 vss.n4132 292.5
R3569 vss.n4134 vss.n4133 292.5
R3570 vss.n4121 vss.n4120 292.5
R3571 vss.n7275 vss.n7274 292.5
R3572 vss.n7290 vss.n7289 292.5
R3573 vss.n7305 vss.n7304 292.5
R3574 vss.n7320 vss.n7319 292.5
R3575 vss.n7335 vss.n7334 292.5
R3576 vss.n7350 vss.n7349 292.5
R3577 vss.n7368 vss.n7367 292.5
R3578 vss.n7389 vss.n7388 292.5
R3579 vss.n7404 vss.n7403 292.5
R3580 vss.n7420 vss.n7419 292.5
R3581 vss.n7435 vss.n7434 292.5
R3582 vss.n7450 vss.n7449 292.5
R3583 vss.n7466 vss.n7465 292.5
R3584 vss.n7489 vss.n7488 292.5
R3585 vss.n7491 vss.n7490 292.5
R3586 vss.n7494 vss.n7493 292.5
R3587 vss.n7496 vss.n7495 292.5
R3588 vss.n7500 vss.n7499 292.5
R3589 vss.n4294 vss.n4293 292.5
R3590 vss.n4293 vss.n4292 292.5
R3591 vss.n4401 vss.n4397 292.5
R3592 vss.n5438 vss.n4397 292.5
R3593 vss.n4509 vss.n4508 292.5
R3594 vss.n4511 vss.n4509 292.5
R3595 vss.n4614 vss.n4610 292.5
R3596 vss.n5197 vss.n4610 292.5
R3597 vss.n4722 vss.n4721 292.5
R3598 vss.n4724 vss.n4722 292.5
R3599 vss.n4827 vss.n4823 292.5
R3600 vss.n4956 vss.n4823 292.5
R3601 vss.n4203 vss.n4192 292.5
R3602 vss.n6965 vss.n4203 292.5
R3603 vss.n5701 vss.n5697 292.5
R3604 vss.n6831 vss.n5697 292.5
R3605 vss.n5801 vss.n5800 292.5
R3606 vss.n5800 vss.n5799 292.5
R3607 vss.n5908 vss.n5904 292.5
R3608 vss.n6584 vss.n5904 292.5
R3609 vss.n6007 vss.n6006 292.5
R3610 vss.n6012 vss.n6006 292.5
R3611 vss.n6115 vss.n6111 292.5
R3612 vss.n6337 vss.n6111 292.5
R3613 vss.n8895 vss.n8894 292.5
R3614 vss.n8881 vss.n8880 292.5
R3615 vss.n8865 vss.n8864 292.5
R3616 vss.n8867 vss.n8866 292.5
R3617 vss.n8844 vss.n8843 292.5
R3618 vss.n8848 vss.n8847 292.5
R3619 vss.n8832 vss.n8831 292.5
R3620 vss.n8818 vss.n8817 292.5
R3621 vss.n8687 vss.n8686 292.5
R3622 vss.n8673 vss.n8672 292.5
R3623 vss.n8657 vss.n8656 292.5
R3624 vss.n8659 vss.n8658 292.5
R3625 vss.n8636 vss.n8635 292.5
R3626 vss.n8640 vss.n8639 292.5
R3627 vss.n8624 vss.n8623 292.5
R3628 vss.n8610 vss.n8609 292.5
R3629 vss.n8479 vss.n8478 292.5
R3630 vss.n8465 vss.n8464 292.5
R3631 vss.n8449 vss.n8448 292.5
R3632 vss.n8451 vss.n8450 292.5
R3633 vss.n8428 vss.n8427 292.5
R3634 vss.n8432 vss.n8431 292.5
R3635 vss.n8416 vss.n8415 292.5
R3636 vss.n8402 vss.n8401 292.5
R3637 vss.n8271 vss.n8270 292.5
R3638 vss.n8257 vss.n8256 292.5
R3639 vss.n8236 vss.n8235 292.5
R3640 vss.n8238 vss.n8237 292.5
R3641 vss.n8221 vss.n8220 292.5
R3642 vss.n8225 vss.n8224 292.5
R3643 vss.n8208 vss.n8207 292.5
R3644 vss.n8194 vss.n8193 292.5
R3645 vss.n8063 vss.n8062 292.5
R3646 vss.n8049 vss.n8048 292.5
R3647 vss.n8033 vss.n8032 292.5
R3648 vss.n8035 vss.n8034 292.5
R3649 vss.n8012 vss.n8011 292.5
R3650 vss.n8016 vss.n8015 292.5
R3651 vss.n8000 vss.n7999 292.5
R3652 vss.n7986 vss.n7985 292.5
R3653 vss.n7855 vss.n7854 292.5
R3654 vss.n7840 vss.n7839 292.5
R3655 vss.n7824 vss.n7823 292.5
R3656 vss.n7826 vss.n7825 292.5
R3657 vss.n7803 vss.n7802 292.5
R3658 vss.n7807 vss.n7806 292.5
R3659 vss.n7791 vss.n7790 292.5
R3660 vss.n7777 vss.n7776 292.5
R3661 vss.n7646 vss.n7645 292.5
R3662 vss.n7632 vss.n7631 292.5
R3663 vss.n7616 vss.n7615 292.5
R3664 vss.n7618 vss.n7617 292.5
R3665 vss.n7595 vss.n7594 292.5
R3666 vss.n7599 vss.n7598 292.5
R3667 vss.n7583 vss.n7582 292.5
R3668 vss.n7569 vss.n7568 292.5
R3669 vss.n1679 vss.n1678 292.5
R3670 vss.n1675 vss.n1674 292.5
R3671 vss.n1673 vss.n1672 292.5
R3672 vss.n1670 vss.n1669 292.5
R3673 vss.n1681 vss.n1680 292.5
R3674 vss.n1689 vss.n1688 292.5
R3675 vss.n1704 vss.n1703 292.5
R3676 vss.n1719 vss.n1718 292.5
R3677 vss.n1734 vss.n1733 292.5
R3678 vss.n1755 vss.n1754 292.5
R3679 vss.n1776 vss.n1775 292.5
R3680 vss.n1793 vss.n1792 292.5
R3681 vss.n1808 vss.n1807 292.5
R3682 vss.n1823 vss.n1822 292.5
R3683 vss.n1838 vss.n1837 292.5
R3684 vss.n1853 vss.n1852 292.5
R3685 vss.n1868 vss.n1867 292.5
R3686 vss.n1645 vss.n1644 292.5
R3687 vss.n1646 vss.n1645 292.5
R3688 vss.n1633 vss.n1632 292.5
R3689 vss.n1634 vss.n1633 292.5
R3690 vss.n1886 vss.n1885 292.5
R3691 vss.n1887 vss.n1886 292.5
R3692 vss.n1902 vss.n1901 292.5
R3693 vss.n1903 vss.n1902 292.5
R3694 vss.n1918 vss.n1917 292.5
R3695 vss.n1919 vss.n1918 292.5
R3696 vss.n1934 vss.n1933 292.5
R3697 vss.n1935 vss.n1934 292.5
R3698 vss.n1950 vss.n1949 292.5
R3699 vss.n1951 vss.n1950 292.5
R3700 vss.n1966 vss.n1965 292.5
R3701 vss.n1967 vss.n1966 292.5
R3702 vss.n1985 vss.n1984 292.5
R3703 vss.n1986 vss.n1985 292.5
R3704 vss.n2015 vss.n2014 292.5
R3705 vss.n2016 vss.n2015 292.5
R3706 vss.n2031 vss.n2030 292.5
R3707 vss.n2032 vss.n2031 292.5
R3708 vss.n2047 vss.n2046 292.5
R3709 vss.n2048 vss.n2047 292.5
R3710 vss.n2063 vss.n2062 292.5
R3711 vss.n2064 vss.n2063 292.5
R3712 vss.n2079 vss.n2078 292.5
R3713 vss.n2080 vss.n2079 292.5
R3714 vss.n2095 vss.n2094 292.5
R3715 vss.n2096 vss.n2095 292.5
R3716 vss.n2112 vss.n2111 292.5
R3717 vss.n2113 vss.n2112 292.5
R3718 vss.n1618 vss.n1617 292.5
R3719 vss.n1619 vss.n1618 292.5
R3720 vss.n1606 vss.n1605 292.5
R3721 vss.n1607 vss.n1606 292.5
R3722 vss.n2130 vss.n2129 292.5
R3723 vss.n2131 vss.n2130 292.5
R3724 vss.n2146 vss.n2145 292.5
R3725 vss.n2147 vss.n2146 292.5
R3726 vss.n2162 vss.n2161 292.5
R3727 vss.n2163 vss.n2162 292.5
R3728 vss.n2178 vss.n2177 292.5
R3729 vss.n2179 vss.n2178 292.5
R3730 vss.n2195 vss.n2194 292.5
R3731 vss.n2196 vss.n2195 292.5
R3732 vss.n2211 vss.n2210 292.5
R3733 vss.n2212 vss.n2211 292.5
R3734 vss.n2230 vss.n2229 292.5
R3735 vss.n2231 vss.n2230 292.5
R3736 vss.n2259 vss.n2258 292.5
R3737 vss.n2260 vss.n2259 292.5
R3738 vss.n2275 vss.n2274 292.5
R3739 vss.n2276 vss.n2275 292.5
R3740 vss.n2291 vss.n2290 292.5
R3741 vss.n2292 vss.n2291 292.5
R3742 vss.n2308 vss.n2307 292.5
R3743 vss.n2309 vss.n2308 292.5
R3744 vss.n2324 vss.n2323 292.5
R3745 vss.n2325 vss.n2324 292.5
R3746 vss.n2340 vss.n2339 292.5
R3747 vss.n2341 vss.n2340 292.5
R3748 vss.n2356 vss.n2355 292.5
R3749 vss.n2357 vss.n2356 292.5
R3750 vss.n1593 vss.n1592 292.5
R3751 vss.n1594 vss.n1593 292.5
R3752 vss.n1581 vss.n1580 292.5
R3753 vss.n1582 vss.n1581 292.5
R3754 vss.n2374 vss.n2373 292.5
R3755 vss.n2375 vss.n2374 292.5
R3756 vss.n2390 vss.n2389 292.5
R3757 vss.n2391 vss.n2390 292.5
R3758 vss.n2407 vss.n2406 292.5
R3759 vss.n2408 vss.n2407 292.5
R3760 vss.n2423 vss.n2422 292.5
R3761 vss.n2424 vss.n2423 292.5
R3762 vss.n2439 vss.n2438 292.5
R3763 vss.n2440 vss.n2439 292.5
R3764 vss.n2455 vss.n2454 292.5
R3765 vss.n2456 vss.n2455 292.5
R3766 vss.n2474 vss.n2473 292.5
R3767 vss.n2475 vss.n2474 292.5
R3768 vss.n2503 vss.n2502 292.5
R3769 vss.n2504 vss.n2503 292.5
R3770 vss.n2520 vss.n2519 292.5
R3771 vss.n2521 vss.n2520 292.5
R3772 vss.n2536 vss.n2535 292.5
R3773 vss.n2537 vss.n2536 292.5
R3774 vss.n2552 vss.n2551 292.5
R3775 vss.n2553 vss.n2552 292.5
R3776 vss.n2568 vss.n2567 292.5
R3777 vss.n2569 vss.n2568 292.5
R3778 vss.n2584 vss.n2583 292.5
R3779 vss.n2585 vss.n2584 292.5
R3780 vss.n2600 vss.n2599 292.5
R3781 vss.n2601 vss.n2600 292.5
R3782 vss.n1568 vss.n1567 292.5
R3783 vss.n1569 vss.n1568 292.5
R3784 vss.n1555 vss.n1554 292.5
R3785 vss.n1556 vss.n1555 292.5
R3786 vss.n2619 vss.n2618 292.5
R3787 vss.n2620 vss.n2619 292.5
R3788 vss.n2635 vss.n2634 292.5
R3789 vss.n2636 vss.n2635 292.5
R3790 vss.n2651 vss.n2650 292.5
R3791 vss.n2652 vss.n2651 292.5
R3792 vss.n2667 vss.n2666 292.5
R3793 vss.n2668 vss.n2667 292.5
R3794 vss.n2683 vss.n2682 292.5
R3795 vss.n2684 vss.n2683 292.5
R3796 vss.n2699 vss.n2698 292.5
R3797 vss.n2700 vss.n2699 292.5
R3798 vss.n2719 vss.n2718 292.5
R3799 vss.n2720 vss.n2719 292.5
R3800 vss.n2748 vss.n2747 292.5
R3801 vss.n2749 vss.n2748 292.5
R3802 vss.n2764 vss.n2763 292.5
R3803 vss.n2765 vss.n2764 292.5
R3804 vss.n2780 vss.n2779 292.5
R3805 vss.n2781 vss.n2780 292.5
R3806 vss.n2796 vss.n2795 292.5
R3807 vss.n2797 vss.n2796 292.5
R3808 vss.n2812 vss.n2811 292.5
R3809 vss.n2827 vss.n2826 292.5
R3810 vss.n2839 vss.n2838 292.5
R3811 vss.n1538 vss.n1537 292.5
R3812 vss.n1539 vss.n1538 292.5
R3813 vss.n1523 vss.n1522 292.5
R3814 vss.n1524 vss.n1523 292.5
R3815 vss.n2857 vss.n2856 292.5
R3816 vss.n2858 vss.n2857 292.5
R3817 vss.n2873 vss.n2872 292.5
R3818 vss.n2874 vss.n2873 292.5
R3819 vss.n2889 vss.n2888 292.5
R3820 vss.n2890 vss.n2889 292.5
R3821 vss.n2905 vss.n2904 292.5
R3822 vss.n2906 vss.n2905 292.5
R3823 vss.n2922 vss.n2921 292.5
R3824 vss.n2923 vss.n2922 292.5
R3825 vss.n2938 vss.n2937 292.5
R3826 vss.n2939 vss.n2938 292.5
R3827 vss.n2957 vss.n2956 292.5
R3828 vss.n2958 vss.n2957 292.5
R3829 vss.n2986 vss.n2985 292.5
R3830 vss.n2987 vss.n2986 292.5
R3831 vss.n3002 vss.n3001 292.5
R3832 vss.n3003 vss.n3002 292.5
R3833 vss.n3019 vss.n3018 292.5
R3834 vss.n3020 vss.n3019 292.5
R3835 vss.n3035 vss.n3034 292.5
R3836 vss.n3036 vss.n3035 292.5
R3837 vss.n3051 vss.n3050 292.5
R3838 vss.n3052 vss.n3051 292.5
R3839 vss.n3067 vss.n3066 292.5
R3840 vss.n3068 vss.n3067 292.5
R3841 vss.n3083 vss.n3082 292.5
R3842 vss.n3084 vss.n3083 292.5
R3843 vss.n1510 vss.n1509 292.5
R3844 vss.n1511 vss.n1510 292.5
R3845 vss.n1498 vss.n1497 292.5
R3846 vss.n1499 vss.n1498 292.5
R3847 vss.n3101 vss.n3100 292.5
R3848 vss.n3102 vss.n3101 292.5
R3849 vss.n3118 vss.n3117 292.5
R3850 vss.n3119 vss.n3118 292.5
R3851 vss.n3134 vss.n3133 292.5
R3852 vss.n3135 vss.n3134 292.5
R3853 vss.n3150 vss.n3149 292.5
R3854 vss.n3151 vss.n3150 292.5
R3855 vss.n3166 vss.n3165 292.5
R3856 vss.n3167 vss.n3166 292.5
R3857 vss.n3182 vss.n3181 292.5
R3858 vss.n3183 vss.n3182 292.5
R3859 vss.n3201 vss.n3200 292.5
R3860 vss.n3202 vss.n3201 292.5
R3861 vss.n3231 vss.n3230 292.5
R3862 vss.n3232 vss.n3231 292.5
R3863 vss.n3247 vss.n3246 292.5
R3864 vss.n3248 vss.n3247 292.5
R3865 vss.n3263 vss.n3262 292.5
R3866 vss.n3264 vss.n3263 292.5
R3867 vss.n3279 vss.n3278 292.5
R3868 vss.n3280 vss.n3279 292.5
R3869 vss.n3295 vss.n3294 292.5
R3870 vss.n3296 vss.n3295 292.5
R3871 vss.n3311 vss.n3310 292.5
R3872 vss.n3312 vss.n3311 292.5
R3873 vss.n3327 vss.n3326 292.5
R3874 vss.n3328 vss.n3327 292.5
R3875 vss.n1483 vss.n1482 292.5
R3876 vss.n1484 vss.n1483 292.5
R3877 vss.n1471 vss.n1470 292.5
R3878 vss.n1472 vss.n1471 292.5
R3879 vss.n3346 vss.n3345 292.5
R3880 vss.n3361 vss.n3360 292.5
R3881 vss.n3376 vss.n3375 292.5
R3882 vss.n3391 vss.n3390 292.5
R3883 vss.n3406 vss.n3405 292.5
R3884 vss.n3421 vss.n3420 292.5
R3885 vss.n15204 vss.n15203 292.5
R3886 vss.n15185 vss.n15184 292.5
R3887 vss.n3462 vss.n3461 292.5
R3888 vss.n3473 vss.n3472 292.5
R3889 vss.n15164 vss.n15163 292.5
R3890 vss.n3485 vss.n3484 292.5
R3891 vss.n15142 vss.n15141 292.5
R3892 vss.n15144 vss.n15143 292.5
R3893 vss.n15147 vss.n15146 292.5
R3894 vss.n15149 vss.n15148 292.5
R3895 vss.n15153 vss.n15152 292.5
R3896 vss.n16486 vss.n16485 292.5
R3897 vss.n16788 vss.n16787 292.5
R3898 vss.n17019 vss.n17018 292.5
R3899 vss.n17257 vss.n17256 292.5
R3900 vss.n16025 vss.n16024 292.5
R3901 vss.n16039 vss.n16038 292.5
R3902 vss.n16053 vss.n16052 292.5
R3903 vss.n16065 vss.n16064 292.5
R3904 vss.n16069 vss.n16068 292.5
R3905 vss.n16083 vss.n16082 292.5
R3906 vss.n16097 vss.n16096 292.5
R3907 vss.n15233 vss.n15232 292.5
R3908 vss.n15539 vss.n15538 292.5
R3909 vss.n15773 vss.n15772 292.5
R3910 vss.n140 vss.n139 292.5
R3911 vss.n136 vss.n135 292.5
R3912 vss.n134 vss.n133 292.5
R3913 vss.n131 vss.n130 292.5
R3914 vss.n142 vss.n141 292.5
R3915 vss.n150 vss.n149 292.5
R3916 vss.n165 vss.n164 292.5
R3917 vss.n180 vss.n179 292.5
R3918 vss.n195 vss.n194 292.5
R3919 vss.n216 vss.n215 292.5
R3920 vss.n237 vss.n236 292.5
R3921 vss.n254 vss.n253 292.5
R3922 vss.n269 vss.n268 292.5
R3923 vss.n284 vss.n283 292.5
R3924 vss.n299 vss.n298 292.5
R3925 vss.n314 vss.n313 292.5
R3926 vss.n329 vss.n328 292.5
R3927 vss.n106 vss.n105 292.5
R3928 vss.n107 vss.n106 292.5
R3929 vss.n94 vss.n93 292.5
R3930 vss.n95 vss.n94 292.5
R3931 vss.n347 vss.n346 292.5
R3932 vss.n348 vss.n347 292.5
R3933 vss.n363 vss.n362 292.5
R3934 vss.n364 vss.n363 292.5
R3935 vss.n379 vss.n378 292.5
R3936 vss.n380 vss.n379 292.5
R3937 vss.n395 vss.n394 292.5
R3938 vss.n396 vss.n395 292.5
R3939 vss.n411 vss.n410 292.5
R3940 vss.n412 vss.n411 292.5
R3941 vss.n427 vss.n426 292.5
R3942 vss.n428 vss.n427 292.5
R3943 vss.n446 vss.n445 292.5
R3944 vss.n447 vss.n446 292.5
R3945 vss.n476 vss.n475 292.5
R3946 vss.n477 vss.n476 292.5
R3947 vss.n492 vss.n491 292.5
R3948 vss.n493 vss.n492 292.5
R3949 vss.n508 vss.n507 292.5
R3950 vss.n509 vss.n508 292.5
R3951 vss.n524 vss.n523 292.5
R3952 vss.n525 vss.n524 292.5
R3953 vss.n540 vss.n539 292.5
R3954 vss.n541 vss.n540 292.5
R3955 vss.n556 vss.n555 292.5
R3956 vss.n557 vss.n556 292.5
R3957 vss.n573 vss.n572 292.5
R3958 vss.n574 vss.n573 292.5
R3959 vss.n79 vss.n78 292.5
R3960 vss.n80 vss.n79 292.5
R3961 vss.n67 vss.n66 292.5
R3962 vss.n68 vss.n67 292.5
R3963 vss.n591 vss.n590 292.5
R3964 vss.n592 vss.n591 292.5
R3965 vss.n607 vss.n606 292.5
R3966 vss.n608 vss.n607 292.5
R3967 vss.n623 vss.n622 292.5
R3968 vss.n624 vss.n623 292.5
R3969 vss.n639 vss.n638 292.5
R3970 vss.n640 vss.n639 292.5
R3971 vss.n656 vss.n655 292.5
R3972 vss.n657 vss.n656 292.5
R3973 vss.n672 vss.n671 292.5
R3974 vss.n673 vss.n672 292.5
R3975 vss.n691 vss.n690 292.5
R3976 vss.n692 vss.n691 292.5
R3977 vss.n720 vss.n719 292.5
R3978 vss.n721 vss.n720 292.5
R3979 vss.n736 vss.n735 292.5
R3980 vss.n737 vss.n736 292.5
R3981 vss.n752 vss.n751 292.5
R3982 vss.n753 vss.n752 292.5
R3983 vss.n769 vss.n768 292.5
R3984 vss.n770 vss.n769 292.5
R3985 vss.n785 vss.n784 292.5
R3986 vss.n786 vss.n785 292.5
R3987 vss.n801 vss.n800 292.5
R3988 vss.n802 vss.n801 292.5
R3989 vss.n817 vss.n816 292.5
R3990 vss.n818 vss.n817 292.5
R3991 vss.n54 vss.n53 292.5
R3992 vss.n55 vss.n54 292.5
R3993 vss.n42 vss.n41 292.5
R3994 vss.n43 vss.n42 292.5
R3995 vss.n835 vss.n834 292.5
R3996 vss.n836 vss.n835 292.5
R3997 vss.n851 vss.n850 292.5
R3998 vss.n852 vss.n851 292.5
R3999 vss.n868 vss.n867 292.5
R4000 vss.n869 vss.n868 292.5
R4001 vss.n884 vss.n883 292.5
R4002 vss.n885 vss.n884 292.5
R4003 vss.n900 vss.n899 292.5
R4004 vss.n901 vss.n900 292.5
R4005 vss.n916 vss.n915 292.5
R4006 vss.n917 vss.n916 292.5
R4007 vss.n935 vss.n934 292.5
R4008 vss.n936 vss.n935 292.5
R4009 vss.n964 vss.n963 292.5
R4010 vss.n965 vss.n964 292.5
R4011 vss.n981 vss.n980 292.5
R4012 vss.n982 vss.n981 292.5
R4013 vss.n997 vss.n996 292.5
R4014 vss.n998 vss.n997 292.5
R4015 vss.n1013 vss.n1012 292.5
R4016 vss.n1014 vss.n1013 292.5
R4017 vss.n1029 vss.n1028 292.5
R4018 vss.n1030 vss.n1029 292.5
R4019 vss.n1045 vss.n1044 292.5
R4020 vss.n1046 vss.n1045 292.5
R4021 vss.n1061 vss.n1060 292.5
R4022 vss.n1062 vss.n1061 292.5
R4023 vss.n29 vss.n28 292.5
R4024 vss.n30 vss.n29 292.5
R4025 vss.n16 vss.n15 292.5
R4026 vss.n17 vss.n16 292.5
R4027 vss.n1080 vss.n1079 292.5
R4028 vss.n1081 vss.n1080 292.5
R4029 vss.n1096 vss.n1095 292.5
R4030 vss.n1097 vss.n1096 292.5
R4031 vss.n1112 vss.n1111 292.5
R4032 vss.n1113 vss.n1112 292.5
R4033 vss.n1128 vss.n1127 292.5
R4034 vss.n1129 vss.n1128 292.5
R4035 vss.n1144 vss.n1143 292.5
R4036 vss.n1145 vss.n1144 292.5
R4037 vss.n1160 vss.n1159 292.5
R4038 vss.n1161 vss.n1160 292.5
R4039 vss.n1180 vss.n1179 292.5
R4040 vss.n1181 vss.n1180 292.5
R4041 vss.n1209 vss.n1208 292.5
R4042 vss.n1210 vss.n1209 292.5
R4043 vss.n1225 vss.n1224 292.5
R4044 vss.n1226 vss.n1225 292.5
R4045 vss.n1241 vss.n1240 292.5
R4046 vss.n1242 vss.n1241 292.5
R4047 vss.n1257 vss.n1256 292.5
R4048 vss.n1258 vss.n1257 292.5
R4049 vss.n1273 vss.n1272 292.5
R4050 vss.n1274 vss.n1273 292.5
R4051 vss.n1290 vss.n1289 292.5
R4052 vss.n1291 vss.n1290 292.5
R4053 vss.n1306 vss.n1305 292.5
R4054 vss.n1307 vss.n1306 292.5
R4055 vss.n1318 vss.n1317 292.5
R4056 vss.n1319 vss.n1318 292.5
R4057 vss.n1330 vss.n1329 292.5
R4058 vss.n1331 vss.n1330 292.5
R4059 vss.n23400 vss.n23399 292.5
R4060 vss.n23401 vss.n23400 292.5
R4061 vss.n23384 vss.n23383 292.5
R4062 vss.n23385 vss.n23384 292.5
R4063 vss.n23368 vss.n23367 292.5
R4064 vss.n23369 vss.n23368 292.5
R4065 vss.n23352 vss.n23351 292.5
R4066 vss.n23353 vss.n23352 292.5
R4067 vss.n23336 vss.n23335 292.5
R4068 vss.n23337 vss.n23336 292.5
R4069 vss.n23320 vss.n23319 292.5
R4070 vss.n23321 vss.n23320 292.5
R4071 vss.n23303 vss.n23302 292.5
R4072 vss.n23304 vss.n23303 292.5
R4073 vss.n23276 vss.n23275 292.5
R4074 vss.n23277 vss.n23276 292.5
R4075 vss.n23256 vss.n23255 292.5
R4076 vss.n23257 vss.n23256 292.5
R4077 vss.n23239 vss.n23238 292.5
R4078 vss.n23240 vss.n23239 292.5
R4079 vss.n23223 vss.n23222 292.5
R4080 vss.n23224 vss.n23223 292.5
R4081 vss.n23207 vss.n23206 292.5
R4082 vss.n23208 vss.n23207 292.5
R4083 vss.n23191 vss.n23190 292.5
R4084 vss.n23192 vss.n23191 292.5
R4085 vss.n23175 vss.n23174 292.5
R4086 vss.n23176 vss.n23175 292.5
R4087 vss.n1344 vss.n1343 292.5
R4088 vss.n1345 vss.n1344 292.5
R4089 vss.n1356 vss.n1355 292.5
R4090 vss.n1357 vss.n1356 292.5
R4091 vss.n23157 vss.n23156 292.5
R4092 vss.n23158 vss.n23157 292.5
R4093 vss.n23140 vss.n23139 292.5
R4094 vss.n23141 vss.n23140 292.5
R4095 vss.n23124 vss.n23123 292.5
R4096 vss.n23125 vss.n23124 292.5
R4097 vss.n23108 vss.n23107 292.5
R4098 vss.n23109 vss.n23108 292.5
R4099 vss.n23092 vss.n23091 292.5
R4100 vss.n23093 vss.n23092 292.5
R4101 vss.n23076 vss.n23075 292.5
R4102 vss.n23077 vss.n23076 292.5
R4103 vss.n23059 vss.n23058 292.5
R4104 vss.n23060 vss.n23059 292.5
R4105 vss.n23031 vss.n23030 292.5
R4106 vss.n23032 vss.n23031 292.5
R4107 vss.n23011 vss.n23010 292.5
R4108 vss.n23012 vss.n23011 292.5
R4109 vss.n22995 vss.n22994 292.5
R4110 vss.n22996 vss.n22995 292.5
R4111 vss.n22979 vss.n22978 292.5
R4112 vss.n22980 vss.n22979 292.5
R4113 vss.n22963 vss.n22962 292.5
R4114 vss.n22964 vss.n22963 292.5
R4115 vss.n22947 vss.n22946 292.5
R4116 vss.n22948 vss.n22947 292.5
R4117 vss.n22931 vss.n22930 292.5
R4118 vss.n22932 vss.n22931 292.5
R4119 vss.n1371 vss.n1370 292.5
R4120 vss.n1372 vss.n1371 292.5
R4121 vss.n1383 vss.n1382 292.5
R4122 vss.n1384 vss.n1383 292.5
R4123 vss.n22913 vss.n22912 292.5
R4124 vss.n22898 vss.n22897 292.5
R4125 vss.n22883 vss.n22882 292.5
R4126 vss.n22868 vss.n22867 292.5
R4127 vss.n22853 vss.n22852 292.5
R4128 vss.n22836 vss.n22835 292.5
R4129 vss.n1397 vss.n1396 292.5
R4130 vss.n22819 vss.n22818 292.5
R4131 vss.n1437 vss.n1436 292.5
R4132 vss.n1448 vss.n1447 292.5
R4133 vss.n22798 vss.n22797 292.5
R4134 vss.n1460 vss.n1459 292.5
R4135 vss.n22776 vss.n22775 292.5
R4136 vss.n22778 vss.n22777 292.5
R4137 vss.n22781 vss.n22780 292.5
R4138 vss.n22783 vss.n22782 292.5
R4139 vss.n22787 vss.n22786 292.5
R4140 vss.n20351 vss.n17575 292.009
R4141 vss.n6961 vss.n4185 292.009
R4142 vss.n20345 vss.n17575 291.03
R4143 vss.n6955 vss.n4185 291.03
R4144 vss.n20338 vss.n17575 290.059
R4145 vss.n6948 vss.n4185 290.059
R4146 vss.n20245 vss.n19069 289.473
R4147 vss.n20197 vss.n19108 289.473
R4148 vss.n20124 vss.n20123 289.473
R4149 vss.n20065 vss.n19209 289.473
R4150 vss.n19998 vss.n19276 289.473
R4151 vss.n19950 vss.n19315 289.473
R4152 vss.n19877 vss.n19876 289.473
R4153 vss.n19818 vss.n19416 289.473
R4154 vss.n19751 vss.n19483 289.473
R4155 vss.n19703 vss.n19522 289.473
R4156 vss.n19630 vss.n19629 289.473
R4157 vss.n20335 vss.n17599 289.473
R4158 vss.n18978 vss.n18977 289.473
R4159 vss.n18919 vss.n17702 289.473
R4160 vss.n18852 vss.n17769 289.473
R4161 vss.n18804 vss.n17808 289.473
R4162 vss.n18737 vss.n17870 289.473
R4163 vss.n18678 vss.n17915 289.473
R4164 vss.n18611 vss.n17982 289.473
R4165 vss.n18563 vss.n18021 289.473
R4166 vss.n18496 vss.n18083 289.473
R4167 vss.n18437 vss.n18128 289.473
R4168 vss.n18370 vss.n18195 289.473
R4169 vss.n18322 vss.n18234 289.473
R4170 vss.n6855 vss.n5679 289.473
R4171 vss.n6807 vss.n5718 289.473
R4172 vss.n6734 vss.n6733 289.473
R4173 vss.n6675 vss.n5819 289.473
R4174 vss.n6608 vss.n5886 289.473
R4175 vss.n6560 vss.n5925 289.473
R4176 vss.n6487 vss.n6486 289.473
R4177 vss.n6428 vss.n6026 289.473
R4178 vss.n6361 vss.n6093 289.473
R4179 vss.n6313 vss.n6132 289.473
R4180 vss.n6240 vss.n6239 289.473
R4181 vss.n6945 vss.n4209 289.473
R4182 vss.n5588 vss.n5587 289.473
R4183 vss.n5529 vss.n4312 289.473
R4184 vss.n5462 vss.n4379 289.473
R4185 vss.n5414 vss.n4418 289.473
R4186 vss.n5347 vss.n4480 289.473
R4187 vss.n5288 vss.n4525 289.473
R4188 vss.n5221 vss.n4592 289.473
R4189 vss.n5173 vss.n4631 289.473
R4190 vss.n5106 vss.n4693 289.473
R4191 vss.n5047 vss.n4738 289.473
R4192 vss.n4980 vss.n4805 289.473
R4193 vss.n4932 vss.n4844 289.473
R4194 vss.n16735 vss.n16734 289.473
R4195 vss.n16832 vss.n16831 289.473
R4196 vss.n16965 vss.n16964 289.473
R4197 vss.n17066 vss.n17065 289.473
R4198 vss.n17201 vss.n17200 289.473
R4199 vss.n17322 vss.n17321 289.473
R4200 vss.n16012 vss.n16011 289.473
R4201 vss.n16112 vss.n16111 289.473
R4202 vss.n15284 vss.n15283 289.473
R4203 vss.n15351 vss.n15350 289.473
R4204 vss.n15485 vss.n15484 289.473
R4205 vss.n15588 vss.n15587 289.473
R4206 vss.n15721 vss.n15720 289.473
R4207 vss.n15812 vss.n15811 289.473
R4208 vss.n16432 vss.n16431 289.473
R4209 vss.n16535 vss.n16534 289.473
R4210 vss.n17600 vss.n17575 289.093
R4211 vss.n4210 vss.n4185 289.093
R4212 vss.n20296 vss.n17556 286.235
R4213 vss.n6906 vss.n4166 286.235
R4214 vss.n22627 vss.n22626 285.714
R4215 vss.n22552 vss.n22551 285.714
R4216 vss.n22419 vss.n22418 285.714
R4217 vss.n22344 vss.n22343 285.714
R4218 vss.n22211 vss.n22210 285.714
R4219 vss.n22136 vss.n22135 285.714
R4220 vss.n21555 vss.n21554 285.714
R4221 vss.n21480 vss.n21479 285.714
R4222 vss.n21347 vss.n21346 285.714
R4223 vss.n21272 vss.n21271 285.714
R4224 vss.n21139 vss.n21138 285.714
R4225 vss.n21064 vss.n21063 285.714
R4226 vss.n20931 vss.n20930 285.714
R4227 vss.n8790 vss.n8789 285.714
R4228 vss.n8715 vss.n8714 285.714
R4229 vss.n8582 vss.n8581 285.714
R4230 vss.n8507 vss.n8506 285.714
R4231 vss.n8374 vss.n8373 285.714
R4232 vss.n8299 vss.n8298 285.714
R4233 vss.n8166 vss.n8165 285.714
R4234 vss.n8091 vss.n8090 285.714
R4235 vss.n7958 vss.n7957 285.714
R4236 vss.n7883 vss.n7882 285.714
R4237 vss.n7749 vss.n7748 285.714
R4238 vss.n7674 vss.n7673 285.714
R4239 vss.n7541 vss.n7540 285.714
R4240 vss.t326 vss.t313 271.232
R4241 vss.t313 vss.t356 271.232
R4242 vss.t356 vss.t214 271.232
R4243 vss.t211 vss.t11 271.232
R4244 vss.t8 vss.t211 271.232
R4245 vss.t321 vss.t8 271.232
R4246 vss.t232 vss.t321 271.232
R4247 vss.t215 vss.t232 271.232
R4248 vss.t226 vss.t215 271.232
R4249 vss.t217 vss.t226 271.232
R4250 vss.t217 vss.t227 271.232
R4251 vss.t227 vss.t212 271.232
R4252 vss.t212 vss.t318 271.232
R4253 vss.t307 vss.t312 271.232
R4254 vss.t330 vss.t307 271.232
R4255 vss.t12 vss.t330 271.232
R4256 vss.t3 vss.t12 271.232
R4257 vss.t216 vss.t3 271.232
R4258 vss.t325 vss.t216 271.232
R4259 vss.t0 vss.t325 271.232
R4260 vss.n20256 vss.n20255 260.526
R4261 vss.n20187 vss.n20186 260.526
R4262 vss.n20136 vss.n20135 260.526
R4263 vss.n19227 vss.n19215 260.526
R4264 vss.n20009 vss.n20008 260.526
R4265 vss.n19940 vss.n19939 260.526
R4266 vss.n19889 vss.n19888 260.526
R4267 vss.n19434 vss.n19422 260.526
R4268 vss.n19762 vss.n19761 260.526
R4269 vss.n19693 vss.n19692 260.526
R4270 vss.n19642 vss.n19641 260.526
R4271 vss.n20329 vss.n20328 260.526
R4272 vss.n18990 vss.n18989 260.526
R4273 vss.n17720 vss.n17708 260.526
R4274 vss.n18863 vss.n18862 260.526
R4275 vss.n18794 vss.n18793 260.526
R4276 vss.n17869 vss.n17860 260.526
R4277 vss.n17933 vss.n17921 260.526
R4278 vss.n18622 vss.n18621 260.526
R4279 vss.n18553 vss.n18552 260.526
R4280 vss.n18082 vss.n18073 260.526
R4281 vss.n18146 vss.n18134 260.526
R4282 vss.n18381 vss.n18380 260.526
R4283 vss.n18312 vss.n18311 260.526
R4284 vss.n6866 vss.n6865 260.526
R4285 vss.n6797 vss.n6796 260.526
R4286 vss.n6746 vss.n6745 260.526
R4287 vss.n5837 vss.n5825 260.526
R4288 vss.n6619 vss.n6618 260.526
R4289 vss.n6550 vss.n6549 260.526
R4290 vss.n6499 vss.n6498 260.526
R4291 vss.n6044 vss.n6032 260.526
R4292 vss.n6372 vss.n6371 260.526
R4293 vss.n6303 vss.n6302 260.526
R4294 vss.n6252 vss.n6251 260.526
R4295 vss.n6939 vss.n6938 260.526
R4296 vss.n5600 vss.n5599 260.526
R4297 vss.n4330 vss.n4318 260.526
R4298 vss.n5473 vss.n5472 260.526
R4299 vss.n5404 vss.n5403 260.526
R4300 vss.n4479 vss.n4470 260.526
R4301 vss.n4543 vss.n4531 260.526
R4302 vss.n5232 vss.n5231 260.526
R4303 vss.n5163 vss.n5162 260.526
R4304 vss.n4692 vss.n4683 260.526
R4305 vss.n4756 vss.n4744 260.526
R4306 vss.n4991 vss.n4990 260.526
R4307 vss.n4922 vss.n4921 260.526
R4308 vss.n16720 vss.n16719 260.526
R4309 vss.n16845 vss.n16844 260.526
R4310 vss.n16950 vss.n16949 260.526
R4311 vss.n17079 vss.n17078 260.526
R4312 vss.n17186 vss.n17185 260.526
R4313 vss.n17281 vss.n17280 260.526
R4314 vss.n15889 vss.n15888 260.526
R4315 vss.n15997 vss.n15996 260.526
R4316 vss.n16125 vss.n16124 260.526
R4317 vss.n16233 vss.n16232 260.526
R4318 vss.n15269 vss.n15268 260.526
R4319 vss.n15365 vss.n15364 260.526
R4320 vss.n15470 vss.n15469 260.526
R4321 vss.n15601 vss.n15600 260.526
R4322 vss.n15706 vss.n15705 260.526
R4323 vss.n15829 vss.n15828 260.526
R4324 vss.n16312 vss.n16311 260.526
R4325 vss.n16417 vss.n16416 260.526
R4326 vss.n16548 vss.n16547 260.526
R4327 vss.n16653 vss.n16652 260.526
R4328 vss.n11812 vss.n11811 259.842
R4329 vss.n15001 vss.n15000 259.842
R4330 vss.n12399 vss.n12398 259.842
R4331 vss.n14709 vss.n14708 259.842
R4332 vss.n13446 vss.n13445 259.842
R4333 vss.n13021 vss.n13020 259.842
R4334 vss.n10578 vss.n10577 259.842
R4335 vss.n10735 vss.n10734 259.842
R4336 vss.n12031 vss.n12030 259.842
R4337 vss.n14573 vss.n14572 259.842
R4338 vss.n13633 vss.n13632 259.842
R4339 vss.n13685 vss.n13684 259.842
R4340 vss.n11382 vss.n11381 259.842
R4341 vss.n11368 vss.n11367 259.842
R4342 vss.n11311 vss.n11310 259.842
R4343 vss.n13959 vss.n13958 259.842
R4344 vss.n22747 vss.n22746 257.142
R4345 vss.n22642 vss.n22641 257.142
R4346 vss.n22539 vss.n22538 257.142
R4347 vss.n22434 vss.n22433 257.142
R4348 vss.n22331 vss.n22330 257.142
R4349 vss.n22226 vss.n22225 257.142
R4350 vss.n22123 vss.n22122 257.142
R4351 vss.n21570 vss.n21569 257.142
R4352 vss.n21467 vss.n21466 257.142
R4353 vss.n21362 vss.n21361 257.142
R4354 vss.n21259 vss.n21258 257.142
R4355 vss.n21154 vss.n21153 257.142
R4356 vss.n21051 vss.n21050 257.142
R4357 vss.n20946 vss.n20945 257.142
R4358 vss.n8910 vss.n8909 257.142
R4359 vss.n8805 vss.n8804 257.142
R4360 vss.n8702 vss.n8701 257.142
R4361 vss.n8597 vss.n8596 257.142
R4362 vss.n8494 vss.n8493 257.142
R4363 vss.n8389 vss.n8388 257.142
R4364 vss.n8286 vss.n8285 257.142
R4365 vss.n8181 vss.n8180 257.142
R4366 vss.n8078 vss.n8077 257.142
R4367 vss.n7973 vss.n7972 257.142
R4368 vss.n7870 vss.n7869 257.142
R4369 vss.n7764 vss.n7763 257.142
R4370 vss.n7661 vss.n7660 257.142
R4371 vss.n7556 vss.n7555 257.142
R4372 vss.n12226 vss.n12225 255.813
R4373 vss.n12020 vss.n12019 255.813
R4374 vss.n11256 vss.n11255 255.813
R4375 vss.n11196 vss.n11195 255.813
R4376 vss.n13913 vss.n13912 255.813
R4377 vss.n14051 vss.n14050 255.813
R4378 vss.n11746 vss.n11745 255.813
R4379 vss.n11073 vss.n11072 255.813
R4380 vss.n14740 vss.n14739 255.813
R4381 vss.n14681 vss.n14680 255.813
R4382 vss.n14468 vss.n14467 255.813
R4383 vss.n14250 vss.n14249 255.813
R4384 vss.n12855 vss.n12854 255.813
R4385 vss.n12913 vss.n12912 255.813
R4386 vss.n12655 vss.n12654 255.813
R4387 vss.n12500 vss.n12499 255.813
R4388 vss.n10244 vss.t311 245.323
R4389 vss.n10268 vss.t224 245.323
R4390 vss.n10288 vss.t355 245.323
R4391 vss.n10311 vss.t360 245.323
R4392 vss.n10329 vss.t223 245.323
R4393 vss.n10371 vss.t85 245.323
R4394 vss.n10403 vss.t319 245.323
R4395 vss.n10437 vss.t225 245.323
R4396 vss.n8938 vss.t308 245.323
R4397 vss.n8956 vss.t317 245.323
R4398 vss.n8993 vss.t86 245.323
R4399 vss.n9023 vss.t320 245.323
R4400 vss.n9054 vss.t329 245.323
R4401 vss.n9085 vss.t213 245.323
R4402 vss.n9104 vss.t324 245.323
R4403 vss.n9134 vss.t222 245.323
R4404 vss.n1647 vss.t67 235.962
R4405 vss.n1473 vss.t29 235.962
R4406 vss.n108 vss.t277 235.962
R4407 vss.n1385 vss.t291 235.962
R4408 vss.n20255 vss.n20254 231.578
R4409 vss.n20188 vss.n20187 231.578
R4410 vss.n20135 vss.n19160 231.578
R4411 vss.n20063 vss.n19215 231.578
R4412 vss.n20008 vss.n20007 231.578
R4413 vss.n19941 vss.n19940 231.578
R4414 vss.n19888 vss.n19367 231.578
R4415 vss.n19816 vss.n19422 231.578
R4416 vss.n19761 vss.n19760 231.578
R4417 vss.n19694 vss.n19693 231.578
R4418 vss.n19641 vss.n19574 231.578
R4419 vss.n20329 vss.n17601 231.578
R4420 vss.n18989 vss.n17653 231.578
R4421 vss.n18917 vss.n17708 231.578
R4422 vss.n18862 vss.n18861 231.578
R4423 vss.n18795 vss.n18794 231.578
R4424 vss.n18739 vss.n17869 231.578
R4425 vss.n18676 vss.n17921 231.578
R4426 vss.n18621 vss.n18620 231.578
R4427 vss.n18554 vss.n18553 231.578
R4428 vss.n18498 vss.n18082 231.578
R4429 vss.n18435 vss.n18134 231.578
R4430 vss.n18380 vss.n18379 231.578
R4431 vss.n18313 vss.n18312 231.578
R4432 vss.n6865 vss.n6864 231.578
R4433 vss.n6798 vss.n6797 231.578
R4434 vss.n6745 vss.n5770 231.578
R4435 vss.n6673 vss.n5825 231.578
R4436 vss.n6618 vss.n6617 231.578
R4437 vss.n6551 vss.n6550 231.578
R4438 vss.n6498 vss.n5977 231.578
R4439 vss.n6426 vss.n6032 231.578
R4440 vss.n6371 vss.n6370 231.578
R4441 vss.n6304 vss.n6303 231.578
R4442 vss.n6251 vss.n6184 231.578
R4443 vss.n6939 vss.n4211 231.578
R4444 vss.n5599 vss.n4263 231.578
R4445 vss.n5527 vss.n4318 231.578
R4446 vss.n5472 vss.n5471 231.578
R4447 vss.n5405 vss.n5404 231.578
R4448 vss.n5349 vss.n4479 231.578
R4449 vss.n5286 vss.n4531 231.578
R4450 vss.n5231 vss.n5230 231.578
R4451 vss.n5164 vss.n5163 231.578
R4452 vss.n5108 vss.n4692 231.578
R4453 vss.n5045 vss.n4744 231.578
R4454 vss.n4990 vss.n4989 231.578
R4455 vss.n4923 vss.n4922 231.578
R4456 vss.n16721 vss.n16720 231.578
R4457 vss.n16846 vss.n16845 231.578
R4458 vss.n16951 vss.n16950 231.578
R4459 vss.n17080 vss.n17079 231.578
R4460 vss.n17187 vss.n17186 231.578
R4461 vss.n17282 vss.n17281 231.578
R4462 vss.n15890 vss.n15889 231.578
R4463 vss.n15998 vss.n15997 231.578
R4464 vss.n16126 vss.n16125 231.578
R4465 vss.n16234 vss.n16233 231.578
R4466 vss.n15270 vss.n15269 231.578
R4467 vss.n15366 vss.n15365 231.578
R4468 vss.n15471 vss.n15470 231.578
R4469 vss.n15602 vss.n15601 231.578
R4470 vss.n15707 vss.n15706 231.578
R4471 vss.n15830 vss.n15829 231.578
R4472 vss.n16313 vss.n16312 231.578
R4473 vss.n16418 vss.n16417 231.578
R4474 vss.n16549 vss.n16548 231.578
R4475 vss.n16654 vss.n16653 231.578
R4476 vss.n22746 vss.n22745 228.571
R4477 vss.n22641 vss.n22640 228.571
R4478 vss.n22538 vss.n22537 228.571
R4479 vss.n22433 vss.n22432 228.571
R4480 vss.n22330 vss.n22329 228.571
R4481 vss.n22225 vss.n22224 228.571
R4482 vss.n22122 vss.n22121 228.571
R4483 vss.n21569 vss.n21568 228.571
R4484 vss.n21466 vss.n21465 228.571
R4485 vss.n21361 vss.n21360 228.571
R4486 vss.n21258 vss.n21257 228.571
R4487 vss.n21153 vss.n21152 228.571
R4488 vss.n21050 vss.n21049 228.571
R4489 vss.n20945 vss.n20944 228.571
R4490 vss.n8909 vss.n8908 228.571
R4491 vss.n8804 vss.n8803 228.571
R4492 vss.n8701 vss.n8700 228.571
R4493 vss.n8596 vss.n8595 228.571
R4494 vss.n8493 vss.n8492 228.571
R4495 vss.n8388 vss.n8387 228.571
R4496 vss.n8285 vss.n8284 228.571
R4497 vss.n8180 vss.n8179 228.571
R4498 vss.n8077 vss.n8076 228.571
R4499 vss.n7972 vss.n7971 228.571
R4500 vss.n7869 vss.n7868 228.571
R4501 vss.n7763 vss.n7762 228.571
R4502 vss.n7660 vss.n7659 228.571
R4503 vss.n7555 vss.n7554 228.571
R4504 vss.n11477 vss.n11476 225.196
R4505 vss.n11695 vss.n11694 225.196
R4506 vss.n13117 vss.n13116 225.196
R4507 vss.n13666 vss.n13665 225.196
R4508 vss.n14982 vss.n14981 225.196
R4509 vss.n13144 vss.n13143 225.196
R4510 vss.n12409 vss.n12408 225.196
R4511 vss.n10672 vss.n10671 225.196
R4512 vss.n12326 vss.n12325 225.196
R4513 vss.n11487 vss.n11486 225.196
R4514 vss.n13375 vss.n13374 225.196
R4515 vss.n13458 vss.n13457 225.196
R4516 vss.n13089 vss.n13088 225.196
R4517 vss.n10642 vss.n10641 225.196
R4518 vss.n12311 vss.n12310 225.196
R4519 vss.n10808 vss.n10807 225.196
R4520 vss.n14563 vss.n14562 225.196
R4521 vss.n14100 vss.n14099 225.196
R4522 vss.n13750 vss.n13749 225.196
R4523 vss.n11447 vss.n11446 225.196
R4524 vss.n11856 vss.n11855 225.196
R4525 vss.n10933 vss.n10932 225.196
R4526 vss.n13653 vss.n13652 225.196
R4527 vss.n14062 vss.n14061 225.196
R4528 vss.n20528 vss.n20527 223.931
R4529 vss.n20556 vss.n20555 223.931
R4530 vss.n20757 vss.n20756 223.931
R4531 vss.n20778 vss.n20777 223.931
R4532 vss.n7138 vss.n7137 223.931
R4533 vss.n7166 vss.n7165 223.931
R4534 vss.n7367 vss.n7366 223.931
R4535 vss.n7388 vss.n7387 223.931
R4536 vss.n1754 vss.n1753 223.931
R4537 vss.n1775 vss.n1774 223.931
R4538 vss.n1985 vss.n1982 223.931
R4539 vss.n2015 vss.n2012 223.931
R4540 vss.n2230 vss.n2227 223.931
R4541 vss.n2259 vss.n2256 223.931
R4542 vss.n2474 vss.n2471 223.931
R4543 vss.n2503 vss.n2500 223.931
R4544 vss.n2719 vss.n2716 223.931
R4545 vss.n2748 vss.n2745 223.931
R4546 vss.n2957 vss.n2954 223.931
R4547 vss.n2986 vss.n2983 223.931
R4548 vss.n3201 vss.n3198 223.931
R4549 vss.n3231 vss.n3228 223.931
R4550 vss.n15203 vss.n15202 223.931
R4551 vss.n15184 vss.n15183 223.931
R4552 vss.n215 vss.n214 223.931
R4553 vss.n236 vss.n235 223.931
R4554 vss.n446 vss.n443 223.931
R4555 vss.n476 vss.n473 223.931
R4556 vss.n691 vss.n688 223.931
R4557 vss.n720 vss.n717 223.931
R4558 vss.n935 vss.n932 223.931
R4559 vss.n964 vss.n961 223.931
R4560 vss.n1180 vss.n1177 223.931
R4561 vss.n1209 vss.n1206 223.931
R4562 vss.n23303 vss.n23300 223.931
R4563 vss.n23276 vss.n23273 223.931
R4564 vss.n23059 vss.n23056 223.931
R4565 vss.n23031 vss.n23028 223.931
R4566 vss.n1396 vss.n1395 223.931
R4567 vss.n22818 vss.n22817 223.931
R4568 vss.n9161 vss.t326 210.958
R4569 vss.n10186 vss.t0 210.958
R4570 vss.n10247 vss.n10241 210.07
R4571 vss.n10271 vss.n10266 210.07
R4572 vss.n10291 vss.n10285 210.07
R4573 vss.n10314 vss.n10308 210.07
R4574 vss.n10332 vss.n10326 210.07
R4575 vss.n10374 vss.n10368 210.07
R4576 vss.n10406 vss.n10400 210.07
R4577 vss.n10440 vss.n10434 210.07
R4578 vss.n8942 vss.n8941 210.07
R4579 vss.n8960 vss.n8959 210.07
R4580 vss.n8996 vss.n8990 210.07
R4581 vss.n9026 vss.n9020 210.07
R4582 vss.n9057 vss.n9051 210.07
R4583 vss.n9088 vss.n9082 210.07
R4584 vss.n9107 vss.n9101 210.07
R4585 vss.n9137 vss.n9131 210.07
R4586 vss.n12888 vss.n12886 208.588
R4587 vss.n12479 vss.n12477 208.588
R4588 vss.n9782 vss.n9779 204.423
R4589 vss.n19069 vss.n19060 202.631
R4590 vss.n19120 vss.n19108 202.631
R4591 vss.n20125 vss.n20124 202.631
R4592 vss.n20065 vss.n20064 202.631
R4593 vss.n19276 vss.n19267 202.631
R4594 vss.n19327 vss.n19315 202.631
R4595 vss.n19878 vss.n19877 202.631
R4596 vss.n19818 vss.n19817 202.631
R4597 vss.n19483 vss.n19474 202.631
R4598 vss.n19534 vss.n19522 202.631
R4599 vss.n19631 vss.n19630 202.631
R4600 vss.n20335 vss.n20334 202.631
R4601 vss.n18979 vss.n18978 202.631
R4602 vss.n18919 vss.n18918 202.631
R4603 vss.n17769 vss.n17760 202.631
R4604 vss.n17820 vss.n17808 202.631
R4605 vss.n18738 vss.n18737 202.631
R4606 vss.n18678 vss.n18677 202.631
R4607 vss.n17982 vss.n17973 202.631
R4608 vss.n18033 vss.n18021 202.631
R4609 vss.n18497 vss.n18496 202.631
R4610 vss.n18437 vss.n18436 202.631
R4611 vss.n18195 vss.n18186 202.631
R4612 vss.n18246 vss.n18234 202.631
R4613 vss.n5679 vss.n5670 202.631
R4614 vss.n5730 vss.n5718 202.631
R4615 vss.n6735 vss.n6734 202.631
R4616 vss.n6675 vss.n6674 202.631
R4617 vss.n5886 vss.n5877 202.631
R4618 vss.n5937 vss.n5925 202.631
R4619 vss.n6488 vss.n6487 202.631
R4620 vss.n6428 vss.n6427 202.631
R4621 vss.n6093 vss.n6084 202.631
R4622 vss.n6144 vss.n6132 202.631
R4623 vss.n6241 vss.n6240 202.631
R4624 vss.n6945 vss.n6944 202.631
R4625 vss.n5589 vss.n5588 202.631
R4626 vss.n5529 vss.n5528 202.631
R4627 vss.n4379 vss.n4370 202.631
R4628 vss.n4430 vss.n4418 202.631
R4629 vss.n5348 vss.n5347 202.631
R4630 vss.n5288 vss.n5287 202.631
R4631 vss.n4592 vss.n4583 202.631
R4632 vss.n4643 vss.n4631 202.631
R4633 vss.n5107 vss.n5106 202.631
R4634 vss.n5047 vss.n5046 202.631
R4635 vss.n4805 vss.n4796 202.631
R4636 vss.n4856 vss.n4844 202.631
R4637 vss.n16734 vss.n16733 202.631
R4638 vss.n16831 vss.n16830 202.631
R4639 vss.n16964 vss.n16963 202.631
R4640 vss.n17065 vss.n17064 202.631
R4641 vss.n17200 vss.n17199 202.631
R4642 vss.n17321 vss.n17320 202.631
R4643 vss.n16011 vss.n16010 202.631
R4644 vss.n16111 vss.n16110 202.631
R4645 vss.n15283 vss.n15282 202.631
R4646 vss.n15350 vss.n15349 202.631
R4647 vss.n15484 vss.n15483 202.631
R4648 vss.n15587 vss.n15586 202.631
R4649 vss.n15720 vss.n15719 202.631
R4650 vss.n15811 vss.n15810 202.631
R4651 vss.n16431 vss.n16430 202.631
R4652 vss.n16534 vss.n16533 202.631
R4653 vss.n20409 vss.n20408 200.702
R4654 vss.n7019 vss.n7018 200.702
R4655 vss.n22628 vss.n22627 200
R4656 vss.n22553 vss.n22552 200
R4657 vss.n22420 vss.n22419 200
R4658 vss.n22345 vss.n22344 200
R4659 vss.n22212 vss.n22211 200
R4660 vss.n22137 vss.n22136 200
R4661 vss.n21556 vss.n21555 200
R4662 vss.n21481 vss.n21480 200
R4663 vss.n21348 vss.n21347 200
R4664 vss.n21273 vss.n21272 200
R4665 vss.n21140 vss.n21139 200
R4666 vss.n21065 vss.n21064 200
R4667 vss.n20932 vss.n20931 200
R4668 vss.n8791 vss.n8790 200
R4669 vss.n8716 vss.n8715 200
R4670 vss.n8583 vss.n8582 200
R4671 vss.n8508 vss.n8507 200
R4672 vss.n8375 vss.n8374 200
R4673 vss.n8300 vss.n8299 200
R4674 vss.n8167 vss.n8166 200
R4675 vss.n8092 vss.n8091 200
R4676 vss.n7959 vss.n7958 200
R4677 vss.n7884 vss.n7883 200
R4678 vss.n7750 vss.n7749 200
R4679 vss.n7675 vss.n7674 200
R4680 vss.n7542 vss.n7541 200
R4681 vss.n9239 vss.n9238 199.152
R4682 vss.n1583 vss.t55 194.321
R4683 vss.n1540 vss.t43 194.321
R4684 vss.n44 vss.t265 194.321
R4685 vss.n1320 vss.t299 194.321
R4686 vss.n9179 vss.n9167 191.246
R4687 vss.n9190 vss.n9165 191.246
R4688 vss.n11549 vss.n11548 190.551
R4689 vss.n11518 vss.n11517 190.551
R4690 vss.n12988 vss.n12987 190.551
R4691 vss.n12978 vss.n12977 190.551
R4692 vss.n12947 vss.n12946 190.551
R4693 vss.n13158 vss.n13157 190.551
R4694 vss.n12388 vss.n12387 190.551
R4695 vss.n12361 vss.n12360 190.551
R4696 vss.n10692 vss.n10691 190.551
R4697 vss.n10702 vss.n10701 190.551
R4698 vss.n13415 vss.n13414 190.551
R4699 vss.n13494 vss.n13493 190.551
R4700 vss.n13074 vss.n13073 190.551
R4701 vss.n10627 vss.n10626 190.551
R4702 vss.n10787 vss.n10786 190.551
R4703 vss.n12295 vss.n12294 190.551
R4704 vss.n14159 vss.n14158 190.551
R4705 vss.n14116 vss.n14115 190.551
R4706 vss.n13735 vss.n13734 190.551
R4707 vss.n11432 vss.n11431 190.551
R4708 vss.n11872 vss.n11871 190.551
R4709 vss.n11908 vss.n11907 190.551
R4710 vss.n13782 vss.n13781 190.551
R4711 vss.n13793 vss.n13792 190.551
R4712 vss.n21745 vss.n21744 185
R4713 vss.n21727 vss.n21718 185
R4714 vss.n21732 vss.n21716 185
R4715 vss.n21741 vss.n21713 185
R4716 vss.n21729 vss.n21728 185
R4717 vss.n21731 vss.n21730 185
R4718 vss.n21733 vss.n21714 185
R4719 vss.n21796 vss.n21662 185
R4720 vss.n21796 vss.n21660 185
R4721 vss.n21796 vss.n21659 185
R4722 vss.n21797 vss.n21796 185
R4723 vss.n3694 vss.n3693 185
R4724 vss.n3676 vss.n3667 185
R4725 vss.n3681 vss.n3665 185
R4726 vss.n3690 vss.n3662 185
R4727 vss.n3678 vss.n3677 185
R4728 vss.n3680 vss.n3679 185
R4729 vss.n3682 vss.n3663 185
R4730 vss.n3745 vss.n3611 185
R4731 vss.n3745 vss.n3609 185
R4732 vss.n3745 vss.n3608 185
R4733 vss.n3746 vss.n3745 185
R4734 vss.n20532 vss.n20525 174.534
R4735 vss.n20559 vss.n20550 174.534
R4736 vss.n20761 vss.n20754 174.534
R4737 vss.n20781 vss.n20772 174.534
R4738 vss.n7142 vss.n7135 174.534
R4739 vss.n7169 vss.n7160 174.534
R4740 vss.n7371 vss.n7364 174.534
R4741 vss.n7391 vss.n7382 174.534
R4742 vss.n1758 vss.n1751 174.534
R4743 vss.n1778 vss.n1769 174.534
R4744 vss.n1989 vss.n1980 174.534
R4745 vss.n2018 vss.n2007 174.534
R4746 vss.n2234 vss.n2225 174.534
R4747 vss.n2262 vss.n2251 174.534
R4748 vss.n2478 vss.n2469 174.534
R4749 vss.n2506 vss.n2495 174.534
R4750 vss.n2723 vss.n2714 174.534
R4751 vss.n2751 vss.n2740 174.534
R4752 vss.n2961 vss.n2952 174.534
R4753 vss.n2989 vss.n2978 174.534
R4754 vss.n3205 vss.n3196 174.534
R4755 vss.n3234 vss.n3223 174.534
R4756 vss.n15207 vss.n15200 174.534
R4757 vss.n15187 vss.n15178 174.534
R4758 vss.n219 vss.n212 174.534
R4759 vss.n239 vss.n230 174.534
R4760 vss.n450 vss.n441 174.534
R4761 vss.n479 vss.n468 174.534
R4762 vss.n695 vss.n686 174.534
R4763 vss.n723 vss.n712 174.534
R4764 vss.n939 vss.n930 174.534
R4765 vss.n967 vss.n956 174.534
R4766 vss.n1184 vss.n1175 174.534
R4767 vss.n1212 vss.n1201 174.534
R4768 vss.n23307 vss.n23298 174.534
R4769 vss.n23279 vss.n23268 174.534
R4770 vss.n23063 vss.n23054 174.534
R4771 vss.n23034 vss.n23023 174.534
R4772 vss.n1400 vss.n1393 174.534
R4773 vss.n22821 vss.n22812 174.534
R4774 vss.n20266 vss.n19050 173.684
R4775 vss.n20176 vss.n19121 173.684
R4776 vss.n20137 vss.n19151 173.684
R4777 vss.n20054 vss.n20053 173.684
R4778 vss.n20019 vss.n19258 173.684
R4779 vss.n19929 vss.n19328 173.684
R4780 vss.n19890 vss.n19358 173.684
R4781 vss.n19807 vss.n19806 173.684
R4782 vss.n19772 vss.n19465 173.684
R4783 vss.n19682 vss.n19535 173.684
R4784 vss.n19643 vss.n19565 173.684
R4785 vss.n20327 vss.n17603 173.684
R4786 vss.n18991 vss.n17644 173.684
R4787 vss.n18908 vss.n18907 173.684
R4788 vss.n18873 vss.n17751 173.684
R4789 vss.n18783 vss.n17821 173.684
R4790 vss.n18749 vss.n18748 173.684
R4791 vss.n18667 vss.n18666 173.684
R4792 vss.n18632 vss.n17964 173.684
R4793 vss.n18542 vss.n18034 173.684
R4794 vss.n18508 vss.n18507 173.684
R4795 vss.n18426 vss.n18425 173.684
R4796 vss.n18391 vss.n18177 173.684
R4797 vss.n18301 vss.n18247 173.684
R4798 vss.n6876 vss.n5660 173.684
R4799 vss.n6786 vss.n5731 173.684
R4800 vss.n6747 vss.n5761 173.684
R4801 vss.n6664 vss.n6663 173.684
R4802 vss.n6629 vss.n5868 173.684
R4803 vss.n6539 vss.n5938 173.684
R4804 vss.n6500 vss.n5968 173.684
R4805 vss.n6417 vss.n6416 173.684
R4806 vss.n6382 vss.n6075 173.684
R4807 vss.n6292 vss.n6145 173.684
R4808 vss.n6253 vss.n6175 173.684
R4809 vss.n6937 vss.n4213 173.684
R4810 vss.n5601 vss.n4254 173.684
R4811 vss.n5518 vss.n5517 173.684
R4812 vss.n5483 vss.n4361 173.684
R4813 vss.n5393 vss.n4431 173.684
R4814 vss.n5359 vss.n5358 173.684
R4815 vss.n5277 vss.n5276 173.684
R4816 vss.n5242 vss.n4574 173.684
R4817 vss.n5152 vss.n4644 173.684
R4818 vss.n5118 vss.n5117 173.684
R4819 vss.n5036 vss.n5035 173.684
R4820 vss.n5001 vss.n4787 173.684
R4821 vss.n4911 vss.n4857 173.684
R4822 vss.n16707 vss.n16706 173.684
R4823 vss.n16858 vss.n16857 173.684
R4824 vss.n16937 vss.n16936 173.684
R4825 vss.n17094 vss.n17093 173.684
R4826 vss.n17173 vss.n17172 173.684
R4827 vss.n17311 vss.n17310 173.684
R4828 vss.n15904 vss.n15903 173.684
R4829 vss.n15984 vss.n15983 173.684
R4830 vss.n16140 vss.n16139 173.684
R4831 vss.n16220 vss.n16219 173.684
R4832 vss.n15256 vss.n15255 173.684
R4833 vss.n15380 vss.n15379 173.684
R4834 vss.n15457 vss.n15456 173.684
R4835 vss.n15616 vss.n15615 173.684
R4836 vss.n15693 vss.n15692 173.684
R4837 vss.n15844 vss.n15843 173.684
R4838 vss.n16327 vss.n16326 173.684
R4839 vss.n16404 vss.n16403 173.684
R4840 vss.n16563 vss.n16562 173.684
R4841 vss.n16640 vss.n16639 173.684
R4842 vss.n14326 vss.n14325 172.549
R4843 vss.n13899 vss.n13898 172.549
R4844 vss.n14457 vss.n14456 172.549
R4845 vss.n14427 vss.n14426 172.549
R4846 vss.n14000 vss.n13999 172.549
R4847 vss.n11592 vss.n11591 172.549
R4848 vss.n11735 vss.n11734 172.549
R4849 vss.n11143 vss.n11142 172.549
R4850 vss.n12454 vss.n12453 172.549
R4851 vss.n12616 vss.n12615 172.549
R4852 vss.n12155 vss.n12154 172.549
R4853 vss.n12212 vss.n12211 172.549
R4854 vss.n14639 vss.n14638 172.549
R4855 vss.n13561 vss.n13560 172.549
R4856 vss.n15032 vss.n15031 172.549
R4857 vss.n10477 vss.n10476 172.549
R4858 vss.n13315 vss.n13314 172.549
R4859 vss.n14752 vss.n14751 172.549
R4860 vss.n14919 vss.n14918 172.549
R4861 vss.n14947 vss.n14946 172.549
R4862 vss.n10845 vss.n10844 172.549
R4863 vss.n10889 vss.n10888 172.549
R4864 vss.n11245 vss.n11244 172.549
R4865 vss.n11210 vss.n11209 172.549
R4866 vss.n22731 vss.n22730 171.428
R4867 vss.n22654 vss.n22653 171.428
R4868 vss.n22523 vss.n22522 171.428
R4869 vss.n22446 vss.n22445 171.428
R4870 vss.n22315 vss.n22314 171.428
R4871 vss.n22238 vss.n22237 171.428
R4872 vss.n22107 vss.n22106 171.428
R4873 vss.n17403 vss.n17402 171.428
R4874 vss.n21451 vss.n21450 171.428
R4875 vss.n21374 vss.n21373 171.428
R4876 vss.n21243 vss.n21242 171.428
R4877 vss.n21166 vss.n21165 171.428
R4878 vss.n21035 vss.n21034 171.428
R4879 vss.n20958 vss.n20957 171.428
R4880 vss.n8894 vss.n8893 171.428
R4881 vss.n8817 vss.n8816 171.428
R4882 vss.n8686 vss.n8685 171.428
R4883 vss.n8609 vss.n8608 171.428
R4884 vss.n8478 vss.n8477 171.428
R4885 vss.n8401 vss.n8400 171.428
R4886 vss.n8270 vss.n8269 171.428
R4887 vss.n8193 vss.n8192 171.428
R4888 vss.n8062 vss.n8061 171.428
R4889 vss.n7985 vss.n7984 171.428
R4890 vss.n7854 vss.n7853 171.428
R4891 vss.n7776 vss.n7775 171.428
R4892 vss.n7645 vss.n7644 171.428
R4893 vss.n7568 vss.n7567 171.428
R4894 vss.n20648 vss.t235 166.561
R4895 vss.n20666 vss.t233 166.561
R4896 vss.n7258 vss.t45 166.561
R4897 vss.n7276 vss.t47 166.561
R4898 vss.n2602 vss.t81 166.561
R4899 vss.n2621 vss.t59 166.561
R4900 vss.n1063 vss.t283 166.561
R4901 vss.n1082 vss.t259 166.561
R4902 vss.n12070 vss.n12069 153.488
R4903 vss.n10799 vss.n10798 153.488
R4904 vss.n10962 vss.n10961 153.488
R4905 vss.n11002 vss.n11001 153.488
R4906 vss.n13852 vss.n13851 153.488
R4907 vss.n14073 vss.n14072 153.488
R4908 vss.n11719 vss.n11718 153.488
R4909 vss.n11063 vss.n11062 153.488
R4910 vss.n13350 vss.n13349 153.488
R4911 vss.n14695 vss.n14694 153.488
R4912 vss.n14188 vss.n14187 153.488
R4913 vss.n14230 vss.n14229 153.488
R4914 vss.n12870 vss.n12869 153.488
R4915 vss.n12919 vss.n12918 153.488
R4916 vss.n12465 vss.n12464 153.488
R4917 vss.n12506 vss.n12505 153.488
R4918 vss.n10272 vss.n10271 148.249
R4919 vss.n8961 vss.n8960 148.246
R4920 vss.n10315 vss.n10314 148.216
R4921 vss.n8943 vss.n8942 148.17
R4922 vss.n10253 vss.n10252 148.17
R4923 vss.n10248 vss.n10247 147.952
R4924 vss.n10292 vss.n10291 147.952
R4925 vss.n10333 vss.n10332 147.813
R4926 vss.n10375 vss.n10374 147.587
R4927 vss.n20244 vss.n20243 144.736
R4928 vss.n20199 vss.n20198 144.736
R4929 vss.n19179 vss.n19170 144.736
R4930 vss.n20076 vss.n20075 144.736
R4931 vss.n19997 vss.n19996 144.736
R4932 vss.n19952 vss.n19951 144.736
R4933 vss.n19386 vss.n19377 144.736
R4934 vss.n19829 vss.n19828 144.736
R4935 vss.n19750 vss.n19749 144.736
R4936 vss.n19705 vss.n19704 144.736
R4937 vss.n19600 vss.n19584 144.736
R4938 vss.n20341 vss.n20340 144.736
R4939 vss.n17672 vss.n17663 144.736
R4940 vss.n18930 vss.n18929 144.736
R4941 vss.n18851 vss.n18850 144.736
R4942 vss.n18806 vss.n18805 144.736
R4943 vss.n18727 vss.n18726 144.736
R4944 vss.n18689 vss.n18688 144.736
R4945 vss.n18610 vss.n18609 144.736
R4946 vss.n18565 vss.n18564 144.736
R4947 vss.n18486 vss.n18485 144.736
R4948 vss.n18448 vss.n18447 144.736
R4949 vss.n18369 vss.n18368 144.736
R4950 vss.n18324 vss.n18323 144.736
R4951 vss.n6854 vss.n6853 144.736
R4952 vss.n6809 vss.n6808 144.736
R4953 vss.n5789 vss.n5780 144.736
R4954 vss.n6686 vss.n6685 144.736
R4955 vss.n6607 vss.n6606 144.736
R4956 vss.n6562 vss.n6561 144.736
R4957 vss.n5996 vss.n5987 144.736
R4958 vss.n6439 vss.n6438 144.736
R4959 vss.n6360 vss.n6359 144.736
R4960 vss.n6315 vss.n6314 144.736
R4961 vss.n6210 vss.n6194 144.736
R4962 vss.n6951 vss.n6950 144.736
R4963 vss.n4282 vss.n4273 144.736
R4964 vss.n5540 vss.n5539 144.736
R4965 vss.n5461 vss.n5460 144.736
R4966 vss.n5416 vss.n5415 144.736
R4967 vss.n5337 vss.n5336 144.736
R4968 vss.n5299 vss.n5298 144.736
R4969 vss.n5220 vss.n5219 144.736
R4970 vss.n5175 vss.n5174 144.736
R4971 vss.n5096 vss.n5095 144.736
R4972 vss.n5058 vss.n5057 144.736
R4973 vss.n4979 vss.n4978 144.736
R4974 vss.n4934 vss.n4933 144.736
R4975 vss.n16748 vss.n16747 144.736
R4976 vss.n16817 vss.n16816 144.736
R4977 vss.n16978 vss.n16977 144.736
R4978 vss.n17051 vss.n17050 144.736
R4979 vss.n17214 vss.n17213 144.736
R4980 vss.n17302 vss.n17301 144.736
R4981 vss.n16024 vss.n16023 144.736
R4982 vss.n16096 vss.n16095 144.736
R4983 vss.n15297 vss.n15296 144.736
R4984 vss.n15336 vss.n15335 144.736
R4985 vss.n15498 vss.n15497 144.736
R4986 vss.n15573 vss.n15572 144.736
R4987 vss.n15734 vss.n15733 144.736
R4988 vss.n15801 vss.n15800 144.736
R4989 vss.n16445 vss.n16444 144.736
R4990 vss.n16520 vss.n16519 144.736
R4991 vss.n9090 vss.n9088 144.668
R4992 vss.n9028 vss.n9026 144.257
R4993 vss.n10441 vss.n10440 143.898
R4994 vss.n8998 vss.n8996 143.704
R4995 vss.n10407 vss.n10406 143.434
R4996 vss.n9059 vss.n9057 143.371
R4997 vss.n9110 vss.n9107 143.006
R4998 vss.n22614 vss.n22613 142.857
R4999 vss.n22567 vss.n22566 142.857
R5000 vss.n22406 vss.n22405 142.857
R5001 vss.n22359 vss.n22358 142.857
R5002 vss.n22198 vss.n22197 142.857
R5003 vss.n22151 vss.n22150 142.857
R5004 vss.n21542 vss.n21541 142.857
R5005 vss.n21495 vss.n21494 142.857
R5006 vss.n21334 vss.n21333 142.857
R5007 vss.n21287 vss.n21286 142.857
R5008 vss.n21126 vss.n21125 142.857
R5009 vss.n21079 vss.n21078 142.857
R5010 vss.n20918 vss.n20917 142.857
R5011 vss.n8777 vss.n8776 142.857
R5012 vss.n8730 vss.n8729 142.857
R5013 vss.n8569 vss.n8568 142.857
R5014 vss.n8522 vss.n8521 142.857
R5015 vss.n8361 vss.n8360 142.857
R5016 vss.n8314 vss.n8313 142.857
R5017 vss.n8153 vss.n8152 142.857
R5018 vss.n8106 vss.n8105 142.857
R5019 vss.n7945 vss.n7944 142.857
R5020 vss.n7898 vss.n7897 142.857
R5021 vss.n7736 vss.n7735 142.857
R5022 vss.n7689 vss.n7688 142.857
R5023 vss.n7528 vss.n7527 142.857
R5024 vss.n9139 vss.n9137 141.54
R5025 vss.n2342 vss.t73 138.801
R5026 vss.n2875 vss.t23 138.801
R5027 vss.n803 vss.t249 138.801
R5028 vss.n23386 vss.t297 138.801
R5029 vss.n21726 vss.n21719 136.669
R5030 vss.n3675 vss.n3668 136.669
R5031 vss.n21773 vss.t196 135.48
R5032 vss.n3722 vss.t112 135.48
R5033 vss.n21998 vss.t143 135.478
R5034 vss.n3947 vss.t121 135.478
R5035 vss.n21998 vss.t140 135.478
R5036 vss.n3947 vss.t149 135.478
R5037 vss.n21773 vss.t192 135.427
R5038 vss.n3722 vss.t183 135.427
R5039 vss.n9185 vss.n9184 127.668
R5040 vss.n21744 vss.n21708 118.524
R5041 vss.n3693 vss.n3657 118.524
R5042 vss.n0 vss.n1 159.639
R5043 vss.n20268 vss.n19040 115.789
R5044 vss.n20174 vss.n19127 115.789
R5045 vss.n20145 vss.n20144 115.789
R5046 vss.n20042 vss.n19228 115.789
R5047 vss.n20021 vss.n19257 115.789
R5048 vss.n19927 vss.n19334 115.789
R5049 vss.n19898 vss.n19897 115.789
R5050 vss.n19795 vss.n19435 115.789
R5051 vss.n19774 vss.n19464 115.789
R5052 vss.n19680 vss.n19541 115.789
R5053 vss.n19651 vss.n19650 115.789
R5054 vss.n20322 vss.n20321 115.789
R5055 vss.n20298 vss.n0 115.789
R5056 vss.n2 vss.n19029 115.789
R5057 vss.n18999 vss.n18998 115.789
R5058 vss.n18896 vss.n17721 115.789
R5059 vss.n18875 vss.n17750 115.789
R5060 vss.n18781 vss.n17827 115.789
R5061 vss.n18760 vss.n17851 115.789
R5062 vss.n18655 vss.n17934 115.789
R5063 vss.n18634 vss.n17963 115.789
R5064 vss.n18540 vss.n18040 115.789
R5065 vss.n18519 vss.n18064 115.789
R5066 vss.n18414 vss.n18147 115.789
R5067 vss.n18393 vss.n18176 115.789
R5068 vss.n18299 vss.n18253 115.789
R5069 vss.n2 vss.n3 159.639
R5070 vss.n4 vss.n5 159.639
R5071 vss.n6878 vss.n5650 115.789
R5072 vss.n6784 vss.n5737 115.789
R5073 vss.n6755 vss.n6754 115.789
R5074 vss.n6652 vss.n5838 115.789
R5075 vss.n6631 vss.n5867 115.789
R5076 vss.n6537 vss.n5944 115.789
R5077 vss.n6508 vss.n6507 115.789
R5078 vss.n6405 vss.n6045 115.789
R5079 vss.n6384 vss.n6074 115.789
R5080 vss.n6290 vss.n6151 115.789
R5081 vss.n6261 vss.n6260 115.789
R5082 vss.n6932 vss.n6931 115.789
R5083 vss.n6908 vss.n4 115.789
R5084 vss.n6 vss.n5639 115.789
R5085 vss.n5609 vss.n5608 115.789
R5086 vss.n5506 vss.n4331 115.789
R5087 vss.n5485 vss.n4360 115.789
R5088 vss.n5391 vss.n4437 115.789
R5089 vss.n5370 vss.n4461 115.789
R5090 vss.n5265 vss.n4544 115.789
R5091 vss.n5244 vss.n4573 115.789
R5092 vss.n5150 vss.n4650 115.789
R5093 vss.n5129 vss.n4674 115.789
R5094 vss.n5024 vss.n4757 115.789
R5095 vss.n5003 vss.n4786 115.789
R5096 vss.n4909 vss.n4863 115.789
R5097 vss.n6 vss.n7 159.639
R5098 vss.n16693 vss.n16692 115.789
R5099 vss.n16872 vss.n16871 115.789
R5100 vss.n16923 vss.n16922 115.789
R5101 vss.n17108 vss.n17107 115.789
R5102 vss.n17159 vss.n17158 115.789
R5103 vss.n17270 vss.n17269 115.789
R5104 vss.n15878 vss.n15877 115.789
R5105 vss.n15918 vss.n15917 115.789
R5106 vss.n15970 vss.n15969 115.789
R5107 vss.n16154 vss.n16153 115.789
R5108 vss.n16206 vss.n16205 115.789
R5109 vss.n16279 vss.n16278 115.789
R5110 vss.n15394 vss.n15393 115.789
R5111 vss.n15443 vss.n15442 115.789
R5112 vss.n15630 vss.n15629 115.789
R5113 vss.n15679 vss.n15678 115.789
R5114 vss.n15858 vss.n15857 115.789
R5115 vss.n16299 vss.n16298 115.789
R5116 vss.n16341 vss.n16340 115.789
R5117 vss.n16390 vss.n16389 115.789
R5118 vss.n16577 vss.n16576 115.789
R5119 vss.n16626 vss.n16625 115.789
R5120 vss.n14358 vss.n14357 115.032
R5121 vss.n13864 vss.n13863 115.032
R5122 vss.n14492 vss.n14491 115.032
R5123 vss.n14399 vss.n14398 115.032
R5124 vss.n13979 vss.n13978 115.032
R5125 vss.n11574 vss.n11573 115.032
R5126 vss.n11761 vss.n11760 115.032
R5127 vss.n11051 vss.n11050 115.032
R5128 vss.n12426 vss.n12425 115.032
R5129 vss.n12599 vss.n12598 115.032
R5130 vss.n12584 vss.n12583 115.032
R5131 vss.n12080 vss.n12079 115.032
R5132 vss.n14662 vss.n14661 115.032
R5133 vss.n13581 vss.n13580 115.032
R5134 vss.n15016 vss.n15015 115.032
R5135 vss.n10507 vss.n10506 115.032
R5136 vss.n13299 vss.n13298 115.032
R5137 vss.n13340 vss.n13339 115.032
R5138 vss.n13241 vss.n13240 115.032
R5139 vss.n14962 vss.n14961 115.032
R5140 vss.n10825 vss.n10824 115.032
R5141 vss.n10899 vss.n10898 115.032
R5142 vss.n10952 vss.n10951 115.032
R5143 vss.n11012 vss.n11011 115.032
R5144 vss.n22717 vss.n22716 114.285
R5145 vss.n22668 vss.n22667 114.285
R5146 vss.n22509 vss.n22508 114.285
R5147 vss.n22460 vss.n22459 114.285
R5148 vss.n22301 vss.n22300 114.285
R5149 vss.n22252 vss.n22251 114.285
R5150 vss.n22093 vss.n22092 114.285
R5151 vss.n21584 vss.n21583 114.285
R5152 vss.n21437 vss.n21436 114.285
R5153 vss.n21388 vss.n21387 114.285
R5154 vss.n21229 vss.n21228 114.285
R5155 vss.n21180 vss.n21179 114.285
R5156 vss.n21021 vss.n21020 114.285
R5157 vss.n20972 vss.n20971 114.285
R5158 vss.n8880 vss.n8879 114.285
R5159 vss.n8831 vss.n8830 114.285
R5160 vss.n8672 vss.n8671 114.285
R5161 vss.n8623 vss.n8622 114.285
R5162 vss.n8464 vss.n8463 114.285
R5163 vss.n8415 vss.n8414 114.285
R5164 vss.n8256 vss.n8255 114.285
R5165 vss.n8207 vss.n8206 114.285
R5166 vss.n8048 vss.n8047 114.285
R5167 vss.n7999 vss.n7998 114.285
R5168 vss.n7839 vss.n7838 114.285
R5169 vss.n7790 vss.n7789 114.285
R5170 vss.n7631 vss.n7630 114.285
R5171 vss.n7582 vss.n7581 114.285
R5172 vss.n17524 vss.n17521 111.041
R5173 vss.n17511 vss.n17509 111.041
R5174 vss.n4134 vss.n4131 111.041
R5175 vss.n4121 vss.n4119 111.041
R5176 vss.n1646 vss.n1643 111.041
R5177 vss.n1634 vss.n1631 111.041
R5178 vss.n2081 vss.t25 111.041
R5179 vss.n1619 vss.n1616 111.041
R5180 vss.n1607 vss.n1604 111.041
R5181 vss.n1594 vss.n1591 111.041
R5182 vss.n1582 vss.n1579 111.041
R5183 vss.n1569 vss.n1566 111.041
R5184 vss.n1556 vss.n1553 111.041
R5185 vss.n1539 vss.n1533 111.041
R5186 vss.n1524 vss.n1521 111.041
R5187 vss.n1511 vss.n1508 111.041
R5188 vss.n1499 vss.n1496 111.041
R5189 vss.n3136 vss.t69 111.041
R5190 vss.n1484 vss.n1481 111.041
R5191 vss.n1472 vss.n1469 111.041
R5192 vss.n107 vss.n104 111.041
R5193 vss.n95 vss.n92 111.041
R5194 vss.n542 vss.t293 111.041
R5195 vss.n80 vss.n77 111.041
R5196 vss.n68 vss.n65 111.041
R5197 vss.n55 vss.n52 111.041
R5198 vss.n43 vss.n40 111.041
R5199 vss.n30 vss.n27 111.041
R5200 vss.n17 vss.n14 111.041
R5201 vss.n1319 vss.n1316 111.041
R5202 vss.n1331 vss.n1328 111.041
R5203 vss.n1345 vss.n1342 111.041
R5204 vss.n1357 vss.n1354 111.041
R5205 vss.n23126 vss.t253 111.041
R5206 vss.n1372 vss.n1369 111.041
R5207 vss.n1384 vss.n1381 111.041
R5208 vss.n9179 vss.n9178 110.305
R5209 vss.n9191 vss.n9190 110.305
R5210 vss.n20437 vss.n20436 105.765
R5211 vss.n20888 vss.n20887 105.765
R5212 vss.n7047 vss.n7046 105.765
R5213 vss.n7498 vss.n7497 105.765
R5214 vss.n1677 vss.n1676 105.765
R5215 vss.n15151 vss.n15150 105.765
R5216 vss.n138 vss.n137 105.765
R5217 vss.n22785 vss.n22784 105.765
R5218 vss.n9185 vss.t9 105.119
R5219 vss.n19020 vss.n17628 104.41
R5220 vss.n19016 vss.n17635 104.41
R5221 vss.n19012 vss.n17635 104.41
R5222 vss.n19008 vss.n17639 104.41
R5223 vss.n18996 vss.n17643 104.41
R5224 vss.n18992 vss.n17652 104.41
R5225 vss.n18980 vss.n17654 104.41
R5226 vss.n18976 vss.n17664 104.41
R5227 vss.n18969 vss.n17671 104.41
R5228 vss.n18957 vss.n17674 104.41
R5229 vss.n18942 vss.n17690 104.41
R5230 vss.n18932 vss.n17696 104.41
R5231 vss.n18928 vss.n17703 104.41
R5232 vss.n18916 vss.n17707 104.41
R5233 vss.n18909 vss.n17718 104.41
R5234 vss.n18905 vss.n17722 104.41
R5235 vss.n18893 vss.n17726 104.41
R5236 vss.n18888 vss.n17736 104.41
R5237 vss.n18888 vss.n17737 104.41
R5238 vss.n17748 vss.n17740 104.41
R5239 vss.n18876 vss.n17746 104.41
R5240 vss.n18864 vss.n17752 104.41
R5241 vss.n18860 vss.n17761 104.41
R5242 vss.n18853 vss.n17768 104.41
R5243 vss.n18841 vss.n17771 104.41
R5244 vss.n18837 vss.n17780 104.41
R5245 vss.n18819 vss.n17799 104.41
R5246 vss.n18815 vss.n17803 104.41
R5247 vss.n18803 vss.n17807 104.41
R5248 vss.n18796 vss.n17818 104.41
R5249 vss.n18792 vss.n17822 104.41
R5250 vss.n18780 vss.n17826 104.41
R5251 vss.n18773 vss.n17837 104.41
R5252 vss.n18769 vss.n17841 104.41
R5253 vss.n17848 vss.n17841 104.41
R5254 vss.n18763 vss.n17847 104.41
R5255 vss.n18751 vss.n17852 104.41
R5256 vss.n18747 vss.n17861 104.41
R5257 vss.n18740 vss.n17868 104.41
R5258 vss.n18728 vss.n17871 104.41
R5259 vss.n18724 vss.n17880 104.41
R5260 vss.n18717 vss.n17887 104.41
R5261 vss.n18701 vss.n17903 104.41
R5262 vss.n18691 vss.n17909 104.41
R5263 vss.n18687 vss.n17916 104.41
R5264 vss.n18675 vss.n17920 104.41
R5265 vss.n18668 vss.n17931 104.41
R5266 vss.n18664 vss.n17935 104.41
R5267 vss.n18652 vss.n17939 104.41
R5268 vss.n18647 vss.n17949 104.41
R5269 vss.n18647 vss.n17950 104.41
R5270 vss.n17961 vss.n17953 104.41
R5271 vss.n18635 vss.n17959 104.41
R5272 vss.n18623 vss.n17965 104.41
R5273 vss.n18619 vss.n17974 104.41
R5274 vss.n18612 vss.n17981 104.41
R5275 vss.n18600 vss.n17984 104.41
R5276 vss.n18596 vss.n17993 104.41
R5277 vss.n18578 vss.n18012 104.41
R5278 vss.n18574 vss.n18016 104.41
R5279 vss.n18562 vss.n18020 104.41
R5280 vss.n18555 vss.n18031 104.41
R5281 vss.n18551 vss.n18035 104.41
R5282 vss.n18539 vss.n18039 104.41
R5283 vss.n18532 vss.n18050 104.41
R5284 vss.n18528 vss.n18054 104.41
R5285 vss.n18061 vss.n18054 104.41
R5286 vss.n18522 vss.n18060 104.41
R5287 vss.n18510 vss.n18065 104.41
R5288 vss.n18506 vss.n18074 104.41
R5289 vss.n18499 vss.n18081 104.41
R5290 vss.n18487 vss.n18084 104.41
R5291 vss.n18483 vss.n18093 104.41
R5292 vss.n18476 vss.n18100 104.41
R5293 vss.n18460 vss.n18116 104.41
R5294 vss.n18450 vss.n18122 104.41
R5295 vss.n18446 vss.n18129 104.41
R5296 vss.n18434 vss.n18133 104.41
R5297 vss.n18427 vss.n18144 104.41
R5298 vss.n18423 vss.n18148 104.41
R5299 vss.n18411 vss.n18152 104.41
R5300 vss.n18406 vss.n18162 104.41
R5301 vss.n18406 vss.n18163 104.41
R5302 vss.n18174 vss.n18166 104.41
R5303 vss.n18394 vss.n18172 104.41
R5304 vss.n18382 vss.n18178 104.41
R5305 vss.n18378 vss.n18187 104.41
R5306 vss.n18371 vss.n18194 104.41
R5307 vss.n18359 vss.n18197 104.41
R5308 vss.n18355 vss.n18206 104.41
R5309 vss.n18337 vss.n18225 104.41
R5310 vss.n18333 vss.n18229 104.41
R5311 vss.n18321 vss.n18233 104.41
R5312 vss.n18314 vss.n18244 104.41
R5313 vss.n18310 vss.n18248 104.41
R5314 vss.n18298 vss.n18252 104.41
R5315 vss.n18291 vss.n18263 104.41
R5316 vss.n18287 vss.n18267 104.41
R5317 vss.n18276 vss.n18267 104.41
R5318 vss.n18281 vss.n18275 104.41
R5319 vss.n20293 vss.n17620 104.41
R5320 vss.n20281 vss.n19035 104.41
R5321 vss.n20281 vss.n19037 104.41
R5322 vss.n20273 vss.n19039 104.41
R5323 vss.n20269 vss.n19049 104.41
R5324 vss.n20257 vss.n19051 104.41
R5325 vss.n20253 vss.n19061 104.41
R5326 vss.n20246 vss.n19068 104.41
R5327 vss.n20234 vss.n19071 104.41
R5328 vss.n20230 vss.n19080 104.41
R5329 vss.n20212 vss.n19099 104.41
R5330 vss.n20208 vss.n19103 104.41
R5331 vss.n20196 vss.n19107 104.41
R5332 vss.n20189 vss.n19118 104.41
R5333 vss.n20185 vss.n19122 104.41
R5334 vss.n20173 vss.n19126 104.41
R5335 vss.n20166 vss.n19137 104.41
R5336 vss.n20162 vss.n19141 104.41
R5337 vss.n20158 vss.n19141 104.41
R5338 vss.n20154 vss.n19146 104.41
R5339 vss.n20142 vss.n19150 104.41
R5340 vss.n20138 vss.n19159 104.41
R5341 vss.n20126 vss.n19161 104.41
R5342 vss.n20122 vss.n19171 104.41
R5343 vss.n20115 vss.n19178 104.41
R5344 vss.n20103 vss.n19181 104.41
R5345 vss.n20088 vss.n19197 104.41
R5346 vss.n20078 vss.n19203 104.41
R5347 vss.n20074 vss.n19210 104.41
R5348 vss.n20062 vss.n19214 104.41
R5349 vss.n20055 vss.n19225 104.41
R5350 vss.n20051 vss.n19229 104.41
R5351 vss.n20039 vss.n19233 104.41
R5352 vss.n20034 vss.n19243 104.41
R5353 vss.n20034 vss.n19244 104.41
R5354 vss.n19255 vss.n19247 104.41
R5355 vss.n20022 vss.n19253 104.41
R5356 vss.n20010 vss.n19259 104.41
R5357 vss.n20006 vss.n19268 104.41
R5358 vss.n19999 vss.n19275 104.41
R5359 vss.n19987 vss.n19278 104.41
R5360 vss.n19983 vss.n19287 104.41
R5361 vss.n19965 vss.n19306 104.41
R5362 vss.n19961 vss.n19310 104.41
R5363 vss.n19949 vss.n19314 104.41
R5364 vss.n19942 vss.n19325 104.41
R5365 vss.n19938 vss.n19329 104.41
R5366 vss.n19926 vss.n19333 104.41
R5367 vss.n19919 vss.n19344 104.41
R5368 vss.n19915 vss.n19348 104.41
R5369 vss.n19911 vss.n19348 104.41
R5370 vss.n19907 vss.n19353 104.41
R5371 vss.n19895 vss.n19357 104.41
R5372 vss.n19891 vss.n19366 104.41
R5373 vss.n19879 vss.n19368 104.41
R5374 vss.n19875 vss.n19378 104.41
R5375 vss.n19868 vss.n19385 104.41
R5376 vss.n19856 vss.n19388 104.41
R5377 vss.n19841 vss.n19404 104.41
R5378 vss.n19831 vss.n19410 104.41
R5379 vss.n19827 vss.n19417 104.41
R5380 vss.n19815 vss.n19421 104.41
R5381 vss.n19808 vss.n19432 104.41
R5382 vss.n19804 vss.n19436 104.41
R5383 vss.n19792 vss.n19440 104.41
R5384 vss.n19787 vss.n19450 104.41
R5385 vss.n19787 vss.n19451 104.41
R5386 vss.n19462 vss.n19454 104.41
R5387 vss.n19775 vss.n19460 104.41
R5388 vss.n19763 vss.n19466 104.41
R5389 vss.n19759 vss.n19475 104.41
R5390 vss.n19752 vss.n19482 104.41
R5391 vss.n19740 vss.n19485 104.41
R5392 vss.n19736 vss.n19494 104.41
R5393 vss.n19718 vss.n19513 104.41
R5394 vss.n19714 vss.n19517 104.41
R5395 vss.n19702 vss.n19521 104.41
R5396 vss.n19695 vss.n19532 104.41
R5397 vss.n19691 vss.n19536 104.41
R5398 vss.n19679 vss.n19540 104.41
R5399 vss.n19672 vss.n19551 104.41
R5400 vss.n19668 vss.n19555 104.41
R5401 vss.n19664 vss.n19555 104.41
R5402 vss.n19660 vss.n19560 104.41
R5403 vss.n19648 vss.n19564 104.41
R5404 vss.n19644 vss.n19573 104.41
R5405 vss.n19632 vss.n19575 104.41
R5406 vss.n19628 vss.n19585 104.41
R5407 vss.n19603 vss.n19602 104.41
R5408 vss.n19610 vss.n19595 104.41
R5409 vss.n20350 vss.n17596 104.41
R5410 vss.n20344 vss.n20343 104.41
R5411 vss.n20339 vss.n20337 104.41
R5412 vss.n20333 vss.n20332 104.41
R5413 vss.n20324 vss.n17605 104.41
R5414 vss.n20319 vss.n17607 104.41
R5415 vss.n20313 vss.n17612 104.41
R5416 vss.n20309 vss.n17612 104.41
R5417 vss.n20301 vss.n17616 104.41
R5418 vss.n5630 vss.n4238 104.41
R5419 vss.n5626 vss.n4245 104.41
R5420 vss.n5622 vss.n4245 104.41
R5421 vss.n5618 vss.n4249 104.41
R5422 vss.n5606 vss.n4253 104.41
R5423 vss.n5602 vss.n4262 104.41
R5424 vss.n5590 vss.n4264 104.41
R5425 vss.n5586 vss.n4274 104.41
R5426 vss.n5579 vss.n4281 104.41
R5427 vss.n5567 vss.n4284 104.41
R5428 vss.n5552 vss.n4300 104.41
R5429 vss.n5542 vss.n4306 104.41
R5430 vss.n5538 vss.n4313 104.41
R5431 vss.n5526 vss.n4317 104.41
R5432 vss.n5519 vss.n4328 104.41
R5433 vss.n5515 vss.n4332 104.41
R5434 vss.n5503 vss.n4336 104.41
R5435 vss.n5498 vss.n4346 104.41
R5436 vss.n5498 vss.n4347 104.41
R5437 vss.n4358 vss.n4350 104.41
R5438 vss.n5486 vss.n4356 104.41
R5439 vss.n5474 vss.n4362 104.41
R5440 vss.n5470 vss.n4371 104.41
R5441 vss.n5463 vss.n4378 104.41
R5442 vss.n5451 vss.n4381 104.41
R5443 vss.n5447 vss.n4390 104.41
R5444 vss.n5429 vss.n4409 104.41
R5445 vss.n5425 vss.n4413 104.41
R5446 vss.n5413 vss.n4417 104.41
R5447 vss.n5406 vss.n4428 104.41
R5448 vss.n5402 vss.n4432 104.41
R5449 vss.n5390 vss.n4436 104.41
R5450 vss.n5383 vss.n4447 104.41
R5451 vss.n5379 vss.n4451 104.41
R5452 vss.n4458 vss.n4451 104.41
R5453 vss.n5373 vss.n4457 104.41
R5454 vss.n5361 vss.n4462 104.41
R5455 vss.n5357 vss.n4471 104.41
R5456 vss.n5350 vss.n4478 104.41
R5457 vss.n5338 vss.n4481 104.41
R5458 vss.n5334 vss.n4490 104.41
R5459 vss.n5327 vss.n4497 104.41
R5460 vss.n5311 vss.n4513 104.41
R5461 vss.n5301 vss.n4519 104.41
R5462 vss.n5297 vss.n4526 104.41
R5463 vss.n5285 vss.n4530 104.41
R5464 vss.n5278 vss.n4541 104.41
R5465 vss.n5274 vss.n4545 104.41
R5466 vss.n5262 vss.n4549 104.41
R5467 vss.n5257 vss.n4559 104.41
R5468 vss.n5257 vss.n4560 104.41
R5469 vss.n4571 vss.n4563 104.41
R5470 vss.n5245 vss.n4569 104.41
R5471 vss.n5233 vss.n4575 104.41
R5472 vss.n5229 vss.n4584 104.41
R5473 vss.n5222 vss.n4591 104.41
R5474 vss.n5210 vss.n4594 104.41
R5475 vss.n5206 vss.n4603 104.41
R5476 vss.n5188 vss.n4622 104.41
R5477 vss.n5184 vss.n4626 104.41
R5478 vss.n5172 vss.n4630 104.41
R5479 vss.n5165 vss.n4641 104.41
R5480 vss.n5161 vss.n4645 104.41
R5481 vss.n5149 vss.n4649 104.41
R5482 vss.n5142 vss.n4660 104.41
R5483 vss.n5138 vss.n4664 104.41
R5484 vss.n4671 vss.n4664 104.41
R5485 vss.n5132 vss.n4670 104.41
R5486 vss.n5120 vss.n4675 104.41
R5487 vss.n5116 vss.n4684 104.41
R5488 vss.n5109 vss.n4691 104.41
R5489 vss.n5097 vss.n4694 104.41
R5490 vss.n5093 vss.n4703 104.41
R5491 vss.n5086 vss.n4710 104.41
R5492 vss.n5070 vss.n4726 104.41
R5493 vss.n5060 vss.n4732 104.41
R5494 vss.n5056 vss.n4739 104.41
R5495 vss.n5044 vss.n4743 104.41
R5496 vss.n5037 vss.n4754 104.41
R5497 vss.n5033 vss.n4758 104.41
R5498 vss.n5021 vss.n4762 104.41
R5499 vss.n5016 vss.n4772 104.41
R5500 vss.n5016 vss.n4773 104.41
R5501 vss.n4784 vss.n4776 104.41
R5502 vss.n5004 vss.n4782 104.41
R5503 vss.n4992 vss.n4788 104.41
R5504 vss.n4988 vss.n4797 104.41
R5505 vss.n4981 vss.n4804 104.41
R5506 vss.n4969 vss.n4807 104.41
R5507 vss.n4965 vss.n4816 104.41
R5508 vss.n4947 vss.n4835 104.41
R5509 vss.n4943 vss.n4839 104.41
R5510 vss.n4931 vss.n4843 104.41
R5511 vss.n4924 vss.n4854 104.41
R5512 vss.n4920 vss.n4858 104.41
R5513 vss.n4908 vss.n4862 104.41
R5514 vss.n4901 vss.n4873 104.41
R5515 vss.n4897 vss.n4877 104.41
R5516 vss.n4886 vss.n4877 104.41
R5517 vss.n4891 vss.n4885 104.41
R5518 vss.n6903 vss.n4230 104.41
R5519 vss.n6891 vss.n5645 104.41
R5520 vss.n6891 vss.n5647 104.41
R5521 vss.n6883 vss.n5649 104.41
R5522 vss.n6879 vss.n5659 104.41
R5523 vss.n6867 vss.n5661 104.41
R5524 vss.n6863 vss.n5671 104.41
R5525 vss.n6856 vss.n5678 104.41
R5526 vss.n6844 vss.n5681 104.41
R5527 vss.n6840 vss.n5690 104.41
R5528 vss.n6822 vss.n5709 104.41
R5529 vss.n6818 vss.n5713 104.41
R5530 vss.n6806 vss.n5717 104.41
R5531 vss.n6799 vss.n5728 104.41
R5532 vss.n6795 vss.n5732 104.41
R5533 vss.n6783 vss.n5736 104.41
R5534 vss.n6776 vss.n5747 104.41
R5535 vss.n6772 vss.n5751 104.41
R5536 vss.n6768 vss.n5751 104.41
R5537 vss.n6764 vss.n5756 104.41
R5538 vss.n6752 vss.n5760 104.41
R5539 vss.n6748 vss.n5769 104.41
R5540 vss.n6736 vss.n5771 104.41
R5541 vss.n6732 vss.n5781 104.41
R5542 vss.n6725 vss.n5788 104.41
R5543 vss.n6713 vss.n5791 104.41
R5544 vss.n6698 vss.n5807 104.41
R5545 vss.n6688 vss.n5813 104.41
R5546 vss.n6684 vss.n5820 104.41
R5547 vss.n6672 vss.n5824 104.41
R5548 vss.n6665 vss.n5835 104.41
R5549 vss.n6661 vss.n5839 104.41
R5550 vss.n6649 vss.n5843 104.41
R5551 vss.n6644 vss.n5853 104.41
R5552 vss.n6644 vss.n5854 104.41
R5553 vss.n5865 vss.n5857 104.41
R5554 vss.n6632 vss.n5863 104.41
R5555 vss.n6620 vss.n5869 104.41
R5556 vss.n6616 vss.n5878 104.41
R5557 vss.n6609 vss.n5885 104.41
R5558 vss.n6597 vss.n5888 104.41
R5559 vss.n6593 vss.n5897 104.41
R5560 vss.n6575 vss.n5916 104.41
R5561 vss.n6571 vss.n5920 104.41
R5562 vss.n6559 vss.n5924 104.41
R5563 vss.n6552 vss.n5935 104.41
R5564 vss.n6548 vss.n5939 104.41
R5565 vss.n6536 vss.n5943 104.41
R5566 vss.n6529 vss.n5954 104.41
R5567 vss.n6525 vss.n5958 104.41
R5568 vss.n6521 vss.n5958 104.41
R5569 vss.n6517 vss.n5963 104.41
R5570 vss.n6505 vss.n5967 104.41
R5571 vss.n6501 vss.n5976 104.41
R5572 vss.n6489 vss.n5978 104.41
R5573 vss.n6485 vss.n5988 104.41
R5574 vss.n6478 vss.n5995 104.41
R5575 vss.n6466 vss.n5998 104.41
R5576 vss.n6451 vss.n6014 104.41
R5577 vss.n6441 vss.n6020 104.41
R5578 vss.n6437 vss.n6027 104.41
R5579 vss.n6425 vss.n6031 104.41
R5580 vss.n6418 vss.n6042 104.41
R5581 vss.n6414 vss.n6046 104.41
R5582 vss.n6402 vss.n6050 104.41
R5583 vss.n6397 vss.n6060 104.41
R5584 vss.n6397 vss.n6061 104.41
R5585 vss.n6072 vss.n6064 104.41
R5586 vss.n6385 vss.n6070 104.41
R5587 vss.n6373 vss.n6076 104.41
R5588 vss.n6369 vss.n6085 104.41
R5589 vss.n6362 vss.n6092 104.41
R5590 vss.n6350 vss.n6095 104.41
R5591 vss.n6346 vss.n6104 104.41
R5592 vss.n6328 vss.n6123 104.41
R5593 vss.n6324 vss.n6127 104.41
R5594 vss.n6312 vss.n6131 104.41
R5595 vss.n6305 vss.n6142 104.41
R5596 vss.n6301 vss.n6146 104.41
R5597 vss.n6289 vss.n6150 104.41
R5598 vss.n6282 vss.n6161 104.41
R5599 vss.n6278 vss.n6165 104.41
R5600 vss.n6274 vss.n6165 104.41
R5601 vss.n6270 vss.n6170 104.41
R5602 vss.n6258 vss.n6174 104.41
R5603 vss.n6254 vss.n6183 104.41
R5604 vss.n6242 vss.n6185 104.41
R5605 vss.n6238 vss.n6195 104.41
R5606 vss.n6213 vss.n6212 104.41
R5607 vss.n6220 vss.n6205 104.41
R5608 vss.n6960 vss.n4206 104.41
R5609 vss.n6954 vss.n6953 104.41
R5610 vss.n6949 vss.n6947 104.41
R5611 vss.n6943 vss.n6942 104.41
R5612 vss.n6934 vss.n4215 104.41
R5613 vss.n6929 vss.n4217 104.41
R5614 vss.n6923 vss.n4222 104.41
R5615 vss.n6919 vss.n4222 104.41
R5616 vss.n6911 vss.n4226 104.41
R5617 vss.n21852 vss.n21851 104.172
R5618 vss.n21734 vss.n21733 104.172
R5619 vss.n21744 vss.n21743 104.172
R5620 vss.n3801 vss.n3800 104.172
R5621 vss.n3683 vss.n3682 104.172
R5622 vss.n3693 vss.n3692 104.172
R5623 vss.n20531 vss.n20529 104.1
R5624 vss.n20558 vss.n20557 104.1
R5625 vss.n20760 vss.n20758 104.1
R5626 vss.n20780 vss.n20779 104.1
R5627 vss.n7141 vss.n7139 104.1
R5628 vss.n7168 vss.n7167 104.1
R5629 vss.n7370 vss.n7368 104.1
R5630 vss.n7390 vss.n7389 104.1
R5631 vss.n1757 vss.n1755 104.1
R5632 vss.n1777 vss.n1776 104.1
R5633 vss.n1988 vss.n1986 104.1
R5634 vss.n1616 vss.t33 104.1
R5635 vss.n2261 vss.n2260 104.1
R5636 vss.n2477 vss.n2475 104.1
R5637 vss.n2505 vss.n2504 104.1
R5638 vss.n2722 vss.n2720 104.1
R5639 vss.n2750 vss.n2749 104.1
R5640 vss.n2960 vss.n2958 104.1
R5641 vss.n1496 vss.t15 104.1
R5642 vss.n3233 vss.n3232 104.1
R5643 vss.n15206 vss.n15204 104.1
R5644 vss.n15186 vss.n15185 104.1
R5645 vss.n218 vss.n216 104.1
R5646 vss.n238 vss.n237 104.1
R5647 vss.n449 vss.n447 104.1
R5648 vss.n77 vss.t237 104.1
R5649 vss.n722 vss.n721 104.1
R5650 vss.n938 vss.n936 104.1
R5651 vss.n966 vss.n965 104.1
R5652 vss.n1183 vss.n1181 104.1
R5653 vss.n1211 vss.n1210 104.1
R5654 vss.n23306 vss.n23304 104.1
R5655 vss.n1354 vss.t257 104.1
R5656 vss.n23033 vss.n23032 104.1
R5657 vss.n1399 vss.n1397 104.1
R5658 vss.n22820 vss.n22819 104.1
R5659 vss.n11550 vss.n11549 103.937
R5660 vss.n11519 vss.n11518 103.937
R5661 vss.n12989 vss.n12988 103.937
R5662 vss.n12979 vss.n12978 103.937
R5663 vss.n12948 vss.n12947 103.937
R5664 vss.n13159 vss.n13158 103.937
R5665 vss.n12389 vss.n12388 103.937
R5666 vss.n12362 vss.n12361 103.937
R5667 vss.n10693 vss.n10692 103.937
R5668 vss.n10703 vss.n10702 103.937
R5669 vss.n13416 vss.n13415 103.937
R5670 vss.n13495 vss.n13494 103.937
R5671 vss.n13075 vss.n13074 103.937
R5672 vss.n10628 vss.n10627 103.937
R5673 vss.n10788 vss.n10787 103.937
R5674 vss.n12296 vss.n12295 103.937
R5675 vss.n14160 vss.n14159 103.937
R5676 vss.n14117 vss.n14116 103.937
R5677 vss.n13736 vss.n13735 103.937
R5678 vss.n11433 vss.n11432 103.937
R5679 vss.n11873 vss.n11872 103.937
R5680 vss.n11909 vss.n11908 103.937
R5681 vss.n13783 vss.n13782 103.937
R5682 vss.n13794 vss.n13793 103.937
R5683 vss.n18953 vss.n17683 102.44
R5684 vss.n18946 vss.n17683 102.44
R5685 vss.n18830 vss.n17787 102.44
R5686 vss.n18826 vss.n17787 102.44
R5687 vss.n17899 vss.n17890 102.44
R5688 vss.n18705 vss.n17899 102.44
R5689 vss.n18589 vss.n18000 102.44
R5690 vss.n18585 vss.n18000 102.44
R5691 vss.n18112 vss.n18103 102.44
R5692 vss.n18464 vss.n18112 102.44
R5693 vss.n18348 vss.n18213 102.44
R5694 vss.n18344 vss.n18213 102.44
R5695 vss.n20223 vss.n19087 102.44
R5696 vss.n20219 vss.n19087 102.44
R5697 vss.n20099 vss.n19190 102.44
R5698 vss.n20092 vss.n19190 102.44
R5699 vss.n19976 vss.n19294 102.44
R5700 vss.n19972 vss.n19294 102.44
R5701 vss.n19852 vss.n19396 102.44
R5702 vss.n19845 vss.n19396 102.44
R5703 vss.n19729 vss.n19501 102.44
R5704 vss.n19725 vss.n19501 102.44
R5705 vss.n20357 vss.n17593 102.44
R5706 vss.n20353 vss.n17593 102.44
R5707 vss.n5563 vss.n4293 102.44
R5708 vss.n5556 vss.n4293 102.44
R5709 vss.n5440 vss.n4397 102.44
R5710 vss.n5436 vss.n4397 102.44
R5711 vss.n4509 vss.n4500 102.44
R5712 vss.n5315 vss.n4509 102.44
R5713 vss.n5199 vss.n4610 102.44
R5714 vss.n5195 vss.n4610 102.44
R5715 vss.n4722 vss.n4713 102.44
R5716 vss.n5074 vss.n4722 102.44
R5717 vss.n4958 vss.n4823 102.44
R5718 vss.n4954 vss.n4823 102.44
R5719 vss.n6833 vss.n5697 102.44
R5720 vss.n6829 vss.n5697 102.44
R5721 vss.n6709 vss.n5800 102.44
R5722 vss.n6702 vss.n5800 102.44
R5723 vss.n6586 vss.n5904 102.44
R5724 vss.n6582 vss.n5904 102.44
R5725 vss.n6462 vss.n6006 102.44
R5726 vss.n6455 vss.n6006 102.44
R5727 vss.n6339 vss.n6111 102.44
R5728 vss.n6335 vss.n6111 102.44
R5729 vss.n6967 vss.n4203 102.44
R5730 vss.n6963 vss.n4203 102.44
R5731 vss.n16794 vss.n16788 102.44
R5732 vss.n17025 vss.n17019 102.44
R5733 vss.n17263 vss.n17257 102.44
R5734 vss.n16071 vss.n16065 102.44
R5735 vss.n15237 vss.n15233 102.44
R5736 vss.n15545 vss.n15539 102.44
R5737 vss.n15779 vss.n15773 102.44
R5738 vss.n16492 vss.n16486 102.44
R5739 vss.n22706 vss.n22704 102.362
R5740 vss.n22687 vss.n22681 102.362
R5741 vss.n22498 vss.n22496 102.362
R5742 vss.n22479 vss.n22473 102.362
R5743 vss.n22290 vss.n22288 102.362
R5744 vss.n22271 vss.n22265 102.362
R5745 vss.n22080 vss.n22078 102.362
R5746 vss.n21601 vss.n21595 102.362
R5747 vss.n21426 vss.n21424 102.362
R5748 vss.n21407 vss.n21401 102.362
R5749 vss.n21218 vss.n21216 102.362
R5750 vss.n21199 vss.n21193 102.362
R5751 vss.n21010 vss.n21008 102.362
R5752 vss.n20991 vss.n20985 102.362
R5753 vss.n8869 vss.n8867 102.362
R5754 vss.n8850 vss.n8844 102.362
R5755 vss.n8661 vss.n8659 102.362
R5756 vss.n8642 vss.n8636 102.362
R5757 vss.n8453 vss.n8451 102.362
R5758 vss.n8434 vss.n8428 102.362
R5759 vss.n8240 vss.n8238 102.362
R5760 vss.n8227 vss.n8221 102.362
R5761 vss.n8037 vss.n8035 102.362
R5762 vss.n8018 vss.n8012 102.362
R5763 vss.n7828 vss.n7826 102.362
R5764 vss.n7809 vss.n7803 102.362
R5765 vss.n7620 vss.n7618 102.362
R5766 vss.n7601 vss.n7595 102.362
R5767 vss.n20647 vss.n20645 97.16
R5768 vss.n20665 vss.n20663 97.16
R5769 vss.n7257 vss.n7255 97.16
R5770 vss.n7275 vss.n7273 97.16
R5771 vss.n1868 vss.n1866 97.16
R5772 vss.n1887 vss.n1884 97.16
R5773 vss.n1904 vss.t53 97.16
R5774 vss.n2113 vss.n2110 97.16
R5775 vss.n2131 vss.n2128 97.16
R5776 vss.n2357 vss.n2354 97.16
R5777 vss.n2375 vss.n2372 97.16
R5778 vss.n2601 vss.n2598 97.16
R5779 vss.n2620 vss.n2617 97.16
R5780 vss.n2839 vss.n2837 97.16
R5781 vss.n2858 vss.n2855 97.16
R5782 vss.n3084 vss.n3081 97.16
R5783 vss.n3102 vss.n3099 97.16
R5784 vss.n3313 vss.t49 97.16
R5785 vss.n3328 vss.n3325 97.16
R5786 vss.n3346 vss.n3344 97.16
R5787 vss.n329 vss.n327 97.16
R5788 vss.n348 vss.n345 97.16
R5789 vss.n365 vss.t263 97.16
R5790 vss.n574 vss.n571 97.16
R5791 vss.n592 vss.n589 97.16
R5792 vss.n818 vss.n815 97.16
R5793 vss.n836 vss.n833 97.16
R5794 vss.n1062 vss.n1059 97.16
R5795 vss.n1081 vss.n1078 97.16
R5796 vss.n1307 vss.n1304 97.16
R5797 vss.n23401 vss.n23398 97.16
R5798 vss.n23176 vss.n23173 97.16
R5799 vss.n23158 vss.n23155 97.16
R5800 vss.n22949 vss.t269 97.16
R5801 vss.n22932 vss.n22929 97.16
R5802 vss.n22913 vss.n22911 97.16
R5803 vss.n12051 vss.n12050 92.705
R5804 vss.n12041 vss.n12040 92.705
R5805 vss.n10970 vss.n10969 92.705
R5806 vss.n10980 vss.n10979 92.705
R5807 vss.n13833 vss.n13832 92.705
R5808 vss.n13823 vss.n13822 92.705
R5809 vss.n11125 vss.n11124 92.705
R5810 vss.n11115 vss.n11114 92.705
R5811 vss.n13364 vss.n13363 92.705
R5812 vss.n13384 vss.n13383 92.705
R5813 vss.n14196 vss.n14195 92.705
R5814 vss.n14206 vss.n14205 92.705
R5815 vss.n12889 vss.n12888 92.705
R5816 vss.n12886 vss.n12884 92.705
R5817 vss.n12480 vss.n12479 92.705
R5818 vss.n12477 vss.n12475 92.705
R5819 vss.n20513 vss.n20512 90.22
R5820 vss.n20573 vss.n20572 90.22
R5821 vss.n20741 vss.n20740 90.22
R5822 vss.n20795 vss.n20794 90.22
R5823 vss.n7123 vss.n7122 90.22
R5824 vss.n7183 vss.n7182 90.22
R5825 vss.n7351 vss.n7350 90.22
R5826 vss.n7405 vss.n7404 90.22
R5827 vss.n1735 vss.n1734 90.22
R5828 vss.n1794 vss.n1793 90.22
R5829 vss.n2033 vss.n2032 90.22
R5830 vss.n2213 vss.n2212 90.22
R5831 vss.n2457 vss.n2456 90.22
R5832 vss.n2522 vss.n2521 90.22
R5833 vss.n2701 vss.n2700 90.22
R5834 vss.n2766 vss.n2765 90.22
R5835 vss.n3004 vss.n3003 90.22
R5836 vss.n3184 vss.n3183 90.22
R5837 vss.n3422 vss.n3421 90.22
R5838 vss.n3463 vss.n3462 90.22
R5839 vss.n196 vss.n195 90.22
R5840 vss.n255 vss.n254 90.22
R5841 vss.n494 vss.n493 90.22
R5842 vss.n674 vss.n673 90.22
R5843 vss.n918 vss.n917 90.22
R5844 vss.n983 vss.n982 90.22
R5845 vss.n1162 vss.n1161 90.22
R5846 vss.n1227 vss.n1226 90.22
R5847 vss.n23258 vss.n23257 90.22
R5848 vss.n23078 vss.n23077 90.22
R5849 vss.n22837 vss.n22836 90.22
R5850 vss.n1438 vss.n1437 90.22
R5851 vss.n17604 vss.n17602 87.419
R5852 vss.n4214 vss.n4212 87.419
R5853 vss.n12120 vss.n12118 86.911
R5854 vss.n12130 vss.n12128 86.911
R5855 vss.n10880 vss.n10878 86.911
R5856 vss.n11948 vss.n11946 86.911
R5857 vss.n14419 vss.n14417 86.911
R5858 vss.n14373 vss.n14371 86.911
R5859 vss.n11637 vss.n11635 86.911
R5860 vss.n11664 vss.n11662 86.911
R5861 vss.n13274 vss.n13272 86.911
R5862 vss.n13258 vss.n13256 86.911
R5863 vss.n13543 vss.n13541 86.911
R5864 vss.n14595 vss.n14593 86.911
R5865 vss.n14835 vss.n14833 86.911
R5866 vss.n14863 vss.n14861 86.911
R5867 vss.n10488 vss.n10486 86.911
R5868 vss.n10518 vss.n10516 86.911
R5869 vss.n20233 vss.n20232 86.842
R5870 vss.n20210 vss.n20209 86.842
R5871 vss.n20113 vss.n20112 86.842
R5872 vss.n19208 vss.n19207 86.842
R5873 vss.n19986 vss.n19985 86.842
R5874 vss.n19963 vss.n19962 86.842
R5875 vss.n19866 vss.n19865 86.842
R5876 vss.n19853 ldomc_0.otaldom_0.nmoslm_0.vss 86.842
R5877 vss.n19415 vss.n19414 86.842
R5878 vss.n19739 vss.n19738 86.842
R5879 vss.n19716 vss.n19715 86.842
R5880 vss.n19607 vss.n19596 86.842
R5881 vss.n20347 vss.n17597 86.842
R5882 vss.n18967 vss.n18966 86.842
R5883 vss.n17701 vss.n17700 86.842
R5884 vss.n18840 vss.n18839 86.842
R5885 vss.n18817 vss.n18816 86.842
R5886 vss.n17888 vss.n17879 86.842
R5887 vss.n17914 vss.n17913 86.842
R5888 vss.n18599 vss.n18598 86.842
R5889 vss.n18576 vss.n18575 86.842
R5890 vss.n18101 vss.n18092 86.842
R5891 vss.n18127 vss.n18126 86.842
R5892 vss.n18358 vss.n18357 86.842
R5893 vss.n18335 vss.n18334 86.842
R5894 vss.n6843 vss.n6842 86.842
R5895 vss.n6820 vss.n6819 86.842
R5896 vss.n6723 vss.n6722 86.842
R5897 vss.n5818 vss.n5817 86.842
R5898 vss.n6596 vss.n6595 86.842
R5899 vss.n6573 vss.n6572 86.842
R5900 vss.n6476 vss.n6475 86.842
R5901 vss.n6463 bandgapmd_0.otam_1.nmoslm_0.vss 86.842
R5902 vss.n6025 vss.n6024 86.842
R5903 vss.n6349 vss.n6348 86.842
R5904 vss.n6326 vss.n6325 86.842
R5905 vss.n6217 vss.n6206 86.842
R5906 vss.n6957 vss.n4207 86.842
R5907 vss.n5577 vss.n5576 86.842
R5908 vss.n4311 vss.n4310 86.842
R5909 vss.n5450 vss.n5449 86.842
R5910 vss.n5427 vss.n5426 86.842
R5911 vss.n4498 vss.n4489 86.842
R5912 vss.n4524 vss.n4523 86.842
R5913 vss.n5209 vss.n5208 86.842
R5914 vss.n5186 vss.n5185 86.842
R5915 vss.n4711 vss.n4702 86.842
R5916 vss.n4737 vss.n4736 86.842
R5917 vss.n4968 vss.n4967 86.842
R5918 vss.n4945 vss.n4944 86.842
R5919 vss.n16762 vss.n16761 86.842
R5920 vss.n16803 vss.n16802 86.842
R5921 vss.n16992 vss.n16991 86.842
R5922 vss.n17037 vss.n17036 86.842
R5923 vss.n17228 vss.n17227 86.842
R5924 vss.n17292 vss.n17291 86.842
R5925 vss.n16038 vss.n16037 86.842
R5926 vss.n16082 vss.n16081 86.842
R5927 vss.n15245 vss.n15244 86.842
R5928 vss.n15223 vss.n15222 86.842
R5929 vss.n15512 vss.n15511 86.842
R5930 vss.n15559 vss.n15558 86.842
R5931 vss.n15748 vss.n15747 86.842
R5932 vss.n15789 vss.n15788 86.842
R5933 vss.n16459 vss.n16458 86.842
R5934 vss.n16506 vss.n16505 86.842
R5935 vss.n1670 vss.n1668 86.211
R5936 vss.n15142 vss.n15139 86.211
R5937 vss.n131 vss.n129 86.211
R5938 vss.n22776 vss.n22773 86.211
R5939 vss.n22600 vss.n22599 85.714
R5940 vss.n22581 vss.n22580 85.714
R5941 vss.n22392 vss.n22391 85.714
R5942 vss.n22373 vss.n22372 85.714
R5943 vss.n22184 vss.n22183 85.714
R5944 vss.n22165 vss.n22164 85.714
R5945 vss.n21528 vss.n21527 85.714
R5946 vss.n21509 vss.n21508 85.714
R5947 vss.n21320 vss.n21319 85.714
R5948 vss.n21301 vss.n21300 85.714
R5949 vss.n21112 vss.n21111 85.714
R5950 vss.n21093 vss.n21092 85.714
R5951 vss.n20904 vss.n20903 85.714
R5952 vss.n8763 vss.n8762 85.714
R5953 vss.n8744 vss.n8743 85.714
R5954 vss.n8555 vss.n8554 85.714
R5955 vss.n8536 vss.n8535 85.714
R5956 vss.n8347 vss.n8346 85.714
R5957 vss.n8328 vss.n8327 85.714
R5958 vss.n8139 vss.n8138 85.714
R5959 vss.n8120 vss.n8119 85.714
R5960 vss.n7931 vss.n7930 85.714
R5961 vss.n7912 vss.n7911 85.714
R5962 vss.n7722 vss.n7721 85.714
R5963 vss.n7703 vss.n7702 85.714
R5964 vss.n7514 vss.n7513 85.714
R5965 vss.n20450 vss.n20448 83.28
R5966 vss.n20632 vss.n20630 83.28
R5967 vss.n20680 vss.n20678 83.28
R5968 vss.n20856 vss.n20854 83.28
R5969 vss.n7060 vss.n7058 83.28
R5970 vss.n7242 vss.n7240 83.28
R5971 vss.n7290 vss.n7288 83.28
R5972 vss.n7466 vss.n7464 83.28
R5973 vss.n1824 vss.t61 83.28
R5974 vss.n1853 vss.n1851 83.28
R5975 vss.n1903 vss.n1900 83.28
R5976 vss.n2096 vss.n2093 83.28
R5977 vss.n2147 vss.n2144 83.28
R5978 vss.n2233 vss.t13 83.28
R5979 vss.n2341 vss.n2338 83.28
R5980 vss.n2391 vss.n2388 83.28
R5981 vss.n2585 vss.n2582 83.28
R5982 vss.n2636 vss.n2633 83.28
R5983 vss.n2827 vss.n2825 83.28
R5984 vss.n2874 vss.n2871 83.28
R5985 vss.n2988 vss.t79 83.28
R5986 vss.n3068 vss.n3065 83.28
R5987 vss.n3119 vss.n3116 83.28
R5988 vss.n3312 vss.n3309 83.28
R5989 vss.n3361 vss.n3359 83.28
R5990 vss.n3392 vss.t77 83.28
R5991 vss.n285 vss.t243 83.28
R5992 vss.n314 vss.n312 83.28
R5993 vss.n364 vss.n361 83.28
R5994 vss.n557 vss.n554 83.28
R5995 vss.n608 vss.n605 83.28
R5996 vss.n694 vss.t303 83.28
R5997 vss.n802 vss.n799 83.28
R5998 vss.n852 vss.n849 83.28
R5999 vss.n1046 vss.n1043 83.28
R6000 vss.n1097 vss.n1094 83.28
R6001 vss.n1291 vss.n1288 83.28
R6002 vss.n23385 vss.n23382 83.28
R6003 vss.n23278 vss.t285 83.28
R6004 vss.n23192 vss.n23189 83.28
R6005 vss.n23141 vss.n23138 83.28
R6006 vss.n22948 vss.n22945 83.28
R6007 vss.n22898 vss.n22896 83.28
R6008 vss.n22869 vss.t287 83.28
R6009 vss.n20430 vss.n20428 83.199
R6010 vss.n20879 vss.n20876 83.199
R6011 vss.n7040 vss.n7038 83.199
R6012 vss.n7489 vss.n7486 83.199
R6013 vss.n12068 vss.n12067 81.117
R6014 vss.n10797 vss.n10796 81.117
R6015 vss.n10960 vss.n10959 81.117
R6016 vss.n11000 vss.n10999 81.117
R6017 vss.n13850 vss.n13849 81.117
R6018 vss.n14071 vss.n14070 81.117
R6019 vss.n11717 vss.n11716 81.117
R6020 vss.n11061 vss.n11060 81.117
R6021 vss.n13348 vss.n13347 81.117
R6022 vss.n14693 vss.n14692 81.117
R6023 vss.n14186 vss.n14185 81.117
R6024 vss.n14228 vss.n14227 81.117
R6025 vss.n12868 vss.n12867 81.117
R6026 vss.n12911 vss.n12910 81.117
R6027 vss.n12463 vss.n12462 81.117
R6028 vss.n12498 vss.n12497 81.117
R6029 vss.n20889 vss.n20888 80.971
R6030 vss.n20438 vss.n20437 80.971
R6031 vss.n20432 vss.n20431 80.971
R6032 vss.n7499 vss.n7498 80.971
R6033 vss.n7048 vss.n7047 80.971
R6034 vss.n7042 vss.n7041 80.971
R6035 vss.n15152 vss.n15151 80.971
R6036 vss.n1678 vss.n1677 80.971
R6037 vss.n1672 vss.n1671 80.971
R6038 vss.n22786 vss.n22785 80.971
R6039 vss.n139 vss.n138 80.971
R6040 vss.n133 vss.n132 80.971
R6041 vss.n9185 vss.t314 78.222
R6042 vss.n20497 vss.n20496 76.34
R6043 vss.n20588 vss.n20587 76.34
R6044 vss.n20726 vss.n20725 76.34
R6045 vss.n20811 vss.n20810 76.34
R6046 vss.n7107 vss.n7106 76.34
R6047 vss.n7198 vss.n7197 76.34
R6048 vss.n7336 vss.n7335 76.34
R6049 vss.n7421 vss.n7420 76.34
R6050 vss.n1809 vss.n1808 76.34
R6051 vss.n1952 vss.n1951 76.34
R6052 vss.n2049 vss.n2048 76.34
R6053 vss.n2197 vss.n2196 76.34
R6054 vss.t65 vss.n2276 76.34
R6055 vss.n2293 vss.n2292 76.34
R6056 vss.n2441 vss.n2440 76.34
R6057 vss.n2538 vss.n2537 76.34
R6058 vss.n2685 vss.n2684 76.34
R6059 vss.n2782 vss.n2781 76.34
R6060 vss.n2924 vss.n2923 76.34
R6061 vss.t31 vss.n2939 76.34
R6062 vss.n3021 vss.n3020 76.34
R6063 vss.n3168 vss.n3167 76.34
R6064 vss.n3265 vss.n3264 76.34
R6065 vss.n3407 vss.n3406 76.34
R6066 vss.n270 vss.n269 76.34
R6067 vss.n413 vss.n412 76.34
R6068 vss.n510 vss.n509 76.34
R6069 vss.n658 vss.n657 76.34
R6070 vss.t255 vss.n737 76.34
R6071 vss.n754 vss.n753 76.34
R6072 vss.n902 vss.n901 76.34
R6073 vss.n999 vss.n998 76.34
R6074 vss.n1146 vss.n1145 76.34
R6075 vss.n1243 vss.n1242 76.34
R6076 vss.n23338 vss.n23337 76.34
R6077 vss.t267 vss.n23321 76.34
R6078 vss.n23241 vss.n23240 76.34
R6079 vss.n23094 vss.n23093 76.34
R6080 vss.n22997 vss.n22996 76.34
R6081 vss.n22854 vss.n22853 76.34
R6082 vss.n12144 vss.n12142 75.323
R6083 vss.n11976 vss.n11974 75.323
R6084 vss.n11922 vss.n11920 75.323
R6085 vss.n14338 vss.n14336 75.323
R6086 vss.n11626 vss.n11624 75.323
R6087 vss.n11675 vss.n11673 75.323
R6088 vss.n14816 vss.n14814 75.323
R6089 vss.n14615 vss.n14613 75.323
R6090 vss.n14555 vss.n14553 75.323
R6091 vss.n14906 vss.n14904 75.323
R6092 vss.n15050 vss.n15048 75.323
R6093 vss.n10548 vss.n10546 75.323
R6094 vss.n9188 vss.n9185 73.333
R6095 vss.n12224 vss.n12223 69.529
R6096 vss.n12018 vss.n12017 69.529
R6097 vss.n11254 vss.n11253 69.529
R6098 vss.n11194 vss.n11193 69.529
R6099 vss.n13911 vss.n13910 69.529
R6100 vss.n14049 vss.n14048 69.529
R6101 vss.n11744 vss.n11743 69.529
R6102 vss.n11071 vss.n11070 69.529
R6103 vss.n14738 vss.n14737 69.529
R6104 vss.n14679 vss.n14678 69.529
R6105 vss.n14466 vss.n14465 69.529
R6106 vss.n14248 vss.n14247 69.529
R6107 vss.n12853 vss.n12852 69.529
R6108 vss.n12917 vss.n12915 69.529
R6109 vss.n12653 vss.n12652 69.529
R6110 vss.n12504 vss.n12502 69.529
R6111 vss.n20466 vss.n20464 69.4
R6112 vss.n20617 vss.n20615 69.4
R6113 vss.n20695 vss.n20693 69.4
R6114 vss.n20840 vss.n20838 69.4
R6115 vss.n7076 vss.n7074 69.4
R6116 vss.n7227 vss.n7225 69.4
R6117 vss.n7305 vss.n7303 69.4
R6118 vss.n7450 vss.n7448 69.4
R6119 vss.n1689 vss.n1687 69.4
R6120 vss.n1838 vss.n1836 69.4
R6121 vss.n1919 vss.n1916 69.4
R6122 vss.n2080 vss.n2077 69.4
R6123 vss.n2163 vss.n2160 69.4
R6124 vss.n2164 vss.t17 69.4
R6125 vss.n2325 vss.n2322 69.4
R6126 vss.n2408 vss.n2405 69.4
R6127 vss.n2569 vss.n2566 69.4
R6128 vss.n2652 vss.n2649 69.4
R6129 vss.n2812 vss.n2810 69.4
R6130 vss.n2890 vss.n2887 69.4
R6131 vss.n3053 vss.t83 69.4
R6132 vss.n3052 vss.n3049 69.4
R6133 vss.n3135 vss.n3132 69.4
R6134 vss.n3296 vss.n3293 69.4
R6135 vss.n3376 vss.n3374 69.4
R6136 vss.n3485 vss.n3483 69.4
R6137 vss.n150 vss.n148 69.4
R6138 vss.n299 vss.n297 69.4
R6139 vss.n380 vss.n377 69.4
R6140 vss.n541 vss.n538 69.4
R6141 vss.n624 vss.n621 69.4
R6142 vss.n625 vss.t281 69.4
R6143 vss.n786 vss.n783 69.4
R6144 vss.n869 vss.n866 69.4
R6145 vss.n1030 vss.n1027 69.4
R6146 vss.n1113 vss.n1110 69.4
R6147 vss.n1274 vss.n1271 69.4
R6148 vss.n23369 vss.n23366 69.4
R6149 vss.n23209 vss.t241 69.4
R6150 vss.n23208 vss.n23205 69.4
R6151 vss.n23125 vss.n23122 69.4
R6152 vss.n22964 vss.n22961 69.4
R6153 vss.n22883 vss.n22881 69.4
R6154 vss.n1460 vss.n1458 69.4
R6155 vss.n11478 vss.n11477 69.291
R6156 vss.n11696 vss.n11695 69.291
R6157 vss.n13118 vss.n13117 69.291
R6158 vss.n13667 vss.n13666 69.291
R6159 vss.n14983 vss.n14982 69.291
R6160 vss.n13145 vss.n13144 69.291
R6161 vss.n12410 vss.n12409 69.291
R6162 vss.n10673 vss.n10672 69.291
R6163 vss.n12327 vss.n12326 69.291
R6164 vss.n11488 vss.n11487 69.291
R6165 vss.n13376 vss.n13375 69.291
R6166 vss.n13459 vss.n13458 69.291
R6167 vss.n13090 vss.n13089 69.291
R6168 vss.n10643 vss.n10642 69.291
R6169 vss.n12312 vss.n12311 69.291
R6170 vss.n10809 vss.n10808 69.291
R6171 vss.n14564 vss.n14563 69.291
R6172 vss.n14101 vss.n14100 69.291
R6173 vss.n13751 vss.n13750 69.291
R6174 vss.n11448 vss.n11447 69.291
R6175 vss.n11857 vss.n11856 69.291
R6176 vss.n10934 vss.n10933 69.291
R6177 vss.n13654 vss.n13653 69.291
R6178 vss.n14063 vss.n14062 69.291
R6179 vss.n9636 vss.n9635 68.223
R6180 vss.n1682 vss.n1681 64.376
R6181 vss.n15154 vss.n15153 64.376
R6182 vss.n143 vss.n142 64.376
R6183 vss.n22788 vss.n22787 64.376
R6184 vss.n12172 vss.n12169 63.735
R6185 vss.n11990 vss.n11987 63.735
R6186 vss.n11324 vss.n11321 63.735
R6187 vss.n14312 vss.n14309 63.735
R6188 vss.n11612 vss.n11609 63.735
R6189 vss.n11825 vss.n11822 63.735
R6190 vss.n14802 vss.n14799 63.735
R6191 vss.n14629 vss.n14626 63.735
R6192 vss.n14540 vss.n14537 63.735
R6193 vss.n14261 vss.n14258 63.735
R6194 vss.n14893 vss.n14890 63.735
R6195 vss.n15055 vss.n15046 63.735
R6196 vss.n12705 vss.n12702 63.735
R6197 vss.n10179 vss.n10178 62.851
R6198 vss.n20482 vss.n20481 62.46
R6199 vss.n20603 vss.n20602 62.46
R6200 vss.n20711 vss.n20710 62.46
R6201 vss.n20826 vss.n20825 62.46
R6202 vss.n7092 vss.n7091 62.46
R6203 vss.n7213 vss.n7212 62.46
R6204 vss.n7321 vss.n7320 62.46
R6205 vss.n7436 vss.n7435 62.46
R6206 vss.n1705 vss.n1704 62.46
R6207 vss.n1824 vss.n1823 62.46
R6208 vss.n1936 vss.n1935 62.46
R6209 vss.t21 vss.n2016 62.46
R6210 vss.n2065 vss.n2064 62.46
R6211 vss.n2180 vss.n2179 62.46
R6212 vss.n2310 vss.n2309 62.46
R6213 vss.n2425 vss.n2424 62.46
R6214 vss.n2554 vss.n2553 62.46
R6215 vss.n2669 vss.n2668 62.46
R6216 vss.n2798 vss.n2797 62.46
R6217 vss.n2907 vss.n2906 62.46
R6218 vss.n3037 vss.n3036 62.46
R6219 vss.n3152 vss.n3151 62.46
R6220 vss.t37 vss.n3202 62.46
R6221 vss.n3281 vss.n3280 62.46
R6222 vss.n3392 vss.n3391 62.46
R6223 vss.n15165 vss.n15164 62.46
R6224 vss.n166 vss.n165 62.46
R6225 vss.n285 vss.n284 62.46
R6226 vss.n397 vss.n396 62.46
R6227 vss.t275 vss.n477 62.46
R6228 vss.n526 vss.n525 62.46
R6229 vss.n641 vss.n640 62.46
R6230 vss.n771 vss.n770 62.46
R6231 vss.n886 vss.n885 62.46
R6232 vss.n1015 vss.n1014 62.46
R6233 vss.n1130 vss.n1129 62.46
R6234 vss.n1259 vss.n1258 62.46
R6235 vss.n23354 vss.n23353 62.46
R6236 vss.n23225 vss.n23224 62.46
R6237 vss.n23110 vss.n23109 62.46
R6238 vss.t245 vss.n23060 62.46
R6239 vss.n22981 vss.n22980 62.46
R6240 vss.n22869 vss.n22868 62.46
R6241 vss.n22799 vss.n22798 62.46
R6242 vss.n20442 vss.n20441 59.858
R6243 vss.n20891 vss.n20890 59.858
R6244 vss.n7052 vss.n7051 59.858
R6245 vss.n7501 vss.n7500 59.858
R6246 vss.n20878 vss.n20877 59.468
R6247 vss.n20883 vss.n20882 59.468
R6248 vss.n7488 vss.n7487 59.468
R6249 vss.n7493 vss.n7492 59.468
R6250 vss.n15141 vss.n15140 59.468
R6251 vss.n15146 vss.n15145 59.468
R6252 vss.n22775 vss.n22774 59.468
R6253 vss.n22780 vss.n22779 59.468
R6254 vss.n12197 vss.n12196 57.941
R6255 vss.n12001 vss.n12000 57.941
R6256 vss.n11280 vss.n11279 57.941
R6257 vss.n11178 vss.n11177 57.941
R6258 vss.n13877 vss.n13876 57.941
R6259 vss.n13987 vss.n13986 57.941
R6260 vss.n11781 vss.n11780 57.941
R6261 vss.n11091 vss.n11090 57.941
R6262 vss.n14771 vss.n14770 57.941
R6263 vss.n13512 vss.n13511 57.941
R6264 vss.n14504 vss.n14503 57.941
R6265 vss.n14218 vss.n14217 57.941
R6266 vss.n12838 vss.n12837 57.941
R6267 vss.n12805 vss.n12804 57.941
R6268 vss.n12669 vss.n12668 57.941
R6269 vss.n12549 vss.n12548 57.941
R6270 vss.n20284 vss.n17619 57.894
R6271 vss.n20276 vss.n20275 57.894
R6272 vss.n20165 vss.n20164 57.894
R6273 vss.n20156 vss.n20155 57.894
R6274 vss.n20040 vss.n19234 57.894
R6275 vss.n20031 vss.n19246 57.894
R6276 vss.n19918 vss.n19917 57.894
R6277 vss.n19909 vss.n19908 57.894
R6278 vss.n19793 vss.n19441 57.894
R6279 vss.n19784 vss.n19453 57.894
R6280 vss.n19671 vss.n19670 57.894
R6281 vss.n19662 vss.n19661 57.894
R6282 vss.n17614 vss.n17613 57.894
R6283 vss.n20300 vss.n17615 57.894
R6284 vss.n19019 vss.n19018 57.894
R6285 vss.n19010 vss.n19009 57.894
R6286 vss.n18894 vss.n17727 57.894
R6287 vss.n18885 vss.n17739 57.894
R6288 vss.n18772 vss.n18771 57.894
R6289 vss.n18762 vss.n17850 57.894
R6290 vss.n18653 vss.n17940 57.894
R6291 vss.n18644 vss.n17952 57.894
R6292 vss.n18531 vss.n18530 57.894
R6293 vss.n18521 vss.n18063 57.894
R6294 vss.n18412 vss.n18153 57.894
R6295 vss.n18403 vss.n18165 57.894
R6296 vss.n18290 vss.n18289 57.894
R6297 vss.n18280 vss.n18278 57.894
R6298 vss.n6894 vss.n4229 57.894
R6299 vss.n6886 vss.n6885 57.894
R6300 vss.n6775 vss.n6774 57.894
R6301 vss.n6766 vss.n6765 57.894
R6302 vss.n6650 vss.n5844 57.894
R6303 vss.n6641 vss.n5856 57.894
R6304 vss.n6528 vss.n6527 57.894
R6305 vss.n6519 vss.n6518 57.894
R6306 vss.n6403 vss.n6051 57.894
R6307 vss.n6394 vss.n6063 57.894
R6308 vss.n6281 vss.n6280 57.894
R6309 vss.n6272 vss.n6271 57.894
R6310 vss.n4224 vss.n4223 57.894
R6311 vss.n6910 vss.n4225 57.894
R6312 vss.n5629 vss.n5628 57.894
R6313 vss.n5620 vss.n5619 57.894
R6314 vss.n5504 vss.n4337 57.894
R6315 vss.n5495 vss.n4349 57.894
R6316 vss.n5382 vss.n5381 57.894
R6317 vss.n5372 vss.n4460 57.894
R6318 vss.n5263 vss.n4550 57.894
R6319 vss.n5254 vss.n4562 57.894
R6320 vss.n5141 vss.n5140 57.894
R6321 vss.n5131 vss.n4673 57.894
R6322 vss.n5022 vss.n4763 57.894
R6323 vss.n5013 vss.n4775 57.894
R6324 vss.n4900 vss.n4899 57.894
R6325 vss.n4890 vss.n4888 57.894
R6326 vss.n16681 vss.n16680 57.894
R6327 vss.n16886 vss.n16885 57.894
R6328 vss.n16909 vss.n16908 57.894
R6329 vss.n17122 vss.n17121 57.894
R6330 vss.n17145 vss.n17144 57.894
R6331 vss.n16262 vss.n16261 57.894
R6332 vss.n15932 vss.n15931 57.894
R6333 vss.n15956 vss.n15955 57.894
R6334 vss.n16168 vss.n16167 57.894
R6335 vss.n16192 vss.n16191 57.894
R6336 vss.n16290 vss.n16289 57.894
R6337 vss.n15408 vss.n15407 57.894
R6338 vss.n15429 vss.n15428 57.894
R6339 vss.n15644 vss.n15643 57.894
R6340 vss.n15665 vss.n15664 57.894
R6341 vss.n15870 vss.n15869 57.894
R6342 vss.n16355 vss.n16354 57.894
R6343 vss.n16376 vss.n16375 57.894
R6344 vss.n16591 vss.n16590 57.894
R6345 vss.n16612 vss.n16611 57.894
R6346 vss.n14276 vss.n14275 57.516
R6347 vss.n11041 vss.n11040 57.516
R6348 vss.n12527 vss.n12526 57.516
R6349 vss.n13227 vss.n13226 57.516
R6350 vss.n22701 vss.n22700 57.142
R6351 vss.n22684 vss.n22683 57.142
R6352 vss.n22493 vss.n22492 57.142
R6353 vss.n22476 vss.n22475 57.142
R6354 vss.n22285 vss.n22284 57.142
R6355 vss.n22268 vss.n22267 57.142
R6356 vss.n22075 vss.n22074 57.142
R6357 vss.n21598 vss.n21597 57.142
R6358 vss.n21421 vss.n21420 57.142
R6359 vss.n21404 vss.n21403 57.142
R6360 vss.n21213 vss.n21212 57.142
R6361 vss.n21196 vss.n21195 57.142
R6362 vss.n21005 vss.n21004 57.142
R6363 vss.n20988 vss.n20987 57.142
R6364 vss.n8864 vss.n8863 57.142
R6365 vss.n8847 vss.n8846 57.142
R6366 vss.n8656 vss.n8655 57.142
R6367 vss.n8639 vss.n8638 57.142
R6368 vss.n8448 vss.n8447 57.142
R6369 vss.n8431 vss.n8430 57.142
R6370 vss.n8235 vss.n8234 57.142
R6371 vss.n8224 vss.n8223 57.142
R6372 vss.n8032 vss.n8031 57.142
R6373 vss.n8015 vss.n8014 57.142
R6374 vss.n7823 vss.n7822 57.142
R6375 vss.n7806 vss.n7805 57.142
R6376 vss.n7615 vss.n7614 57.142
R6377 vss.n7598 vss.n7597 57.142
R6378 vss.n20481 vss.n20479 55.52
R6379 vss.n20602 vss.n20600 55.52
R6380 vss.n20710 vss.n20708 55.52
R6381 vss.n20825 vss.n20823 55.52
R6382 vss.n7091 vss.n7089 55.52
R6383 vss.n7212 vss.n7210 55.52
R6384 vss.n7320 vss.n7318 55.52
R6385 vss.n7435 vss.n7433 55.52
R6386 vss.n1704 vss.n1702 55.52
R6387 vss.n1823 vss.n1821 55.52
R6388 vss.n1935 vss.n1932 55.52
R6389 vss.n1968 vss.t75 55.52
R6390 vss.n2064 vss.n2061 55.52
R6391 vss.n2179 vss.n2176 55.52
R6392 vss.n2309 vss.n2306 55.52
R6393 vss.n2424 vss.n2421 55.52
R6394 vss.n2553 vss.n2550 55.52
R6395 vss.n2668 vss.n2665 55.52
R6396 vss.n2797 vss.n2794 55.52
R6397 vss.n2906 vss.n2903 55.52
R6398 vss.n3036 vss.n3033 55.52
R6399 vss.n3151 vss.n3148 55.52
R6400 vss.n3249 vss.t41 55.52
R6401 vss.n3280 vss.n3277 55.52
R6402 vss.n3391 vss.n3389 55.52
R6403 vss.n15164 vss.n15162 55.52
R6404 vss.n165 vss.n163 55.52
R6405 vss.n284 vss.n282 55.52
R6406 vss.n396 vss.n393 55.52
R6407 vss.n429 vss.t261 55.52
R6408 vss.n525 vss.n522 55.52
R6409 vss.n640 vss.n637 55.52
R6410 vss.n770 vss.n767 55.52
R6411 vss.n885 vss.n882 55.52
R6412 vss.n1014 vss.n1011 55.52
R6413 vss.n1129 vss.n1126 55.52
R6414 vss.n1258 vss.n1255 55.52
R6415 vss.n23353 vss.n23350 55.52
R6416 vss.n23224 vss.n23221 55.52
R6417 vss.n23109 vss.n23106 55.52
R6418 vss.n23013 vss.t273 55.52
R6419 vss.n22980 vss.n22977 55.52
R6420 vss.n22868 vss.n22866 55.52
R6421 vss.n22798 vss.n22796 55.52
R6422 vss.t170 vss.n14174 52.79
R6423 vss.t174 vss.n11231 52.79
R6424 vss.t174 vss.n11230 52.79
R6425 vss.n10865 vss.n10860 52.79
R6426 vss.t172 vss.n12439 52.79
R6427 vss.t172 vss.n12440 52.79
R6428 vss.t168 vss.n13203 52.79
R6429 vss.t198 vss.n12954 52.79
R6430 vss.t198 vss.n12955 52.79
R6431 vss.t168 vss.n13204 52.79
R6432 vss.t110 vss.n10861 52.79
R6433 vss.t176 vss.n13057 52.79
R6434 vss.t147 vss.n12783 52.79
R6435 vss.t166 vss.n14016 52.79
R6436 vss.t166 vss.n14017 52.79
R6437 vss.n17520 vss.n17519 52.689
R6438 vss.n17508 vss.n17507 52.689
R6439 vss.n4130 vss.n4129 52.689
R6440 vss.n4118 vss.n4117 52.689
R6441 vss.n1642 vss.n1641 52.689
R6442 vss.n1630 vss.n1629 52.689
R6443 vss.n1615 vss.n1614 52.689
R6444 vss.n1603 vss.n1602 52.689
R6445 vss.n1590 vss.n1589 52.689
R6446 vss.n1578 vss.n1577 52.689
R6447 vss.n1565 vss.n1564 52.689
R6448 vss.n1552 vss.n1551 52.689
R6449 vss.n1532 vss.n1531 52.689
R6450 vss.n1520 vss.n1519 52.689
R6451 vss.n1507 vss.n1506 52.689
R6452 vss.n1495 vss.n1494 52.689
R6453 vss.n1480 vss.n1479 52.689
R6454 vss.n1468 vss.n1467 52.689
R6455 vss.n103 vss.n102 52.689
R6456 vss.n91 vss.n90 52.689
R6457 vss.n76 vss.n75 52.689
R6458 vss.n64 vss.n63 52.689
R6459 vss.n51 vss.n50 52.689
R6460 vss.n39 vss.n38 52.689
R6461 vss.n26 vss.n25 52.689
R6462 vss.n13 vss.n12 52.689
R6463 vss.n1315 vss.n1314 52.689
R6464 vss.n1327 vss.n1326 52.689
R6465 vss.n1341 vss.n1340 52.689
R6466 vss.n1353 vss.n1352 52.689
R6467 vss.n1368 vss.n1367 52.689
R6468 vss.n1380 vss.n1379 52.689
R6469 vss.n12186 vss.n12183 52.147
R6470 vss.n10856 vss.n10853 52.147
R6471 vss.n11299 vss.n11296 52.147
R6472 vss.n11160 vss.n11157 52.147
R6473 vss.n14298 vss.n14295 52.147
R6474 vss.n14011 vss.n14008 52.147
R6475 vss.n11800 vss.n11797 52.147
R6476 vss.n11084 vss.n11081 52.147
R6477 vss.n14788 vss.n14785 52.147
R6478 vss.n13532 vss.n13529 52.147
R6479 vss.n14523 vss.n14520 52.147
R6480 vss.n14241 vss.n14238 52.147
R6481 vss.n14878 vss.n14875 52.147
R6482 vss.n12809 vss.n12808 52.147
R6483 vss.n12689 vss.n12686 52.147
R6484 vss.n12553 vss.n12552 52.147
R6485 vss.n12053 vss.n12052 51.162
R6486 vss.n12043 vss.n12042 51.162
R6487 vss.n10972 vss.n10971 51.162
R6488 vss.n10982 vss.n10981 51.162
R6489 vss.n13835 vss.n13834 51.162
R6490 vss.n13825 vss.n13824 51.162
R6491 vss.n11127 vss.n11126 51.162
R6492 vss.n11117 vss.n11116 51.162
R6493 vss.n13366 vss.n13365 51.162
R6494 vss.n13386 vss.n13385 51.162
R6495 vss.n14198 vss.n14197 51.162
R6496 vss.n14208 vss.n14207 51.162
R6497 vss.n12891 vss.n12890 51.162
R6498 vss.n12882 vss.n12881 51.162
R6499 vss.n12482 vss.n12481 51.162
R6500 vss.n12473 vss.n12472 51.162
R6501 vss.n20532 vss.n20524 49.396
R6502 vss.n20559 vss.n20552 49.396
R6503 vss.n20761 vss.n20753 49.396
R6504 vss.n20781 vss.n20774 49.396
R6505 vss.n7142 vss.n7134 49.396
R6506 vss.n7169 vss.n7162 49.396
R6507 vss.n7371 vss.n7363 49.396
R6508 vss.n7391 vss.n7384 49.396
R6509 vss.n1758 vss.n1750 49.396
R6510 vss.n1778 vss.n1771 49.396
R6511 vss.n1989 vss.n1979 49.396
R6512 vss.n2018 vss.n2009 49.396
R6513 vss.n2234 vss.n2224 49.396
R6514 vss.n2262 vss.n2253 49.396
R6515 vss.n2478 vss.n2468 49.396
R6516 vss.n2506 vss.n2497 49.396
R6517 vss.n2723 vss.n2713 49.396
R6518 vss.n2751 vss.n2742 49.396
R6519 vss.n2961 vss.n2951 49.396
R6520 vss.n2989 vss.n2980 49.396
R6521 vss.n3205 vss.n3195 49.396
R6522 vss.n3234 vss.n3225 49.396
R6523 vss.n15207 vss.n15199 49.396
R6524 vss.n15187 vss.n15180 49.396
R6525 vss.n219 vss.n211 49.396
R6526 vss.n239 vss.n232 49.396
R6527 vss.n450 vss.n440 49.396
R6528 vss.n479 vss.n470 49.396
R6529 vss.n695 vss.n685 49.396
R6530 vss.n723 vss.n714 49.396
R6531 vss.n939 vss.n929 49.396
R6532 vss.n967 vss.n958 49.396
R6533 vss.n1184 vss.n1174 49.396
R6534 vss.n1212 vss.n1203 49.396
R6535 vss.n23307 vss.n23297 49.396
R6536 vss.n23279 vss.n23270 49.396
R6537 vss.n23063 vss.n23053 49.396
R6538 vss.n23034 vss.n23025 49.396
R6539 vss.n1400 vss.n1392 49.396
R6540 vss.n22821 vss.n22814 49.396
R6541 vss.n20467 vss.n20466 48.58
R6542 vss.n20618 vss.n20617 48.58
R6543 vss.n20696 vss.n20695 48.58
R6544 vss.n20841 vss.n20840 48.58
R6545 vss.n7077 vss.n7076 48.58
R6546 vss.n7228 vss.n7227 48.58
R6547 vss.n7306 vss.n7305 48.58
R6548 vss.n7451 vss.n7450 48.58
R6549 vss.n1690 vss.n1689 48.58
R6550 vss.t136 vss.n1719 48.58
R6551 vss.n1772 vss.t101 48.58
R6552 vss.n1839 vss.n1838 48.58
R6553 vss.n1920 vss.n1919 48.58
R6554 vss.n2081 vss.n2080 48.58
R6555 vss.n2164 vss.n2163 48.58
R6556 vss.n2326 vss.n2325 48.58
R6557 vss.n2409 vss.n2408 48.58
R6558 vss.n2570 vss.n2569 48.58
R6559 vss.n2653 vss.n2652 48.58
R6560 vss.n2813 vss.n2812 48.58
R6561 vss.n2891 vss.n2890 48.58
R6562 vss.n3053 vss.n3052 48.58
R6563 vss.n3136 vss.n3135 48.58
R6564 vss.n3297 vss.n3296 48.58
R6565 vss.n3377 vss.n3376 48.58
R6566 vss.n15205 vss.t203 48.58
R6567 vss.t88 vss.n3473 48.58
R6568 vss.n3486 vss.n3485 48.58
R6569 vss.n151 vss.n150 48.58
R6570 vss.t188 vss.n180 48.58
R6571 vss.n233 vss.t117 48.58
R6572 vss.n300 vss.n299 48.58
R6573 vss.n381 vss.n380 48.58
R6574 vss.n542 vss.n541 48.58
R6575 vss.n625 vss.n624 48.58
R6576 vss.n787 vss.n786 48.58
R6577 vss.n870 vss.n869 48.58
R6578 vss.n1031 vss.n1030 48.58
R6579 vss.n1114 vss.n1113 48.58
R6580 vss.n1275 vss.n1274 48.58
R6581 vss.n23370 vss.n23369 48.58
R6582 vss.n23209 vss.n23208 48.58
R6583 vss.n23126 vss.n23125 48.58
R6584 vss.n22965 vss.n22964 48.58
R6585 vss.n22884 vss.n22883 48.58
R6586 vss.n1398 vss.t106 48.58
R6587 vss.t97 vss.n1448 48.58
R6588 vss.n1461 vss.n1460 48.58
R6589 vss.n12183 vss.n12182 46.352
R6590 vss.n10853 vss.n10852 46.352
R6591 vss.n11296 vss.n11295 46.352
R6592 vss.n11157 vss.n11156 46.352
R6593 vss.n14295 vss.n14294 46.352
R6594 vss.n14008 vss.n14007 46.352
R6595 vss.n11797 vss.n11796 46.352
R6596 vss.n11081 vss.n11080 46.352
R6597 vss.n14785 vss.n14784 46.352
R6598 vss.n13529 vss.n13528 46.352
R6599 vss.n14520 vss.n14519 46.352
R6600 vss.n14238 vss.n14237 46.352
R6601 vss.n14875 vss.n14874 46.352
R6602 vss.n12811 vss.n12809 46.352
R6603 vss.n12686 vss.n12685 46.352
R6604 vss.n12555 vss.n12553 46.352
R6605 vss.n20644 vss.n20643 46.103
R6606 vss.n20662 vss.n20661 46.103
R6607 vss.n7254 vss.n7253 46.103
R6608 vss.n7272 vss.n7271 46.103
R6609 vss.n1865 vss.n1864 46.103
R6610 vss.n1883 vss.n1882 46.103
R6611 vss.n2109 vss.n2108 46.103
R6612 vss.n2127 vss.n2126 46.103
R6613 vss.n2353 vss.n2352 46.103
R6614 vss.n2371 vss.n2370 46.103
R6615 vss.n2597 vss.n2596 46.103
R6616 vss.n2616 vss.n2615 46.103
R6617 vss.n2836 vss.n2835 46.103
R6618 vss.n2854 vss.n2853 46.103
R6619 vss.n3080 vss.n3079 46.103
R6620 vss.n3098 vss.n3097 46.103
R6621 vss.n3324 vss.n3323 46.103
R6622 vss.n3343 vss.n3342 46.103
R6623 vss.n326 vss.n325 46.103
R6624 vss.n344 vss.n343 46.103
R6625 vss.n570 vss.n569 46.103
R6626 vss.n588 vss.n587 46.103
R6627 vss.n814 vss.n813 46.103
R6628 vss.n832 vss.n831 46.103
R6629 vss.n1058 vss.n1057 46.103
R6630 vss.n1077 vss.n1076 46.103
R6631 vss.n1303 vss.n1302 46.103
R6632 vss.n23397 vss.n23396 46.103
R6633 vss.n23172 vss.n23171 46.103
R6634 vss.n23154 vss.n23153 46.103
R6635 vss.n22928 vss.n22927 46.103
R6636 vss.n22910 vss.n22909 46.103
R6637 vss.n20514 vss.n20509 42.81
R6638 vss.n20574 vss.n20569 42.81
R6639 vss.n20742 vss.n20737 42.81
R6640 vss.n20796 vss.n20791 42.81
R6641 vss.n7124 vss.n7119 42.81
R6642 vss.n7184 vss.n7179 42.81
R6643 vss.n7352 vss.n7347 42.81
R6644 vss.n7406 vss.n7401 42.81
R6645 vss.n1736 vss.n1731 42.81
R6646 vss.n1795 vss.n1790 42.81
R6647 vss.n1969 vss.n1963 42.81
R6648 vss.n2034 vss.n2028 42.81
R6649 vss.n2214 vss.n2208 42.81
R6650 vss.n2278 vss.n2272 42.81
R6651 vss.n2458 vss.n2452 42.81
R6652 vss.n2523 vss.n2517 42.81
R6653 vss.n2702 vss.n2696 42.81
R6654 vss.n2767 vss.n2761 42.81
R6655 vss.n2941 vss.n2935 42.81
R6656 vss.n3005 vss.n2999 42.81
R6657 vss.n3185 vss.n3179 42.81
R6658 vss.n3250 vss.n3244 42.81
R6659 vss.n3423 vss.n3418 42.81
R6660 vss.n3464 vss.n3459 42.81
R6661 vss.n197 vss.n192 42.81
R6662 vss.n256 vss.n251 42.81
R6663 vss.n430 vss.n424 42.81
R6664 vss.n495 vss.n489 42.81
R6665 vss.n675 vss.n669 42.81
R6666 vss.n739 vss.n733 42.81
R6667 vss.n919 vss.n913 42.81
R6668 vss.n984 vss.n978 42.81
R6669 vss.n1163 vss.n1157 42.81
R6670 vss.n1228 vss.n1222 42.81
R6671 vss.n23323 vss.n23317 42.81
R6672 vss.n23259 vss.n23253 42.81
R6673 vss.n23079 vss.n23073 42.81
R6674 vss.n23014 vss.n23008 42.81
R6675 vss.n22838 vss.n22833 42.81
R6676 vss.n1439 vss.n1434 42.81
R6677 vss.n20482 vss.t158 41.64
R6678 vss.n20496 vss.n20494 41.64
R6679 vss.n20587 vss.n20585 41.64
R6680 vss.n20725 vss.n20723 41.64
R6681 vss.n20810 vss.n20808 41.64
R6682 vss.n20826 vss.t163 41.64
R6683 vss.n7092 vss.t179 41.64
R6684 vss.n7106 vss.n7104 41.64
R6685 vss.n7197 vss.n7195 41.64
R6686 vss.n7335 vss.n7333 41.64
R6687 vss.n7420 vss.n7418 41.64
R6688 vss.n7436 vss.t208 41.64
R6689 vss.n1719 vss.n1717 41.64
R6690 vss.n1808 vss.n1806 41.64
R6691 vss.n1951 vss.n1948 41.64
R6692 vss.n2017 vss.t21 41.64
R6693 vss.n2048 vss.n2045 41.64
R6694 vss.n2196 vss.n2193 41.64
R6695 vss.n2292 vss.n2289 41.64
R6696 vss.n2425 vss.t19 41.64
R6697 vss.n2440 vss.n2437 41.64
R6698 vss.n2537 vss.n2534 41.64
R6699 vss.n2684 vss.n2681 41.64
R6700 vss.n2781 vss.n2778 41.64
R6701 vss.n2798 vss.t39 41.64
R6702 vss.n2923 vss.n2920 41.64
R6703 vss.n3020 vss.n3017 41.64
R6704 vss.n3167 vss.n3164 41.64
R6705 vss.n3204 vss.t37 41.64
R6706 vss.n3264 vss.n3261 41.64
R6707 vss.n3406 vss.n3404 41.64
R6708 vss.n3473 vss.n3471 41.64
R6709 vss.n180 vss.n178 41.64
R6710 vss.n269 vss.n267 41.64
R6711 vss.n412 vss.n409 41.64
R6712 vss.n478 vss.t275 41.64
R6713 vss.n509 vss.n506 41.64
R6714 vss.n657 vss.n654 41.64
R6715 vss.n753 vss.n750 41.64
R6716 vss.n886 vss.t271 41.64
R6717 vss.n901 vss.n898 41.64
R6718 vss.n998 vss.n995 41.64
R6719 vss.n1145 vss.n1142 41.64
R6720 vss.n1242 vss.n1239 41.64
R6721 vss.n1259 vss.t247 41.64
R6722 vss.n23337 vss.n23334 41.64
R6723 vss.n23240 vss.n23237 41.64
R6724 vss.n23093 vss.n23090 41.64
R6725 vss.n23062 vss.t245 41.64
R6726 vss.n22996 vss.n22993 41.64
R6727 vss.n22853 vss.n22851 41.64
R6728 vss.n1448 vss.n1446 41.64
R6729 vss.n12200 vss.n12197 40.558
R6730 vss.n12004 vss.n12001 40.558
R6731 vss.n11283 vss.n11280 40.558
R6732 vss.n11181 vss.n11178 40.558
R6733 vss.n13880 vss.n13877 40.558
R6734 vss.n13990 vss.n13987 40.558
R6735 vss.n11784 vss.n11781 40.558
R6736 vss.n11094 vss.n11091 40.558
R6737 vss.n14774 vss.n14771 40.558
R6738 vss.n13515 vss.n13512 40.558
R6739 vss.n14507 vss.n14504 40.558
R6740 vss.n14221 vss.n14218 40.558
R6741 vss.n12841 vss.n12838 40.558
R6742 vss.n12814 vss.n12805 40.558
R6743 vss.n12672 vss.n12669 40.558
R6744 vss.n12558 vss.n12549 40.558
R6745 vss.n20447 vss.n20446 39.517
R6746 vss.n20629 vss.n20628 39.517
R6747 vss.n20677 vss.n20676 39.517
R6748 vss.n20853 vss.n20852 39.517
R6749 vss.n7057 vss.n7056 39.517
R6750 vss.n7239 vss.n7238 39.517
R6751 vss.n7287 vss.n7286 39.517
R6752 vss.n7463 vss.n7462 39.517
R6753 vss.n1850 vss.n1849 39.517
R6754 vss.n1899 vss.n1898 39.517
R6755 vss.n2092 vss.n2091 39.517
R6756 vss.n2143 vss.n2142 39.517
R6757 vss.n2337 vss.n2336 39.517
R6758 vss.n2387 vss.n2386 39.517
R6759 vss.n2581 vss.n2580 39.517
R6760 vss.n2632 vss.n2631 39.517
R6761 vss.n2824 vss.n2823 39.517
R6762 vss.n2870 vss.n2869 39.517
R6763 vss.n3064 vss.n3063 39.517
R6764 vss.n3115 vss.n3114 39.517
R6765 vss.n3308 vss.n3307 39.517
R6766 vss.n3358 vss.n3357 39.517
R6767 vss.n311 vss.n310 39.517
R6768 vss.n360 vss.n359 39.517
R6769 vss.n553 vss.n552 39.517
R6770 vss.n604 vss.n603 39.517
R6771 vss.n798 vss.n797 39.517
R6772 vss.n848 vss.n847 39.517
R6773 vss.n1042 vss.n1041 39.517
R6774 vss.n1093 vss.n1092 39.517
R6775 vss.n1287 vss.n1286 39.517
R6776 vss.n23381 vss.n23380 39.517
R6777 vss.n23188 vss.n23187 39.517
R6778 vss.n23137 vss.n23136 39.517
R6779 vss.n22944 vss.n22943 39.517
R6780 vss.n22895 vss.n22894 39.517
R6781 vss.n3429 vss.t202 39.079
R6782 vss.n1404 vss.t105 39.079
R6783 vss.n1653 vss.t100 39.078
R6784 vss.n114 vss.t116 39.078
R6785 vss.n3429 vss.t87 39.075
R6786 vss.n1404 vss.t96 39.075
R6787 vss.n17531 vss.t152 39.067
R6788 vss.n4141 vss.t91 39.067
R6789 vss.n17486 vss.t130 39.061
R6790 vss.n4096 vss.t125 39.061
R6791 vss.n1743 vss.t135 39.06
R6792 vss.n204 vss.t187 39.06
R6793 vss.n17486 vss.t162 39.048
R6794 vss.n4096 vss.t207 39.048
R6795 vss.n17531 vss.t157 39.037
R6796 vss.n4141 vss.t178 39.037
R6797 vss.n20498 vss.n20493 36.224
R6798 vss.n20589 vss.n20584 36.224
R6799 vss.n20727 vss.n20722 36.224
R6800 vss.n20812 vss.n20807 36.224
R6801 vss.n7108 vss.n7103 36.224
R6802 vss.n7199 vss.n7194 36.224
R6803 vss.n7337 vss.n7332 36.224
R6804 vss.n7422 vss.n7417 36.224
R6805 vss.n1721 vss.n1716 36.224
R6806 vss.n1810 vss.n1805 36.224
R6807 vss.n1953 vss.n1947 36.224
R6808 vss.n2050 vss.n2044 36.224
R6809 vss.n2198 vss.n2192 36.224
R6810 vss.n2294 vss.n2288 36.224
R6811 vss.n2442 vss.n2436 36.224
R6812 vss.n2539 vss.n2533 36.224
R6813 vss.n2686 vss.n2680 36.224
R6814 vss.n2783 vss.n2777 36.224
R6815 vss.n2925 vss.n2919 36.224
R6816 vss.n3022 vss.n3016 36.224
R6817 vss.n3169 vss.n3163 36.224
R6818 vss.n3266 vss.n3260 36.224
R6819 vss.n3408 vss.n3403 36.224
R6820 vss.n3475 vss.n3470 36.224
R6821 vss.n182 vss.n177 36.224
R6822 vss.n271 vss.n266 36.224
R6823 vss.n414 vss.n408 36.224
R6824 vss.n511 vss.n505 36.224
R6825 vss.n659 vss.n653 36.224
R6826 vss.n755 vss.n749 36.224
R6827 vss.n903 vss.n897 36.224
R6828 vss.n1000 vss.n994 36.224
R6829 vss.n1147 vss.n1141 36.224
R6830 vss.n1244 vss.n1238 36.224
R6831 vss.n23339 vss.n23333 36.224
R6832 vss.n23242 vss.n23236 36.224
R6833 vss.n23095 vss.n23089 36.224
R6834 vss.n22998 vss.n22992 36.224
R6835 vss.n22855 vss.n22850 36.224
R6836 vss.n1450 vss.n1445 36.224
R6837 vss.n21838 vss.t142 35.379
R6838 vss.n21728 vss.n21691 35.379
R6839 vss.n21731 vss.n21691 35.379
R6840 vss.n3787 vss.t151 35.379
R6841 vss.n3677 vss.n3640 35.379
R6842 vss.n3680 vss.n3640 35.379
R6843 vss.n12169 vss.n12168 34.764
R6844 vss.n11987 vss.n11986 34.764
R6845 vss.n11321 vss.n11320 34.764
R6846 vss.n14309 vss.n14308 34.764
R6847 vss.n11609 vss.n11608 34.764
R6848 vss.n11822 vss.n11821 34.764
R6849 vss.n14799 vss.n14798 34.764
R6850 vss.n14626 vss.n14625 34.764
R6851 vss.n14537 vss.n14536 34.764
R6852 vss.n14258 vss.n14257 34.764
R6853 vss.n14890 vss.n14889 34.764
R6854 vss.n15046 vss.n15045 34.764
R6855 vss.n12702 vss.n12701 34.764
R6856 vss.n20451 vss.n20450 34.7
R6857 vss.n20633 vss.n20632 34.7
R6858 vss.n20681 vss.n20680 34.7
R6859 vss.n20857 vss.n20856 34.7
R6860 vss.n7061 vss.n7060 34.7
R6861 vss.n7243 vss.n7242 34.7
R6862 vss.n7291 vss.n7290 34.7
R6863 vss.n7467 vss.n7466 34.7
R6864 vss.n1854 vss.n1853 34.7
R6865 vss.n1904 vss.n1903 34.7
R6866 vss.t75 vss.n1967 34.7
R6867 vss.n2097 vss.n2096 34.7
R6868 vss.n2148 vss.n2147 34.7
R6869 vss.n2342 vss.n2341 34.7
R6870 vss.n2392 vss.n2391 34.7
R6871 vss.n2586 vss.n2585 34.7
R6872 vss.n2637 vss.n2636 34.7
R6873 vss.n2828 vss.n2827 34.7
R6874 vss.n2875 vss.n2874 34.7
R6875 vss.n3069 vss.n3068 34.7
R6876 vss.n3120 vss.n3119 34.7
R6877 vss.t41 vss.n3248 34.7
R6878 vss.n3313 vss.n3312 34.7
R6879 vss.n3362 vss.n3361 34.7
R6880 vss.n315 vss.n314 34.7
R6881 vss.n365 vss.n364 34.7
R6882 vss.t261 vss.n428 34.7
R6883 vss.n558 vss.n557 34.7
R6884 vss.n609 vss.n608 34.7
R6885 vss.n803 vss.n802 34.7
R6886 vss.n853 vss.n852 34.7
R6887 vss.n1047 vss.n1046 34.7
R6888 vss.n1098 vss.n1097 34.7
R6889 vss.n1292 vss.n1291 34.7
R6890 vss.n23386 vss.n23385 34.7
R6891 vss.n23193 vss.n23192 34.7
R6892 vss.n23142 vss.n23141 34.7
R6893 vss.t273 vss.n23012 34.7
R6894 vss.n22949 vss.n22948 34.7
R6895 vss.n22899 vss.n22898 34.7
R6896 vss.n11813 vss.n11812 34.645
R6897 vss.n15002 vss.n15001 34.645
R6898 vss.n12400 vss.n12399 34.645
R6899 vss.n14710 vss.n14709 34.645
R6900 vss.n13447 vss.n13446 34.645
R6901 vss.n13022 vss.n13021 34.645
R6902 vss.n10579 vss.n10578 34.645
R6903 vss.n10736 vss.n10735 34.645
R6904 vss.n12032 vss.n12031 34.645
R6905 vss.n14574 vss.n14573 34.645
R6906 vss.n13634 vss.n13633 34.645
R6907 vss.n13686 vss.n13685 34.645
R6908 vss.n11383 vss.n11382 34.645
R6909 vss.n11369 vss.n11368 34.645
R6910 vss.n11312 vss.n11311 34.645
R6911 vss.n13960 vss.n13959 34.645
R6912 vss.n16249 vss.n16248 33.624
R6913 vss.n16672 vss.n16671 33.624
R6914 vss.n16899 vss.n16896 33.49
R6915 vss.n17135 vss.n17132 33.49
R6916 vss.n15944 vss.n15941 33.49
R6917 vss.n16180 vss.n16177 33.49
R6918 vss.n15420 vss.n15417 33.49
R6919 vss.n15656 vss.n15653 33.49
R6920 vss.n16367 vss.n16364 33.49
R6921 vss.n16603 vss.n16600 33.49
R6922 vss.n21859 vss.n21858 33.413
R6923 vss.n3808 vss.n3807 33.413
R6924 vss.n20463 vss.n20462 32.931
R6925 vss.n20614 vss.n20613 32.931
R6926 vss.n20692 vss.n20691 32.931
R6927 vss.n20837 vss.n20836 32.931
R6928 vss.n7073 vss.n7072 32.931
R6929 vss.n7224 vss.n7223 32.931
R6930 vss.n7302 vss.n7301 32.931
R6931 vss.n7447 vss.n7446 32.931
R6932 vss.n1686 vss.n1685 32.931
R6933 vss.n1835 vss.n1834 32.931
R6934 vss.n1915 vss.n1914 32.931
R6935 vss.n2076 vss.n2075 32.931
R6936 vss.n2159 vss.n2158 32.931
R6937 vss.n2321 vss.n2320 32.931
R6938 vss.n2404 vss.n2403 32.931
R6939 vss.n2565 vss.n2564 32.931
R6940 vss.n2648 vss.n2647 32.931
R6941 vss.n2809 vss.n2808 32.931
R6942 vss.n2886 vss.n2885 32.931
R6943 vss.n3048 vss.n3047 32.931
R6944 vss.n3131 vss.n3130 32.931
R6945 vss.n3292 vss.n3291 32.931
R6946 vss.n3373 vss.n3372 32.931
R6947 vss.n3482 vss.n3481 32.931
R6948 vss.n147 vss.n146 32.931
R6949 vss.n296 vss.n295 32.931
R6950 vss.n376 vss.n375 32.931
R6951 vss.n537 vss.n536 32.931
R6952 vss.n620 vss.n619 32.931
R6953 vss.n782 vss.n781 32.931
R6954 vss.n865 vss.n864 32.931
R6955 vss.n1026 vss.n1025 32.931
R6956 vss.n1109 vss.n1108 32.931
R6957 vss.n1270 vss.n1269 32.931
R6958 vss.n23365 vss.n23364 32.931
R6959 vss.n23204 vss.n23203 32.931
R6960 vss.n23121 vss.n23120 32.931
R6961 vss.n22960 vss.n22959 32.931
R6962 vss.n22880 vss.n22879 32.931
R6963 vss.n1457 vss.n1456 32.931
R6964 vss.n9272 vss.n9269 31.623
R6965 vss.n18953 vss.n17681 31.52
R6966 vss.n18946 vss.n17688 31.52
R6967 vss.n18830 vss.n17786 31.52
R6968 vss.n18826 vss.n17790 31.52
R6969 vss.n18713 vss.n17890 31.52
R6970 vss.n18705 vss.n17900 31.52
R6971 vss.n18589 vss.n17999 31.52
R6972 vss.n18585 vss.n18003 31.52
R6973 vss.n18472 vss.n18103 31.52
R6974 vss.n18464 vss.n18113 31.52
R6975 vss.n18348 vss.n18212 31.52
R6976 vss.n18344 vss.n18216 31.52
R6977 vss.n20223 vss.n19086 31.52
R6978 vss.n20219 vss.n19090 31.52
R6979 vss.n20099 vss.n19188 31.52
R6980 vss.n20092 vss.n19195 31.52
R6981 vss.n19976 vss.n19293 31.52
R6982 vss.n19972 vss.n19297 31.52
R6983 vss.n19852 vss.n19395 31.52
R6984 vss.n19845 vss.n19401 31.52
R6985 vss.n19729 vss.n19500 31.52
R6986 vss.n19725 vss.n19504 31.52
R6987 vss.n20357 vss.n17592 31.52
R6988 vss.n20353 vss.n20352 31.52
R6989 vss.n5563 vss.n4291 31.52
R6990 vss.n5556 vss.n4298 31.52
R6991 vss.n5440 vss.n4396 31.52
R6992 vss.n5436 vss.n4400 31.52
R6993 vss.n5323 vss.n4500 31.52
R6994 vss.n5315 vss.n4510 31.52
R6995 vss.n5199 vss.n4609 31.52
R6996 vss.n5195 vss.n4613 31.52
R6997 vss.n5082 vss.n4713 31.52
R6998 vss.n5074 vss.n4723 31.52
R6999 vss.n4958 vss.n4822 31.52
R7000 vss.n4954 vss.n4826 31.52
R7001 vss.n6833 vss.n5696 31.52
R7002 vss.n6829 vss.n5700 31.52
R7003 vss.n6709 vss.n5798 31.52
R7004 vss.n6702 vss.n5805 31.52
R7005 vss.n6586 vss.n5903 31.52
R7006 vss.n6582 vss.n5907 31.52
R7007 vss.n6462 vss.n6005 31.52
R7008 vss.n6455 vss.n6011 31.52
R7009 vss.n6339 vss.n6110 31.52
R7010 vss.n6335 vss.n6114 31.52
R7011 vss.n6967 vss.n4202 31.52
R7012 vss.n6963 vss.n6962 31.52
R7013 vss.n16776 vss.n16772 31.52
R7014 vss.n16794 vss.n16790 31.52
R7015 vss.n17008 vss.n17004 31.52
R7016 vss.n17025 vss.n17021 31.52
R7017 vss.n17244 vss.n17240 31.52
R7018 vss.n17263 vss.n17259 31.52
R7019 vss.n16055 vss.n16053 31.52
R7020 vss.n16071 vss.n16069 31.52
R7021 vss.n15237 vss.n15231 31.52
R7022 vss.n15320 vss.n15316 31.52
R7023 vss.n15528 vss.n15524 31.52
R7024 vss.n15545 vss.n15541 31.52
R7025 vss.n15764 vss.n15760 31.52
R7026 vss.n15779 vss.n15775 31.52
R7027 vss.n16475 vss.n16471 31.52
R7028 vss.n16492 vss.n16488 31.52
R7029 vss.n21832 vss.n21831 31.448
R7030 vss.n21839 vss.n21838 31.448
R7031 vss.n21728 vss.n21727 31.448
R7032 vss.n21732 vss.n21731 31.448
R7033 vss.n3781 vss.n3780 31.448
R7034 vss.n3788 vss.n3787 31.448
R7035 vss.n3677 vss.n3676 31.448
R7036 vss.n3681 vss.n3680 31.448
R7037 vss.n17335 vss.n17334 30.901
R7038 vss.n17346 vss.n17345 30.901
R7039 vss.n17357 vss.n17356 30.901
R7040 vss.n17368 vss.n17367 30.901
R7041 vss.n17379 vss.n17378 30.901
R7042 vss.n17390 vss.n17389 30.901
R7043 vss.n17412 vss.n17411 30.901
R7044 vss.n17423 vss.n17422 30.901
R7045 vss.n17434 vss.n17433 30.901
R7046 vss.n17445 vss.n17444 30.901
R7047 vss.n17456 vss.n17455 30.901
R7048 vss.n17467 vss.n17466 30.901
R7049 vss.n17478 vss.n17477 30.901
R7050 vss.n3493 vss.n3492 30.901
R7051 vss.n3504 vss.n3503 30.901
R7052 vss.n3515 vss.n3514 30.901
R7053 vss.n3526 vss.n3525 30.901
R7054 vss.n3537 vss.n3536 30.901
R7055 vss.n3548 vss.n3547 30.901
R7056 vss.n4022 vss.n4021 30.901
R7057 vss.n4033 vss.n4032 30.901
R7058 vss.n4044 vss.n4043 30.901
R7059 vss.n4055 vss.n4054 30.901
R7060 vss.n4066 vss.n4065 30.901
R7061 vss.n4077 vss.n4076 30.901
R7062 vss.n4088 vss.n4087 30.901
R7063 vss.n20483 vss.n20478 29.637
R7064 vss.n20604 vss.n20599 29.637
R7065 vss.n20712 vss.n20707 29.637
R7066 vss.n20827 vss.n20822 29.637
R7067 vss.n7093 vss.n7088 29.637
R7068 vss.n7214 vss.n7209 29.637
R7069 vss.n7322 vss.n7317 29.637
R7070 vss.n7437 vss.n7432 29.637
R7071 vss.n1706 vss.n1701 29.637
R7072 vss.n1825 vss.n1820 29.637
R7073 vss.n1937 vss.n1931 29.637
R7074 vss.n2066 vss.n2060 29.637
R7075 vss.n2181 vss.n2175 29.637
R7076 vss.n2311 vss.n2305 29.637
R7077 vss.n2426 vss.n2420 29.637
R7078 vss.n2555 vss.n2549 29.637
R7079 vss.n2670 vss.n2664 29.637
R7080 vss.n2799 vss.n2793 29.637
R7081 vss.n2908 vss.n2902 29.637
R7082 vss.n3038 vss.n3032 29.637
R7083 vss.n3153 vss.n3147 29.637
R7084 vss.n3282 vss.n3276 29.637
R7085 vss.n3393 vss.n3388 29.637
R7086 vss.n15166 vss.n15161 29.637
R7087 vss.n167 vss.n162 29.637
R7088 vss.n286 vss.n281 29.637
R7089 vss.n398 vss.n392 29.637
R7090 vss.n527 vss.n521 29.637
R7091 vss.n642 vss.n636 29.637
R7092 vss.n772 vss.n766 29.637
R7093 vss.n887 vss.n881 29.637
R7094 vss.n1016 vss.n1010 29.637
R7095 vss.n1131 vss.n1125 29.637
R7096 vss.n1260 vss.n1254 29.637
R7097 vss.n23355 vss.n23349 29.637
R7098 vss.n23226 vss.n23220 29.637
R7099 vss.n23111 vss.n23105 29.637
R7100 vss.n22982 vss.n22976 29.637
R7101 vss.n22870 vss.n22865 29.637
R7102 vss.n22800 vss.n22795 29.637
R7103 vss.n19016 vss.n17633 29.55
R7104 vss.n19012 vss.n17637 29.55
R7105 vss.n17736 vss.n17728 29.55
R7106 vss.n18884 vss.n17737 29.55
R7107 vss.n18769 vss.n17838 29.55
R7108 vss.n17848 vss.n17846 29.55
R7109 vss.n17949 vss.n17941 29.55
R7110 vss.n18643 vss.n17950 29.55
R7111 vss.n18528 vss.n18051 29.55
R7112 vss.n18061 vss.n18059 29.55
R7113 vss.n18162 vss.n18154 29.55
R7114 vss.n18402 vss.n18163 29.55
R7115 vss.n18287 vss.n18264 29.55
R7116 vss.n18276 vss.n18272 29.55
R7117 vss.n20285 vss.n19035 29.55
R7118 vss.n20277 vss.n19037 29.55
R7119 vss.n20162 vss.n19138 29.55
R7120 vss.n20158 vss.n19144 29.55
R7121 vss.n19243 vss.n19235 29.55
R7122 vss.n20030 vss.n19244 29.55
R7123 vss.n19915 vss.n19345 29.55
R7124 vss.n19911 vss.n19351 29.55
R7125 vss.n19450 vss.n19442 29.55
R7126 vss.n19783 vss.n19451 29.55
R7127 vss.n19668 vss.n19552 29.55
R7128 vss.n19664 vss.n19558 29.55
R7129 vss.n20313 vss.n17611 29.55
R7130 vss.n20309 vss.n20302 29.55
R7131 vss.n5626 vss.n4243 29.55
R7132 vss.n5622 vss.n4247 29.55
R7133 vss.n4346 vss.n4338 29.55
R7134 vss.n5494 vss.n4347 29.55
R7135 vss.n5379 vss.n4448 29.55
R7136 vss.n4458 vss.n4456 29.55
R7137 vss.n4559 vss.n4551 29.55
R7138 vss.n5253 vss.n4560 29.55
R7139 vss.n5138 vss.n4661 29.55
R7140 vss.n4671 vss.n4669 29.55
R7141 vss.n4772 vss.n4764 29.55
R7142 vss.n5012 vss.n4773 29.55
R7143 vss.n4897 vss.n4874 29.55
R7144 vss.n4886 vss.n4882 29.55
R7145 vss.n6895 vss.n5645 29.55
R7146 vss.n6887 vss.n5647 29.55
R7147 vss.n6772 vss.n5748 29.55
R7148 vss.n6768 vss.n5754 29.55
R7149 vss.n5853 vss.n5845 29.55
R7150 vss.n6640 vss.n5854 29.55
R7151 vss.n6525 vss.n5955 29.55
R7152 vss.n6521 vss.n5961 29.55
R7153 vss.n6060 vss.n6052 29.55
R7154 vss.n6393 vss.n6061 29.55
R7155 vss.n6278 vss.n6162 29.55
R7156 vss.n6274 vss.n6168 29.55
R7157 vss.n6923 vss.n4221 29.55
R7158 vss.n6919 vss.n6912 29.55
R7159 vss.n16679 vss.n16678 29.55
R7160 vss.n16883 vss.n16882 29.55
R7161 vss.n16906 vss.n16905 29.55
R7162 vss.n17119 vss.n17118 29.55
R7163 vss.n17142 vss.n17141 29.55
R7164 vss.n16260 vss.n16259 29.55
R7165 vss.n15929 vss.n15928 29.55
R7166 vss.n15953 vss.n15952 29.55
R7167 vss.n16165 vss.n16164 29.55
R7168 vss.n16189 vss.n16188 29.55
R7169 vss.n16244 vss.n16243 29.55
R7170 vss.n16288 vss.n16287 29.55
R7171 vss.n15405 vss.n15404 29.55
R7172 vss.n15426 vss.n15425 29.55
R7173 vss.n15641 vss.n15640 29.55
R7174 vss.n15662 vss.n15661 29.55
R7175 vss.n15868 vss.n15867 29.55
R7176 vss.n16352 vss.n16351 29.55
R7177 vss.n16373 vss.n16372 29.55
R7178 vss.n16588 vss.n16587 29.55
R7179 vss.n16609 vss.n16608 29.55
R7180 vss.n16667 vss.n16666 29.55
R7181 vss.n12524 vss.n12523 29.257
R7182 vss.n13224 vss.n13223 29.257
R7183 vss.n14273 vss.n14272 29.257
R7184 vss.n11038 vss.n11037 29.257
R7185 vss.n22706 vss.n22702 28.97
R7186 vss.n22687 vss.n22685 28.97
R7187 vss.n22498 vss.n22494 28.97
R7188 vss.n22479 vss.n22477 28.97
R7189 vss.n22290 vss.n22286 28.97
R7190 vss.n22271 vss.n22269 28.97
R7191 vss.n22080 vss.n22076 28.97
R7192 vss.n21601 vss.n21599 28.97
R7193 vss.n21426 vss.n21422 28.97
R7194 vss.n21407 vss.n21405 28.97
R7195 vss.n21218 vss.n21214 28.97
R7196 vss.n21199 vss.n21197 28.97
R7197 vss.n21010 vss.n21006 28.97
R7198 vss.n20991 vss.n20989 28.97
R7199 vss.n12227 vss.n12224 28.97
R7200 vss.n12021 vss.n12018 28.97
R7201 vss.n11257 vss.n11254 28.97
R7202 vss.n11197 vss.n11194 28.97
R7203 vss.n13914 vss.n13911 28.97
R7204 vss.n14052 vss.n14049 28.97
R7205 vss.n11747 vss.n11744 28.97
R7206 vss.n11074 vss.n11071 28.97
R7207 vss.n14741 vss.n14738 28.97
R7208 vss.n14682 vss.n14679 28.97
R7209 vss.n14469 vss.n14466 28.97
R7210 vss.n14251 vss.n14248 28.97
R7211 vss.n12856 vss.n12853 28.97
R7212 vss.n12915 vss.n12914 28.97
R7213 vss.n12656 vss.n12653 28.97
R7214 vss.n12502 vss.n12501 28.97
R7215 vss.n8869 vss.n8865 28.97
R7216 vss.n8850 vss.n8848 28.97
R7217 vss.n8661 vss.n8657 28.97
R7218 vss.n8642 vss.n8640 28.97
R7219 vss.n8453 vss.n8449 28.97
R7220 vss.n8434 vss.n8432 28.97
R7221 vss.n8240 vss.n8236 28.97
R7222 vss.n8227 vss.n8225 28.97
R7223 vss.n8037 vss.n8033 28.97
R7224 vss.n8018 vss.n8016 28.97
R7225 vss.n7828 vss.n7824 28.97
R7226 vss.n7809 vss.n7807 28.97
R7227 vss.n7620 vss.n7616 28.97
R7228 vss.n7601 vss.n7599 28.97
R7229 vss.n19088 vss.n19079 28.947
R7230 vss.n19101 vss.n19089 28.947
R7231 vss.n20102 vss.n20101 28.947
R7232 vss.n20090 vss.n20089 28.947
R7233 vss.n19295 vss.n19286 28.947
R7234 vss.n19308 vss.n19296 28.947
R7235 vss.n19855 vss.n19854 28.947
R7236 vss.n19843 vss.n19842 28.947
R7237 vss.n19502 vss.n19493 28.947
R7238 vss.n19515 vss.n19503 28.947
R7239 vss.n19609 vss.n17594 28.947
R7240 vss.n20349 vss.n17595 28.947
R7241 vss.n18956 vss.n18955 28.947
R7242 vss.n18944 vss.n18943 28.947
R7243 vss.n17788 vss.n17779 28.947
R7244 vss.n17801 vss.n17789 28.947
R7245 vss.n18715 vss.n18714 28.947
R7246 vss.n18703 vss.n18702 28.947
R7247 vss.n18001 vss.n17992 28.947
R7248 vss.n18014 vss.n18002 28.947
R7249 vss.n18474 vss.n18473 28.947
R7250 vss.n18462 vss.n18461 28.947
R7251 vss.n18214 vss.n18205 28.947
R7252 vss.n18227 vss.n18215 28.947
R7253 vss.n5698 vss.n5689 28.947
R7254 vss.n5711 vss.n5699 28.947
R7255 vss.n6712 vss.n6711 28.947
R7256 vss.n6700 vss.n6699 28.947
R7257 vss.n5905 vss.n5896 28.947
R7258 vss.n5918 vss.n5906 28.947
R7259 vss.n6465 vss.n6464 28.947
R7260 vss.n6453 vss.n6452 28.947
R7261 vss.n6112 vss.n6103 28.947
R7262 vss.n6125 vss.n6113 28.947
R7263 vss.n6219 vss.n4204 28.947
R7264 vss.n6959 vss.n4205 28.947
R7265 vss.n5566 vss.n5565 28.947
R7266 vss.n5554 vss.n5553 28.947
R7267 vss.n4398 vss.n4389 28.947
R7268 vss.n4411 vss.n4399 28.947
R7269 vss.n5325 vss.n5324 28.947
R7270 vss.n5313 vss.n5312 28.947
R7271 vss.n4611 vss.n4602 28.947
R7272 vss.n4624 vss.n4612 28.947
R7273 vss.n5084 vss.n5083 28.947
R7274 vss.n5072 vss.n5071 28.947
R7275 vss.n4824 vss.n4815 28.947
R7276 vss.n4837 vss.n4825 28.947
R7277 vss.n16774 vss.n16773 28.947
R7278 vss.n16792 vss.n16791 28.947
R7279 vss.n17006 vss.n17005 28.947
R7280 vss.n17023 vss.n17022 28.947
R7281 vss.n17242 vss.n17241 28.947
R7282 vss.n17261 vss.n17260 28.947
R7283 vss.n16052 vss.n16051 28.947
R7284 vss.n16068 vss.n16067 28.947
R7285 vss.n16248 vss.n16247 28.947
R7286 vss.n15235 vss.n15234 28.947
R7287 vss.n15318 vss.n15317 28.947
R7288 vss.n15526 vss.n15525 28.947
R7289 vss.n15543 vss.n15542 28.947
R7290 vss.n15762 vss.n15761 28.947
R7291 vss.n15777 vss.n15776 28.947
R7292 vss.n16473 vss.n16472 28.947
R7293 vss.n16490 vss.n16489 28.947
R7294 vss.n16671 vss.n16670 28.947
R7295 vss.n9193 vss.t361 28.577
R7296 vss.n17338 vss.n17337 28.571
R7297 vss.n17349 vss.n17348 28.571
R7298 vss.n17360 vss.n17359 28.571
R7299 vss.n17371 vss.n17370 28.571
R7300 vss.n17382 vss.n17381 28.571
R7301 vss.n17393 vss.n17392 28.571
R7302 vss.n17415 vss.n17414 28.571
R7303 vss.n17426 vss.n17425 28.571
R7304 vss.n17437 vss.n17436 28.571
R7305 vss.n17448 vss.n17447 28.571
R7306 vss.n17459 vss.n17458 28.571
R7307 vss.n17470 vss.n17469 28.571
R7308 vss.n17481 vss.n17480 28.571
R7309 vss.n3496 vss.n3495 28.571
R7310 vss.n3507 vss.n3506 28.571
R7311 vss.n3518 vss.n3517 28.571
R7312 vss.n3529 vss.n3528 28.571
R7313 vss.n3540 vss.n3539 28.571
R7314 vss.n3551 vss.n3550 28.571
R7315 vss.n4025 vss.n4024 28.571
R7316 vss.n4036 vss.n4035 28.571
R7317 vss.n4047 vss.n4046 28.571
R7318 vss.n4058 vss.n4057 28.571
R7319 vss.n4069 vss.n4068 28.571
R7320 vss.n4080 vss.n4079 28.571
R7321 vss.n4091 vss.n4090 28.571
R7322 vss.n14177 vss.n14176 28.333
R7323 vss.n11234 vss.n11233 28.333
R7324 vss.n11709 vss.n11708 28.333
R7325 vss.n11334 vss.n11333 28.333
R7326 vss.n10868 vss.n10867 28.333
R7327 vss.n11341 vss.n11340 28.333
R7328 vss.n10765 vss.n10764 28.333
R7329 vss.n12444 vss.n12443 28.333
R7330 vss.n13050 vss.n13049 28.333
R7331 vss.n13281 vss.n13280 28.333
R7332 vss.n13393 vss.n13391 28.333
R7333 vss.n12958 vss.n12957 28.333
R7334 vss.n14147 vss.n14146 28.333
R7335 vss.n13484 vss.n13483 28.333
R7336 vss.n13722 vss.n13721 28.333
R7337 vss.n13715 vss.n13714 28.333
R7338 vss.n14022 vss.n14021 28.333
R7339 vss.n20512 vss.n20510 27.76
R7340 vss.n20572 vss.n20570 27.76
R7341 vss.n20740 vss.n20738 27.76
R7342 vss.n20794 vss.n20792 27.76
R7343 vss.n7122 vss.n7120 27.76
R7344 vss.n7182 vss.n7180 27.76
R7345 vss.n7350 vss.n7348 27.76
R7346 vss.n7404 vss.n7402 27.76
R7347 vss.n1720 vss.t136 27.76
R7348 vss.n1734 vss.n1732 27.76
R7349 vss.n1793 vss.n1791 27.76
R7350 vss.n1967 vss.n1964 27.76
R7351 vss.n2032 vss.n2029 27.76
R7352 vss.n2212 vss.n2209 27.76
R7353 vss.n2276 vss.n2273 27.76
R7354 vss.n2456 vss.n2453 27.76
R7355 vss.n2521 vss.n2518 27.76
R7356 vss.n2700 vss.n2697 27.76
R7357 vss.n2765 vss.n2762 27.76
R7358 vss.n2939 vss.n2936 27.76
R7359 vss.n3003 vss.n3000 27.76
R7360 vss.n3183 vss.n3180 27.76
R7361 vss.n3248 vss.n3245 27.76
R7362 vss.n3421 vss.n3419 27.76
R7363 vss.n3462 vss.n3460 27.76
R7364 vss.n3474 vss.t88 27.76
R7365 vss.n181 vss.t188 27.76
R7366 vss.n195 vss.n193 27.76
R7367 vss.n254 vss.n252 27.76
R7368 vss.n428 vss.n425 27.76
R7369 vss.n493 vss.n490 27.76
R7370 vss.n673 vss.n670 27.76
R7371 vss.n737 vss.n734 27.76
R7372 vss.n917 vss.n914 27.76
R7373 vss.n982 vss.n979 27.76
R7374 vss.n1161 vss.n1158 27.76
R7375 vss.n1226 vss.n1223 27.76
R7376 vss.n23321 vss.n23318 27.76
R7377 vss.n23257 vss.n23254 27.76
R7378 vss.n23077 vss.n23074 27.76
R7379 vss.n23012 vss.n23009 27.76
R7380 vss.n22836 vss.n22834 27.76
R7381 vss.n1437 vss.n1435 27.76
R7382 vss.n1449 vss.t97 27.76
R7383 vss.n18965 vss.n17674 27.58
R7384 vss.n17699 vss.n17690 27.58
R7385 vss.n18837 vss.n17778 27.58
R7386 vss.n18819 vss.n17800 27.58
R7387 vss.n18717 vss.n17886 27.58
R7388 vss.n17912 vss.n17903 27.58
R7389 vss.n18596 vss.n17991 27.58
R7390 vss.n18578 vss.n18013 27.58
R7391 vss.n18476 vss.n18099 27.58
R7392 vss.n18125 vss.n18116 27.58
R7393 vss.n18355 vss.n18204 27.58
R7394 vss.n18337 vss.n18226 27.58
R7395 vss.n20230 vss.n19078 27.58
R7396 vss.n20212 vss.n19100 27.58
R7397 vss.n20111 vss.n19181 27.58
R7398 vss.n19206 vss.n19197 27.58
R7399 vss.n19983 vss.n19285 27.58
R7400 vss.n19965 vss.n19307 27.58
R7401 vss.n19864 vss.n19388 27.58
R7402 vss.n19413 vss.n19404 27.58
R7403 vss.n19736 vss.n19492 27.58
R7404 vss.n19718 vss.n19514 27.58
R7405 vss.n19606 vss.n19595 27.58
R7406 vss.n20346 vss.n17596 27.58
R7407 vss.n5575 vss.n4284 27.58
R7408 vss.n4309 vss.n4300 27.58
R7409 vss.n5447 vss.n4388 27.58
R7410 vss.n5429 vss.n4410 27.58
R7411 vss.n5327 vss.n4496 27.58
R7412 vss.n4522 vss.n4513 27.58
R7413 vss.n5206 vss.n4601 27.58
R7414 vss.n5188 vss.n4623 27.58
R7415 vss.n5086 vss.n4709 27.58
R7416 vss.n4735 vss.n4726 27.58
R7417 vss.n4965 vss.n4814 27.58
R7418 vss.n4947 vss.n4836 27.58
R7419 vss.n6840 vss.n5688 27.58
R7420 vss.n6822 vss.n5710 27.58
R7421 vss.n6721 vss.n5791 27.58
R7422 vss.n5816 vss.n5807 27.58
R7423 vss.n6593 vss.n5895 27.58
R7424 vss.n6575 vss.n5917 27.58
R7425 vss.n6474 vss.n5998 27.58
R7426 vss.n6023 vss.n6014 27.58
R7427 vss.n6346 vss.n6102 27.58
R7428 vss.n6328 vss.n6124 27.58
R7429 vss.n6216 vss.n6205 27.58
R7430 vss.n6956 vss.n4206 27.58
R7431 vss.n16764 vss.n16760 27.58
R7432 vss.n16805 vss.n16801 27.58
R7433 vss.n16994 vss.n16990 27.58
R7434 vss.n17039 vss.n17035 27.58
R7435 vss.n17230 vss.n17226 27.58
R7436 vss.n17294 vss.n17290 27.58
R7437 vss.n16041 vss.n16039 27.58
R7438 vss.n16085 vss.n16083 27.58
R7439 vss.n15247 vss.n15243 27.58
R7440 vss.n15225 vss.n15221 27.58
R7441 vss.n15514 vss.n15510 27.58
R7442 vss.n15561 vss.n15557 27.58
R7443 vss.n15750 vss.n15746 27.58
R7444 vss.n15791 vss.n15787 27.58
R7445 vss.n16461 vss.n16457 27.58
R7446 vss.n16508 vss.n16504 27.58
R7447 vss.n21850 vss.n21849 27.517
R7448 vss.n21733 vss.n21713 27.517
R7449 vss.n3799 vss.n3798 27.517
R7450 vss.n3682 vss.n3662 27.517
R7451 vss.n22597 vss.n22596 27.039
R7452 vss.n22578 vss.n22577 27.039
R7453 vss.n22389 vss.n22388 27.039
R7454 vss.n22370 vss.n22369 27.039
R7455 vss.n22181 vss.n22180 27.039
R7456 vss.n22162 vss.n22161 27.039
R7457 vss.n21525 vss.n21524 27.039
R7458 vss.n21506 vss.n21505 27.039
R7459 vss.n21317 vss.n21316 27.039
R7460 vss.n21298 vss.n21297 27.039
R7461 vss.n21109 vss.n21108 27.039
R7462 vss.n21090 vss.n21089 27.039
R7463 vss.n20901 vss.n20900 27.039
R7464 vss.n8760 vss.n8759 27.039
R7465 vss.n8741 vss.n8740 27.039
R7466 vss.n8552 vss.n8551 27.039
R7467 vss.n8533 vss.n8532 27.039
R7468 vss.n8344 vss.n8343 27.039
R7469 vss.n8325 vss.n8324 27.039
R7470 vss.n8136 vss.n8135 27.039
R7471 vss.n8117 vss.n8116 27.039
R7472 vss.n7928 vss.n7927 27.039
R7473 vss.n7909 vss.n7908 27.039
R7474 vss.n7719 vss.n7718 27.039
R7475 vss.n7700 vss.n7699 27.039
R7476 vss.n7511 vss.n7510 27.039
R7477 vss.n13889 vss.n13888 26.666
R7478 vss.n14435 vss.n14434 26.666
R7479 vss.n11105 vss.n11104 26.666
R7480 vss.n11895 vss.n11894 26.666
R7481 vss.n11962 vss.n11961 26.666
R7482 vss.n11888 vss.n11887 26.666
R7483 vss.n10774 vss.n10773 26.666
R7484 vss.n12625 vss.n12624 26.666
R7485 vss.n10615 vss.n10614 26.666
R7486 vss.n14760 vss.n14759 26.666
R7487 vss.n14933 vss.n14932 26.666
R7488 vss.n13402 vss.n13401 26.666
R7489 vss.n14127 vss.n14126 26.666
R7490 vss.n13474 vss.n13473 26.666
R7491 vss.n11412 vss.n11411 26.666
R7492 vss.n13803 vss.n13802 26.666
R7493 vss.n11420 vss.n11419 26.666
R7494 vss.n11600 vss.n11599 26.666
R7495 vss.n9815 vss.n9812 26.352
R7496 vss.n20478 vss.n20477 26.344
R7497 vss.n20599 vss.n20598 26.344
R7498 vss.n20707 vss.n20706 26.344
R7499 vss.n20822 vss.n20821 26.344
R7500 vss.n7088 vss.n7087 26.344
R7501 vss.n7209 vss.n7208 26.344
R7502 vss.n7317 vss.n7316 26.344
R7503 vss.n7432 vss.n7431 26.344
R7504 vss.n1701 vss.n1700 26.344
R7505 vss.n1820 vss.n1819 26.344
R7506 vss.n1931 vss.n1930 26.344
R7507 vss.n2060 vss.n2059 26.344
R7508 vss.n2175 vss.n2174 26.344
R7509 vss.n2305 vss.n2304 26.344
R7510 vss.n2420 vss.n2419 26.344
R7511 vss.n2549 vss.n2548 26.344
R7512 vss.n2664 vss.n2663 26.344
R7513 vss.n2793 vss.n2792 26.344
R7514 vss.n2902 vss.n2901 26.344
R7515 vss.n3032 vss.n3031 26.344
R7516 vss.n3147 vss.n3146 26.344
R7517 vss.n3276 vss.n3275 26.344
R7518 vss.n3388 vss.n3387 26.344
R7519 vss.n15161 vss.n15160 26.344
R7520 vss.n162 vss.n161 26.344
R7521 vss.n281 vss.n280 26.344
R7522 vss.n392 vss.n391 26.344
R7523 vss.n521 vss.n520 26.344
R7524 vss.n636 vss.n635 26.344
R7525 vss.n766 vss.n765 26.344
R7526 vss.n881 vss.n880 26.344
R7527 vss.n1010 vss.n1009 26.344
R7528 vss.n1125 vss.n1124 26.344
R7529 vss.n1254 vss.n1253 26.344
R7530 vss.n23349 vss.n23348 26.344
R7531 vss.n23220 vss.n23219 26.344
R7532 vss.n23105 vss.n23104 26.344
R7533 vss.n22976 vss.n22975 26.344
R7534 vss.n22865 vss.n22864 26.344
R7535 vss.n22795 vss.n22794 26.344
R7536 vss.n19028 vss.n17628 25.61
R7537 vss.n19000 vss.n17639 25.61
R7538 vss.n18897 vss.n17726 25.61
R7539 vss.n17748 vss.n17745 25.61
R7540 vss.n17837 vss.n17828 25.61
R7541 vss.n18759 vss.n17847 25.61
R7542 vss.n18656 vss.n17939 25.61
R7543 vss.n17961 vss.n17958 25.61
R7544 vss.n18050 vss.n18041 25.61
R7545 vss.n18518 vss.n18060 25.61
R7546 vss.n18415 vss.n18152 25.61
R7547 vss.n18174 vss.n18171 25.61
R7548 vss.n18263 vss.n18254 25.61
R7549 vss.n18275 vss.n17625 25.61
R7550 vss.n20293 vss.n17617 25.61
R7551 vss.n20273 vss.n19041 25.61
R7552 vss.n19137 vss.n19128 25.61
R7553 vss.n20146 vss.n19146 25.61
R7554 vss.n20043 vss.n19233 25.61
R7555 vss.n19255 vss.n19252 25.61
R7556 vss.n19344 vss.n19335 25.61
R7557 vss.n19899 vss.n19353 25.61
R7558 vss.n19796 vss.n19440 25.61
R7559 vss.n19462 vss.n19459 25.61
R7560 vss.n19551 vss.n19542 25.61
R7561 vss.n19652 vss.n19560 25.61
R7562 vss.n20320 vss.n20319 25.61
R7563 vss.n5638 vss.n4238 25.61
R7564 vss.n5610 vss.n4249 25.61
R7565 vss.n5507 vss.n4336 25.61
R7566 vss.n4358 vss.n4355 25.61
R7567 vss.n4447 vss.n4438 25.61
R7568 vss.n5369 vss.n4457 25.61
R7569 vss.n5266 vss.n4549 25.61
R7570 vss.n4571 vss.n4568 25.61
R7571 vss.n4660 vss.n4651 25.61
R7572 vss.n5128 vss.n4670 25.61
R7573 vss.n5025 vss.n4762 25.61
R7574 vss.n4784 vss.n4781 25.61
R7575 vss.n4873 vss.n4864 25.61
R7576 vss.n4885 vss.n4235 25.61
R7577 vss.n6903 vss.n4227 25.61
R7578 vss.n6883 vss.n5651 25.61
R7579 vss.n5747 vss.n5738 25.61
R7580 vss.n6756 vss.n5756 25.61
R7581 vss.n6653 vss.n5843 25.61
R7582 vss.n5865 vss.n5862 25.61
R7583 vss.n5954 vss.n5945 25.61
R7584 vss.n6509 vss.n5963 25.61
R7585 vss.n6406 vss.n6050 25.61
R7586 vss.n6072 vss.n6069 25.61
R7587 vss.n6161 vss.n6152 25.61
R7588 vss.n6262 vss.n6170 25.61
R7589 vss.n6930 vss.n6929 25.61
R7590 vss.n16690 vss.n16689 25.61
R7591 vss.n16869 vss.n16868 25.61
R7592 vss.n16920 vss.n16919 25.61
R7593 vss.n17105 vss.n17104 25.61
R7594 vss.n17156 vss.n17155 25.61
R7595 vss.n17267 vss.n17266 25.61
R7596 vss.n15915 vss.n15914 25.61
R7597 vss.n15967 vss.n15966 25.61
R7598 vss.n16151 vss.n16150 25.61
R7599 vss.n16203 vss.n16202 25.61
R7600 vss.n16276 vss.n16275 25.61
R7601 vss.n15391 vss.n15390 25.61
R7602 vss.n15440 vss.n15439 25.61
R7603 vss.n15627 vss.n15626 25.61
R7604 vss.n15676 vss.n15675 25.61
R7605 vss.n15855 vss.n15854 25.61
R7606 vss.n16338 vss.n16337 25.61
R7607 vss.n16387 vss.n16386 25.61
R7608 vss.n16574 vss.n16573 25.61
R7609 vss.n16623 vss.n16622 25.61
R7610 vss.n20433 vss.n20430 25.6
R7611 vss.n20435 vss.n20433 25.6
R7612 vss.n20439 vss.n20435 25.6
R7613 vss.n20441 vss.n20439 25.6
R7614 vss.n20428 vss.n20427 25.6
R7615 vss.n20427 vss.n20426 25.6
R7616 vss.n20426 vss.n20425 25.6
R7617 vss.n20425 vss.n20424 25.6
R7618 vss.n20424 vss.n20423 25.6
R7619 vss.n20423 vss.n20422 25.6
R7620 vss.n20422 vss.n20421 25.6
R7621 vss.n20421 vss.n20420 25.6
R7622 vss.n20420 vss.n20419 25.6
R7623 vss.n20419 vss.n20418 25.6
R7624 vss.n20418 vss.n20417 25.6
R7625 vss.n20417 vss.n20416 25.6
R7626 vss.n20416 vss.n20415 25.6
R7627 vss.n20415 vss.n20414 25.6
R7628 vss.n20862 vss.n20861 25.6
R7629 vss.n20863 vss.n20862 25.6
R7630 vss.n20864 vss.n20863 25.6
R7631 vss.n20865 vss.n20864 25.6
R7632 vss.n20866 vss.n20865 25.6
R7633 vss.n20867 vss.n20866 25.6
R7634 vss.n20868 vss.n20867 25.6
R7635 vss.n20869 vss.n20868 25.6
R7636 vss.n20870 vss.n20869 25.6
R7637 vss.n20871 vss.n20870 25.6
R7638 vss.n20872 vss.n20871 25.6
R7639 vss.n20873 vss.n20872 25.6
R7640 vss.n20874 vss.n20873 25.6
R7641 vss.n20875 vss.n20874 25.6
R7642 vss.n20876 vss.n20875 25.6
R7643 vss.n20881 vss.n20879 25.6
R7644 vss.n20884 vss.n20881 25.6
R7645 vss.n20886 vss.n20884 25.6
R7646 vss.n20890 vss.n20886 25.6
R7647 vss.n9635 vss.n9632 25.6
R7648 vss.n9632 vss.n9629 25.6
R7649 vss.n9629 vss.n9626 25.6
R7650 vss.n9626 vss.n9623 25.6
R7651 vss.n9623 vss.n9620 25.6
R7652 vss.n9620 vss.n9617 25.6
R7653 vss.n9617 vss.n9614 25.6
R7654 vss.n9614 vss.n9611 25.6
R7655 vss.n9611 vss.n9608 25.6
R7656 vss.n9608 vss.n9605 25.6
R7657 vss.n9605 vss.n9602 25.6
R7658 vss.n9602 vss.n9599 25.6
R7659 vss.n9599 vss.n9596 25.6
R7660 vss.n9596 vss.n9593 25.6
R7661 vss.n9593 vss.n9590 25.6
R7662 vss.n9590 vss.n9587 25.6
R7663 vss.n9587 vss.n9584 25.6
R7664 vss.n9584 vss.n9581 25.6
R7665 vss.n9581 vss.n9578 25.6
R7666 vss.n9578 vss.n9575 25.6
R7667 vss.n9575 vss.n9572 25.6
R7668 vss.n9572 vss.n9569 25.6
R7669 vss.n9569 vss.n9566 25.6
R7670 vss.n9566 vss.n9563 25.6
R7671 vss.n9563 vss.n9560 25.6
R7672 vss.n9560 vss.n9557 25.6
R7673 vss.n9557 vss.n9554 25.6
R7674 vss.n9554 vss.n9551 25.6
R7675 vss.n9551 vss.n9548 25.6
R7676 vss.n9548 vss.n9545 25.6
R7677 vss.n9545 vss.n9542 25.6
R7678 vss.n9542 vss.n9539 25.6
R7679 vss.n9539 vss.n9536 25.6
R7680 vss.n9536 vss.n9533 25.6
R7681 vss.n9533 vss.n9530 25.6
R7682 vss.n9530 vss.n9527 25.6
R7683 vss.n9527 vss.n9524 25.6
R7684 vss.n9524 vss.n9521 25.6
R7685 vss.n9521 vss.n9518 25.6
R7686 vss.n9518 vss.n9515 25.6
R7687 vss.n9515 vss.n9512 25.6
R7688 vss.n9512 vss.n9509 25.6
R7689 vss.n9509 vss.n9506 25.6
R7690 vss.n9506 vss.n9503 25.6
R7691 vss.n9503 vss.n9500 25.6
R7692 vss.n9500 vss.n9497 25.6
R7693 vss.n9497 vss.n9494 25.6
R7694 vss.n9494 vss.n9491 25.6
R7695 vss.n9491 vss.n9488 25.6
R7696 vss.n9488 vss.n9485 25.6
R7697 vss.n9485 vss.n9482 25.6
R7698 vss.n9482 vss.n9479 25.6
R7699 vss.n9479 vss.n9476 25.6
R7700 vss.n9476 vss.n9473 25.6
R7701 vss.n9473 vss.n9470 25.6
R7702 vss.n9470 vss.n9467 25.6
R7703 vss.n9467 vss.n9464 25.6
R7704 vss.n9464 vss.n9461 25.6
R7705 vss.n9461 vss.n9458 25.6
R7706 vss.n9458 vss.n9455 25.6
R7707 vss.n9455 vss.n9452 25.6
R7708 vss.n9452 vss.n9449 25.6
R7709 vss.n9449 vss.n9446 25.6
R7710 vss.n9446 vss.n9443 25.6
R7711 vss.n9443 vss.n9440 25.6
R7712 vss.n9440 vss.n9437 25.6
R7713 vss.n9437 vss.n9434 25.6
R7714 vss.n9434 vss.n9431 25.6
R7715 vss.n9431 vss.n9428 25.6
R7716 vss.n9428 vss.n9425 25.6
R7717 vss.n9425 vss.n9422 25.6
R7718 vss.n9422 vss.n9419 25.6
R7719 vss.n9419 vss.n9416 25.6
R7720 vss.n9416 vss.n9413 25.6
R7721 vss.n9413 vss.n9410 25.6
R7722 vss.n9410 vss.n9407 25.6
R7723 vss.n9407 vss.n9404 25.6
R7724 vss.n9404 vss.n9401 25.6
R7725 vss.n9401 vss.n9398 25.6
R7726 vss.n9398 vss.n9395 25.6
R7727 vss.n9395 vss.n9392 25.6
R7728 vss.n9392 vss.n9389 25.6
R7729 vss.n9389 vss.n9386 25.6
R7730 vss.n9386 vss.n9383 25.6
R7731 vss.n9383 vss.n9380 25.6
R7732 vss.n9380 vss.n9377 25.6
R7733 vss.n9377 vss.n9374 25.6
R7734 vss.n9374 vss.n9371 25.6
R7735 vss.n9371 vss.n9368 25.6
R7736 vss.n9368 vss.n9365 25.6
R7737 vss.n9365 vss.n9362 25.6
R7738 vss.n9362 vss.n9359 25.6
R7739 vss.n9359 vss.n9356 25.6
R7740 vss.n9356 vss.n9353 25.6
R7741 vss.n9353 vss.n9350 25.6
R7742 vss.n9350 vss.n9347 25.6
R7743 vss.n9347 vss.n9344 25.6
R7744 vss.n9344 vss.n9341 25.6
R7745 vss.n9341 vss.n9338 25.6
R7746 vss.n9338 vss.n9335 25.6
R7747 vss.n9335 vss.n9332 25.6
R7748 vss.n9332 vss.n9329 25.6
R7749 vss.n9329 vss.n9326 25.6
R7750 vss.n9326 vss.n9323 25.6
R7751 vss.n9323 vss.n9320 25.6
R7752 vss.n9320 vss.n9317 25.6
R7753 vss.n9317 vss.n9314 25.6
R7754 vss.n9314 vss.n9311 25.6
R7755 vss.n9311 vss.n9308 25.6
R7756 vss.n9308 vss.n9305 25.6
R7757 vss.n9305 vss.n9302 25.6
R7758 vss.n9302 vss.n9299 25.6
R7759 vss.n9299 vss.n9296 25.6
R7760 vss.n9296 vss.n9293 25.6
R7761 vss.n9293 vss.n9290 25.6
R7762 vss.n9290 vss.n9287 25.6
R7763 vss.n9287 vss.n9284 25.6
R7764 vss.n9284 vss.n9281 25.6
R7765 vss.n9281 vss.n9278 25.6
R7766 vss.n9278 vss.n9275 25.6
R7767 vss.n9275 vss.n9272 25.6
R7768 vss.n9269 vss.n9266 25.6
R7769 vss.n9266 vss.n9263 25.6
R7770 vss.n9263 vss.n9260 25.6
R7771 vss.n9260 vss.n9257 25.6
R7772 vss.n9257 vss.n9254 25.6
R7773 vss.n9254 vss.n9251 25.6
R7774 vss.n9251 vss.n9248 25.6
R7775 vss.n9248 vss.n9245 25.6
R7776 vss.n9245 vss.n9242 25.6
R7777 vss.n9242 vss.n9239 25.6
R7778 vss.n9238 vss.n9235 25.6
R7779 vss.n9235 vss.n9232 25.6
R7780 vss.n9232 vss.n9229 25.6
R7781 vss.n9229 vss.n9226 25.6
R7782 vss.n9226 vss.n9223 25.6
R7783 vss.n9223 vss.n9220 25.6
R7784 vss.n9220 vss.n9217 25.6
R7785 vss.n9217 vss.n9214 25.6
R7786 vss.n9214 vss.n9211 25.6
R7787 vss.n9211 vss.n9208 25.6
R7788 vss.n9752 vss.n9749 25.6
R7789 vss.n9755 vss.n9752 25.6
R7790 vss.n9758 vss.n9755 25.6
R7791 vss.n9761 vss.n9758 25.6
R7792 vss.n9764 vss.n9761 25.6
R7793 vss.n9767 vss.n9764 25.6
R7794 vss.n9770 vss.n9767 25.6
R7795 vss.n9773 vss.n9770 25.6
R7796 vss.n9776 vss.n9773 25.6
R7797 vss.n9779 vss.n9776 25.6
R7798 vss.n10178 vss.n10175 25.6
R7799 vss.n10175 vss.n10172 25.6
R7800 vss.n10172 vss.n10169 25.6
R7801 vss.n10169 vss.n10166 25.6
R7802 vss.n10166 vss.n10163 25.6
R7803 vss.n10163 vss.n10160 25.6
R7804 vss.n10160 vss.n10157 25.6
R7805 vss.n10157 vss.n10154 25.6
R7806 vss.n10154 vss.n10151 25.6
R7807 vss.n10151 vss.n10148 25.6
R7808 vss.n10148 vss.n10145 25.6
R7809 vss.n10145 vss.n10142 25.6
R7810 vss.n10142 vss.n10139 25.6
R7811 vss.n10139 vss.n10136 25.6
R7812 vss.n10136 vss.n10133 25.6
R7813 vss.n10133 vss.n10130 25.6
R7814 vss.n10130 vss.n10127 25.6
R7815 vss.n10127 vss.n10124 25.6
R7816 vss.n10124 vss.n10121 25.6
R7817 vss.n10121 vss.n10118 25.6
R7818 vss.n10118 vss.n10115 25.6
R7819 vss.n10115 vss.n10112 25.6
R7820 vss.n10112 vss.n10109 25.6
R7821 vss.n10109 vss.n10106 25.6
R7822 vss.n10106 vss.n10103 25.6
R7823 vss.n10103 vss.n10100 25.6
R7824 vss.n10100 vss.n10097 25.6
R7825 vss.n10097 vss.n10094 25.6
R7826 vss.n10094 vss.n10091 25.6
R7827 vss.n10091 vss.n10088 25.6
R7828 vss.n10088 vss.n10085 25.6
R7829 vss.n10085 vss.n10082 25.6
R7830 vss.n10082 vss.n10079 25.6
R7831 vss.n10079 vss.n10076 25.6
R7832 vss.n10076 vss.n10073 25.6
R7833 vss.n10073 vss.n10070 25.6
R7834 vss.n10070 vss.n10067 25.6
R7835 vss.n10067 vss.n10064 25.6
R7836 vss.n10064 vss.n10061 25.6
R7837 vss.n10061 vss.n10058 25.6
R7838 vss.n10058 vss.n10055 25.6
R7839 vss.n10055 vss.n10052 25.6
R7840 vss.n10052 vss.n10049 25.6
R7841 vss.n10049 vss.n10046 25.6
R7842 vss.n10046 vss.n10043 25.6
R7843 vss.n10043 vss.n10040 25.6
R7844 vss.n10040 vss.n10037 25.6
R7845 vss.n10037 vss.n10034 25.6
R7846 vss.n10034 vss.n10031 25.6
R7847 vss.n10031 vss.n10028 25.6
R7848 vss.n10028 vss.n10025 25.6
R7849 vss.n10025 vss.n10022 25.6
R7850 vss.n10022 vss.n10019 25.6
R7851 vss.n10019 vss.n10016 25.6
R7852 vss.n10016 vss.n10013 25.6
R7853 vss.n10013 vss.n10010 25.6
R7854 vss.n10010 vss.n10007 25.6
R7855 vss.n10007 vss.n10004 25.6
R7856 vss.n10004 vss.n10001 25.6
R7857 vss.n10001 vss.n9998 25.6
R7858 vss.n9998 vss.n9995 25.6
R7859 vss.n9995 vss.n9992 25.6
R7860 vss.n9992 vss.n9989 25.6
R7861 vss.n9989 vss.n9986 25.6
R7862 vss.n9986 vss.n9983 25.6
R7863 vss.n9983 vss.n9980 25.6
R7864 vss.n9980 vss.n9977 25.6
R7865 vss.n9977 vss.n9974 25.6
R7866 vss.n9974 vss.n9971 25.6
R7867 vss.n9971 vss.n9968 25.6
R7868 vss.n9968 vss.n9965 25.6
R7869 vss.n9965 vss.n9962 25.6
R7870 vss.n9962 vss.n9959 25.6
R7871 vss.n9959 vss.n9956 25.6
R7872 vss.n9956 vss.n9953 25.6
R7873 vss.n9953 vss.n9950 25.6
R7874 vss.n9950 vss.n9947 25.6
R7875 vss.n9947 vss.n9944 25.6
R7876 vss.n9944 vss.n9941 25.6
R7877 vss.n9941 vss.n9938 25.6
R7878 vss.n9938 vss.n9935 25.6
R7879 vss.n9935 vss.n9932 25.6
R7880 vss.n9932 vss.n9929 25.6
R7881 vss.n9929 vss.n9926 25.6
R7882 vss.n9926 vss.n9923 25.6
R7883 vss.n9923 vss.n9920 25.6
R7884 vss.n9920 vss.n9917 25.6
R7885 vss.n9917 vss.n9914 25.6
R7886 vss.n9914 vss.n9911 25.6
R7887 vss.n9911 vss.n9908 25.6
R7888 vss.n9908 vss.n9905 25.6
R7889 vss.n9905 vss.n9902 25.6
R7890 vss.n9902 vss.n9899 25.6
R7891 vss.n9899 vss.n9896 25.6
R7892 vss.n9896 vss.n9893 25.6
R7893 vss.n9893 vss.n9890 25.6
R7894 vss.n9890 vss.n9887 25.6
R7895 vss.n9887 vss.n9884 25.6
R7896 vss.n9884 vss.n9881 25.6
R7897 vss.n9881 vss.n9878 25.6
R7898 vss.n9878 vss.n9875 25.6
R7899 vss.n9875 vss.n9872 25.6
R7900 vss.n9872 vss.n9869 25.6
R7901 vss.n9869 vss.n9866 25.6
R7902 vss.n9866 vss.n9863 25.6
R7903 vss.n9863 vss.n9860 25.6
R7904 vss.n9860 vss.n9857 25.6
R7905 vss.n9857 vss.n9854 25.6
R7906 vss.n9854 vss.n9851 25.6
R7907 vss.n9851 vss.n9848 25.6
R7908 vss.n9848 vss.n9845 25.6
R7909 vss.n9845 vss.n9842 25.6
R7910 vss.n9842 vss.n9839 25.6
R7911 vss.n9839 vss.n9836 25.6
R7912 vss.n9836 vss.n9833 25.6
R7913 vss.n9833 vss.n9830 25.6
R7914 vss.n9830 vss.n9827 25.6
R7915 vss.n9827 vss.n9824 25.6
R7916 vss.n9824 vss.n9821 25.6
R7917 vss.n9821 vss.n9818 25.6
R7918 vss.n9818 vss.n9815 25.6
R7919 vss.n9812 vss.n9809 25.6
R7920 vss.n9809 vss.n9806 25.6
R7921 vss.n9806 vss.n9803 25.6
R7922 vss.n9803 vss.n9800 25.6
R7923 vss.n9800 vss.n9797 25.6
R7924 vss.n9797 vss.n9794 25.6
R7925 vss.n9794 vss.n9791 25.6
R7926 vss.n9791 vss.n9788 25.6
R7927 vss.n9788 vss.n9785 25.6
R7928 vss.n9785 vss.n9782 25.6
R7929 vss.n7043 vss.n7040 25.6
R7930 vss.n7045 vss.n7043 25.6
R7931 vss.n7049 vss.n7045 25.6
R7932 vss.n7051 vss.n7049 25.6
R7933 vss.n7038 vss.n7037 25.6
R7934 vss.n7037 vss.n7036 25.6
R7935 vss.n7036 vss.n7035 25.6
R7936 vss.n7035 vss.n7034 25.6
R7937 vss.n7034 vss.n7033 25.6
R7938 vss.n7033 vss.n7032 25.6
R7939 vss.n7032 vss.n7031 25.6
R7940 vss.n7031 vss.n7030 25.6
R7941 vss.n7030 vss.n7029 25.6
R7942 vss.n7029 vss.n7028 25.6
R7943 vss.n7028 vss.n7027 25.6
R7944 vss.n7027 vss.n7026 25.6
R7945 vss.n7026 vss.n7025 25.6
R7946 vss.n7025 vss.n7024 25.6
R7947 vss.n7472 vss.n7471 25.6
R7948 vss.n7473 vss.n7472 25.6
R7949 vss.n7474 vss.n7473 25.6
R7950 vss.n7475 vss.n7474 25.6
R7951 vss.n7476 vss.n7475 25.6
R7952 vss.n7477 vss.n7476 25.6
R7953 vss.n7478 vss.n7477 25.6
R7954 vss.n7479 vss.n7478 25.6
R7955 vss.n7480 vss.n7479 25.6
R7956 vss.n7481 vss.n7480 25.6
R7957 vss.n7482 vss.n7481 25.6
R7958 vss.n7483 vss.n7482 25.6
R7959 vss.n7484 vss.n7483 25.6
R7960 vss.n7485 vss.n7484 25.6
R7961 vss.n7486 vss.n7485 25.6
R7962 vss.n7491 vss.n7489 25.6
R7963 vss.n7494 vss.n7491 25.6
R7964 vss.n7496 vss.n7494 25.6
R7965 vss.n7500 vss.n7496 25.6
R7966 vss.n1673 vss.n1670 25.6
R7967 vss.n1675 vss.n1673 25.6
R7968 vss.n1679 vss.n1675 25.6
R7969 vss.n1681 vss.n1679 25.6
R7970 vss.n1668 vss.n1667 25.6
R7971 vss.n1667 vss.n1666 25.6
R7972 vss.n1666 vss.n1665 25.6
R7973 vss.n1665 vss.n1664 25.6
R7974 vss.n1664 vss.n1663 25.6
R7975 vss.n1663 vss.n1662 25.6
R7976 vss.n1662 vss.n1661 25.6
R7977 vss.n1661 vss.n1660 25.6
R7978 vss.n1660 vss.n1659 25.6
R7979 vss.n1659 vss.n1658 25.6
R7980 vss.n1658 vss.n1657 25.6
R7981 vss.n1657 vss.n1656 25.6
R7982 vss.n1656 vss.n1655 25.6
R7983 vss.n1984 vss.n1983 25.6
R7984 vss.n2014 vss.n2013 25.6
R7985 vss.n2229 vss.n2228 25.6
R7986 vss.n2258 vss.n2257 25.6
R7987 vss.n2473 vss.n2472 25.6
R7988 vss.n2502 vss.n2501 25.6
R7989 vss.n2718 vss.n2717 25.6
R7990 vss.n2747 vss.n2746 25.6
R7991 vss.n1535 vss.n1534 25.6
R7992 vss.n1536 vss.n1535 25.6
R7993 vss.n1537 vss.n1536 25.6
R7994 vss.n2956 vss.n2955 25.6
R7995 vss.n2985 vss.n2984 25.6
R7996 vss.n3200 vss.n3199 25.6
R7997 vss.n3230 vss.n3229 25.6
R7998 vss.n15127 vss.n15126 25.6
R7999 vss.n15128 vss.n15127 25.6
R8000 vss.n15129 vss.n15128 25.6
R8001 vss.n15130 vss.n15129 25.6
R8002 vss.n15131 vss.n15130 25.6
R8003 vss.n15132 vss.n15131 25.6
R8004 vss.n15133 vss.n15132 25.6
R8005 vss.n15134 vss.n15133 25.6
R8006 vss.n15135 vss.n15134 25.6
R8007 vss.n15136 vss.n15135 25.6
R8008 vss.n15137 vss.n15136 25.6
R8009 vss.n15138 vss.n15137 25.6
R8010 vss.n15139 vss.n15138 25.6
R8011 vss.n15144 vss.n15142 25.6
R8012 vss.n15147 vss.n15144 25.6
R8013 vss.n15149 vss.n15147 25.6
R8014 vss.n15153 vss.n15149 25.6
R8015 vss.n134 vss.n131 25.6
R8016 vss.n136 vss.n134 25.6
R8017 vss.n140 vss.n136 25.6
R8018 vss.n142 vss.n140 25.6
R8019 vss.n129 vss.n128 25.6
R8020 vss.n128 vss.n127 25.6
R8021 vss.n127 vss.n126 25.6
R8022 vss.n126 vss.n125 25.6
R8023 vss.n125 vss.n124 25.6
R8024 vss.n124 vss.n123 25.6
R8025 vss.n123 vss.n122 25.6
R8026 vss.n122 vss.n121 25.6
R8027 vss.n121 vss.n120 25.6
R8028 vss.n120 vss.n119 25.6
R8029 vss.n119 vss.n118 25.6
R8030 vss.n118 vss.n117 25.6
R8031 vss.n117 vss.n116 25.6
R8032 vss.n445 vss.n444 25.6
R8033 vss.n475 vss.n474 25.6
R8034 vss.n690 vss.n689 25.6
R8035 vss.n719 vss.n718 25.6
R8036 vss.n934 vss.n933 25.6
R8037 vss.n963 vss.n962 25.6
R8038 vss.n1179 vss.n1178 25.6
R8039 vss.n1208 vss.n1207 25.6
R8040 vss.n23302 vss.n23301 25.6
R8041 vss.n23275 vss.n23274 25.6
R8042 vss.n23058 vss.n23057 25.6
R8043 vss.n23030 vss.n23029 25.6
R8044 vss.n22761 vss.n22760 25.6
R8045 vss.n22762 vss.n22761 25.6
R8046 vss.n22763 vss.n22762 25.6
R8047 vss.n22764 vss.n22763 25.6
R8048 vss.n22765 vss.n22764 25.6
R8049 vss.n22766 vss.n22765 25.6
R8050 vss.n22767 vss.n22766 25.6
R8051 vss.n22768 vss.n22767 25.6
R8052 vss.n22769 vss.n22768 25.6
R8053 vss.n22770 vss.n22769 25.6
R8054 vss.n22771 vss.n22770 25.6
R8055 vss.n22772 vss.n22771 25.6
R8056 vss.n22773 vss.n22772 25.6
R8057 vss.n22778 vss.n22776 25.6
R8058 vss.n22781 vss.n22778 25.6
R8059 vss.n22783 vss.n22781 25.6
R8060 vss.n22787 vss.n22783 25.6
R8061 vss.n12423 vss.n12422 25.356
R8062 vss.n12596 vss.n12595 25.356
R8063 vss.n14489 vss.n14488 25.356
R8064 vss.n14396 vss.n14395 25.356
R8065 vss.n14659 vss.n14658 25.356
R8066 vss.n13578 vss.n13577 25.356
R8067 vss.n15013 vss.n15012 25.356
R8068 vss.n10504 vss.n10503 25.356
R8069 vss.n13296 vss.n13295 25.356
R8070 vss.n13337 vss.n13336 25.356
R8071 vss.n13238 vss.n13237 25.356
R8072 vss.n14959 vss.n14958 25.356
R8073 vss.n14355 vss.n14354 25.356
R8074 vss.n13861 vss.n13860 25.356
R8075 vss.n13976 vss.n13975 25.356
R8076 vss.n11571 vss.n11570 25.356
R8077 vss.n11758 vss.n11757 25.356
R8078 vss.n11048 vss.n11047 25.356
R8079 vss.n10822 vss.n10821 25.356
R8080 vss.n10896 vss.n10895 25.356
R8081 vss.n10949 vss.n10948 25.356
R8082 vss.n11009 vss.n11008 25.356
R8083 vss.n12581 vss.n12580 25.356
R8084 vss.n12077 vss.n12076 25.356
R8085 vss.n22720 vss.n22718 25.107
R8086 vss.n22671 vss.n22669 25.107
R8087 vss.n22512 vss.n22510 25.107
R8088 vss.n22463 vss.n22461 25.107
R8089 vss.n22304 vss.n22302 25.107
R8090 vss.n22255 vss.n22253 25.107
R8091 vss.n22096 vss.n22094 25.107
R8092 vss.n21587 vss.n21585 25.107
R8093 vss.n21440 vss.n21438 25.107
R8094 vss.n21391 vss.n21389 25.107
R8095 vss.n21232 vss.n21230 25.107
R8096 vss.n21183 vss.n21181 25.107
R8097 vss.n21024 vss.n21022 25.107
R8098 vss.n20975 vss.n20973 25.107
R8099 vss.n8883 vss.n8881 25.107
R8100 vss.n8834 vss.n8832 25.107
R8101 vss.n8675 vss.n8673 25.107
R8102 vss.n8626 vss.n8624 25.107
R8103 vss.n8467 vss.n8465 25.107
R8104 vss.n8418 vss.n8416 25.107
R8105 vss.n8259 vss.n8257 25.107
R8106 vss.n8210 vss.n8208 25.107
R8107 vss.n8051 vss.n8049 25.107
R8108 vss.n8002 vss.n8000 25.107
R8109 vss.n7842 vss.n7840 25.107
R8110 vss.n7793 vss.n7791 25.107
R8111 vss.n7634 vss.n7632 25.107
R8112 vss.n7585 vss.n7583 25.107
R8113 vss.n11772 vss.n11771 25
R8114 vss.n11349 vss.n11348 25
R8115 vss.n11357 vss.n11356 25
R8116 vss.n10746 vss.n10745 25
R8117 vss.n12434 vss.n12433 25
R8118 vss.n13216 vss.n13215 25
R8119 vss.n13327 vss.n13326 25
R8120 vss.n13570 vss.n13569 25
R8121 vss.n14651 vss.n14650 25
R8122 vss.n14034 vss.n14033 25
R8123 vss.n18969 vss.n17670 23.64
R8124 vss.n18932 vss.n17697 23.64
R8125 vss.n18849 vss.n17771 23.64
R8126 vss.n18807 vss.n17803 23.64
R8127 vss.n18724 vss.n17878 23.64
R8128 vss.n18691 vss.n17910 23.64
R8129 vss.n18608 vss.n17984 23.64
R8130 vss.n18566 vss.n18016 23.64
R8131 vss.n18483 vss.n18091 23.64
R8132 vss.n18450 vss.n18123 23.64
R8133 vss.n18367 vss.n18197 23.64
R8134 vss.n18325 vss.n18229 23.64
R8135 vss.n20242 vss.n19071 23.64
R8136 vss.n20200 vss.n19103 23.64
R8137 vss.n20115 vss.n19177 23.64
R8138 vss.n20078 vss.n19204 23.64
R8139 vss.n19995 vss.n19278 23.64
R8140 vss.n19953 vss.n19310 23.64
R8141 vss.n19868 vss.n19384 23.64
R8142 vss.n19831 vss.n19411 23.64
R8143 vss.n19748 vss.n19485 23.64
R8144 vss.n19706 vss.n19517 23.64
R8145 vss.n19602 vss.n19599 23.64
R8146 vss.n20343 vss.n17598 23.64
R8147 vss.n5579 vss.n4280 23.64
R8148 vss.n5542 vss.n4307 23.64
R8149 vss.n5459 vss.n4381 23.64
R8150 vss.n5417 vss.n4413 23.64
R8151 vss.n5334 vss.n4488 23.64
R8152 vss.n5301 vss.n4520 23.64
R8153 vss.n5218 vss.n4594 23.64
R8154 vss.n5176 vss.n4626 23.64
R8155 vss.n5093 vss.n4701 23.64
R8156 vss.n5060 vss.n4733 23.64
R8157 vss.n4977 vss.n4807 23.64
R8158 vss.n4935 vss.n4839 23.64
R8159 vss.n6852 vss.n5681 23.64
R8160 vss.n6810 vss.n5713 23.64
R8161 vss.n6725 vss.n5787 23.64
R8162 vss.n6688 vss.n5814 23.64
R8163 vss.n6605 vss.n5888 23.64
R8164 vss.n6563 vss.n5920 23.64
R8165 vss.n6478 vss.n5994 23.64
R8166 vss.n6441 vss.n6021 23.64
R8167 vss.n6358 vss.n6095 23.64
R8168 vss.n6316 vss.n6127 23.64
R8169 vss.n6212 vss.n6209 23.64
R8170 vss.n6953 vss.n4208 23.64
R8171 vss.n16750 vss.n16746 23.64
R8172 vss.n16819 vss.n16815 23.64
R8173 vss.n16980 vss.n16976 23.64
R8174 vss.n17053 vss.n17049 23.64
R8175 vss.n17216 vss.n17212 23.64
R8176 vss.n17304 vss.n17300 23.64
R8177 vss.n16027 vss.n16025 23.64
R8178 vss.n16099 vss.n16097 23.64
R8179 vss.n15299 vss.n15295 23.64
R8180 vss.n15338 vss.n15334 23.64
R8181 vss.n15500 vss.n15496 23.64
R8182 vss.n15575 vss.n15571 23.64
R8183 vss.n15736 vss.n15732 23.64
R8184 vss.n15803 vss.n15799 23.64
R8185 vss.n16447 vss.n16443 23.64
R8186 vss.n16522 vss.n16518 23.64
R8187 vss.n14285 vss.n14284 23.634
R8188 vss.n13602 vss.n13601 23.634
R8189 vss.n12284 vss.n12283 23.634
R8190 vss.n12784 vss.n12780 23.634
R8191 vss.n13207 vss.n13202 23.634
R8192 vss.n13060 vss.n13056 23.634
R8193 vss.n13771 vss.n13770 23.592
R8194 vss.n12098 vss.n12097 23.592
R8195 vss.n13521 vss.n13520 23.592
R8196 vss.n13809 vss.n13808 23.544
R8197 vss.n10914 vss.n10913 23.333
R8198 vss.n10834 vss.n10833 23.333
R8199 vss.n10596 vss.n10595 23.333
R8200 vss.n10494 vss.n10493 23.333
R8201 vss.n10587 vss.n10586 23.333
R8202 vss.n11401 vss.n11400 23.333
R8203 vss.n20412 vss.n20411 23.316
R8204 vss.n7022 vss.n7021 23.316
R8205 vss.n20457 vss.n17546 23.222
R8206 vss.n20845 vss.t165 23.222
R8207 vss.n7067 vss.n4156 23.222
R8208 vss.n7455 vss.t210 23.222
R8209 vss.n15175 vss.t90 23.185
R8210 vss.n22809 vss.t99 23.185
R8211 vss.n22611 vss.n22610 23.176
R8212 vss.n22564 vss.n22563 23.176
R8213 vss.n22403 vss.n22402 23.176
R8214 vss.n22356 vss.n22355 23.176
R8215 vss.n22195 vss.n22194 23.176
R8216 vss.n22148 vss.n22147 23.176
R8217 vss.n21539 vss.n21538 23.176
R8218 vss.n21492 vss.n21491 23.176
R8219 vss.n21331 vss.n21330 23.176
R8220 vss.n21284 vss.n21283 23.176
R8221 vss.n21123 vss.n21122 23.176
R8222 vss.n21076 vss.n21075 23.176
R8223 vss.n20915 vss.n20914 23.176
R8224 vss.n12142 vss.n12140 23.176
R8225 vss.n11974 vss.n11972 23.176
R8226 vss.n11920 vss.n11918 23.176
R8227 vss.n14336 vss.n14334 23.176
R8228 vss.n11624 vss.n11622 23.176
R8229 vss.n11673 vss.n11671 23.176
R8230 vss.n14814 vss.n14812 23.176
R8231 vss.n14613 vss.n14611 23.176
R8232 vss.n14553 vss.n14551 23.176
R8233 vss.n14904 vss.n14902 23.176
R8234 vss.n15052 vss.n15050 23.176
R8235 vss.n10546 vss.n10544 23.176
R8236 vss.n8774 vss.n8773 23.176
R8237 vss.n8727 vss.n8726 23.176
R8238 vss.n8566 vss.n8565 23.176
R8239 vss.n8519 vss.n8518 23.176
R8240 vss.n8358 vss.n8357 23.176
R8241 vss.n8311 vss.n8310 23.176
R8242 vss.n8150 vss.n8149 23.176
R8243 vss.n8103 vss.n8102 23.176
R8244 vss.n7942 vss.n7941 23.176
R8245 vss.n7895 vss.n7894 23.176
R8246 vss.n7733 vss.n7732 23.176
R8247 vss.n7686 vss.n7685 23.176
R8248 vss.n7525 vss.n7524 23.176
R8249 vss.n20468 vss.n20463 23.051
R8250 vss.n20619 vss.n20614 23.051
R8251 vss.n20697 vss.n20692 23.051
R8252 vss.n20842 vss.n20837 23.051
R8253 vss.n7078 vss.n7073 23.051
R8254 vss.n7229 vss.n7224 23.051
R8255 vss.n7307 vss.n7302 23.051
R8256 vss.n7452 vss.n7447 23.051
R8257 vss.n1691 vss.n1686 23.051
R8258 vss.n1840 vss.n1835 23.051
R8259 vss.n1921 vss.n1915 23.051
R8260 vss.n2082 vss.n2076 23.051
R8261 vss.n2165 vss.n2159 23.051
R8262 vss.n2327 vss.n2321 23.051
R8263 vss.n2410 vss.n2404 23.051
R8264 vss.n2571 vss.n2565 23.051
R8265 vss.n2654 vss.n2648 23.051
R8266 vss.n2814 vss.n2809 23.051
R8267 vss.n2892 vss.n2886 23.051
R8268 vss.n3054 vss.n3048 23.051
R8269 vss.n3137 vss.n3131 23.051
R8270 vss.n3298 vss.n3292 23.051
R8271 vss.n3378 vss.n3373 23.051
R8272 vss.n3487 vss.n3482 23.051
R8273 vss.n152 vss.n147 23.051
R8274 vss.n301 vss.n296 23.051
R8275 vss.n382 vss.n376 23.051
R8276 vss.n543 vss.n537 23.051
R8277 vss.n626 vss.n620 23.051
R8278 vss.n788 vss.n782 23.051
R8279 vss.n871 vss.n865 23.051
R8280 vss.n1032 vss.n1026 23.051
R8281 vss.n1115 vss.n1109 23.051
R8282 vss.n1276 vss.n1270 23.051
R8283 vss.n23371 vss.n23365 23.051
R8284 vss.n23210 vss.n23204 23.051
R8285 vss.n23127 vss.n23121 23.051
R8286 vss.n22966 vss.n22960 23.051
R8287 vss.n22885 vss.n22880 23.051
R8288 vss.n1462 vss.n1457 23.051
R8289 vss.n1695 vss.n1654 23.007
R8290 vss.n156 vss.n115 23.007
R8291 vss.n21788 vss.n21690 22.141
R8292 vss.n3737 vss.n3639 22.141
R8293 vss.n21790 vss.n21689 21.97
R8294 vss.n3739 vss.n3638 21.97
R8295 vss.n18996 vss.n17645 21.67
R8296 vss.n18905 vss.n17719 21.67
R8297 vss.n18872 vss.n17746 21.67
R8298 vss.n18784 vss.n17826 21.67
R8299 vss.n18751 vss.n17859 21.67
R8300 vss.n18664 vss.n17932 21.67
R8301 vss.n18631 vss.n17959 21.67
R8302 vss.n18543 vss.n18039 21.67
R8303 vss.n18510 vss.n18072 21.67
R8304 vss.n18423 vss.n18145 21.67
R8305 vss.n18390 vss.n18172 21.67
R8306 vss.n18302 vss.n18252 21.67
R8307 vss.n20265 vss.n19049 21.67
R8308 vss.n20177 vss.n19126 21.67
R8309 vss.n20142 vss.n19152 21.67
R8310 vss.n20051 vss.n19226 21.67
R8311 vss.n20018 vss.n19253 21.67
R8312 vss.n19930 vss.n19333 21.67
R8313 vss.n19895 vss.n19359 21.67
R8314 vss.n19804 vss.n19433 21.67
R8315 vss.n19771 vss.n19460 21.67
R8316 vss.n19683 vss.n19540 21.67
R8317 vss.n19648 vss.n19566 21.67
R8318 vss.n20325 vss.n20324 21.67
R8319 vss.n5606 vss.n4255 21.67
R8320 vss.n5515 vss.n4329 21.67
R8321 vss.n5482 vss.n4356 21.67
R8322 vss.n5394 vss.n4436 21.67
R8323 vss.n5361 vss.n4469 21.67
R8324 vss.n5274 vss.n4542 21.67
R8325 vss.n5241 vss.n4569 21.67
R8326 vss.n5153 vss.n4649 21.67
R8327 vss.n5120 vss.n4682 21.67
R8328 vss.n5033 vss.n4755 21.67
R8329 vss.n5000 vss.n4782 21.67
R8330 vss.n4912 vss.n4862 21.67
R8331 vss.n6875 vss.n5659 21.67
R8332 vss.n6787 vss.n5736 21.67
R8333 vss.n6752 vss.n5762 21.67
R8334 vss.n6661 vss.n5836 21.67
R8335 vss.n6628 vss.n5863 21.67
R8336 vss.n6540 vss.n5943 21.67
R8337 vss.n6505 vss.n5969 21.67
R8338 vss.n6414 vss.n6043 21.67
R8339 vss.n6381 vss.n6070 21.67
R8340 vss.n6293 vss.n6150 21.67
R8341 vss.n6258 vss.n6176 21.67
R8342 vss.n6935 vss.n6934 21.67
R8343 vss.n16704 vss.n16703 21.67
R8344 vss.n16855 vss.n16854 21.67
R8345 vss.n16934 vss.n16933 21.67
R8346 vss.n17091 vss.n17090 21.67
R8347 vss.n17170 vss.n17169 21.67
R8348 vss.n17308 vss.n17307 21.67
R8349 vss.n15901 vss.n15900 21.67
R8350 vss.n15981 vss.n15980 21.67
R8351 vss.n16137 vss.n16136 21.67
R8352 vss.n16217 vss.n16216 21.67
R8353 vss.n15253 vss.n15252 21.67
R8354 vss.n15377 vss.n15376 21.67
R8355 vss.n15454 vss.n15453 21.67
R8356 vss.n15613 vss.n15612 21.67
R8357 vss.n15690 vss.n15689 21.67
R8358 vss.n15841 vss.n15840 21.67
R8359 vss.n16324 vss.n16323 21.67
R8360 vss.n16401 vss.n16400 21.67
R8361 vss.n16560 vss.n16559 21.67
R8362 vss.n16637 vss.n16636 21.67
R8363 vss.n21795 vss.n21664 21.645
R8364 vss.n3744 vss.n3613 21.645
R8365 vss.n21872 vss.n21871 21.62
R8366 vss.n3821 vss.n3820 21.62
R8367 vss.n12451 vss.n12450 21.455
R8368 vss.n12613 vss.n12612 21.455
R8369 vss.n14454 vss.n14453 21.455
R8370 vss.n14424 vss.n14423 21.455
R8371 vss.n14636 vss.n14635 21.455
R8372 vss.n13558 vss.n13557 21.455
R8373 vss.n15029 vss.n15028 21.455
R8374 vss.n10474 vss.n10473 21.455
R8375 vss.n13312 vss.n13311 21.455
R8376 vss.n14749 vss.n14748 21.455
R8377 vss.n14916 vss.n14915 21.455
R8378 vss.n14944 vss.n14943 21.455
R8379 vss.n14323 vss.n14322 21.455
R8380 vss.n13896 vss.n13895 21.455
R8381 vss.n13997 vss.n13996 21.455
R8382 vss.n11589 vss.n11588 21.455
R8383 vss.n11732 vss.n11731 21.455
R8384 vss.n11140 vss.n11139 21.455
R8385 vss.n10842 vss.n10841 21.455
R8386 vss.n10886 vss.n10885 21.455
R8387 vss.n11242 vss.n11241 21.455
R8388 vss.n11207 vss.n11206 21.455
R8389 vss.n12152 vss.n12151 21.455
R8390 vss.n12209 vss.n12208 21.455
R8391 vss.n22734 vss.n22732 21.245
R8392 vss.n22657 vss.n22655 21.245
R8393 vss.n22526 vss.n22524 21.245
R8394 vss.n22449 vss.n22447 21.245
R8395 vss.n22318 vss.n22316 21.245
R8396 vss.n22241 vss.n22239 21.245
R8397 vss.n22110 vss.n22108 21.245
R8398 vss.n17406 vss.n17404 21.245
R8399 vss.n21454 vss.n21452 21.245
R8400 vss.n21377 vss.n21375 21.245
R8401 vss.n21246 vss.n21244 21.245
R8402 vss.n21169 vss.n21167 21.245
R8403 vss.n21038 vss.n21036 21.245
R8404 vss.n20961 vss.n20959 21.245
R8405 vss.n8897 vss.n8895 21.245
R8406 vss.n8820 vss.n8818 21.245
R8407 vss.n8689 vss.n8687 21.245
R8408 vss.n8612 vss.n8610 21.245
R8409 vss.n8481 vss.n8479 21.245
R8410 vss.n8404 vss.n8402 21.245
R8411 vss.n8273 vss.n8271 21.245
R8412 vss.n8196 vss.n8194 21.245
R8413 vss.n8065 vss.n8063 21.245
R8414 vss.n7988 vss.n7986 21.245
R8415 vss.n7857 vss.n7855 21.245
R8416 vss.n7779 vss.n7777 21.245
R8417 vss.n7648 vss.n7646 21.245
R8418 vss.n7571 vss.n7569 21.245
R8419 vss.n21658 vss.n21657 21.219
R8420 vss.n3607 vss.n3606 21.219
R8421 vss.n20648 vss.n20647 20.82
R8422 vss.n20666 vss.n20665 20.82
R8423 vss.n7258 vss.n7257 20.82
R8424 vss.n7276 vss.n7275 20.82
R8425 vss.n1869 vss.n1868 20.82
R8426 vss.n1888 vss.n1887 20.82
R8427 vss.n2114 vss.n2113 20.82
R8428 vss.n2132 vss.n2131 20.82
R8429 vss.t13 vss.n2231 20.82
R8430 vss.n2358 vss.n2357 20.82
R8431 vss.n2376 vss.n2375 20.82
R8432 vss.n2602 vss.n2601 20.82
R8433 vss.n2621 vss.n2620 20.82
R8434 vss.n2840 vss.n2839 20.82
R8435 vss.n2859 vss.n2858 20.82
R8436 vss.t79 vss.n2987 20.82
R8437 vss.n3085 vss.n3084 20.82
R8438 vss.n3103 vss.n3102 20.82
R8439 vss.n3329 vss.n3328 20.82
R8440 vss.n3347 vss.n3346 20.82
R8441 vss.n330 vss.n329 20.82
R8442 vss.n349 vss.n348 20.82
R8443 vss.n575 vss.n574 20.82
R8444 vss.n593 vss.n592 20.82
R8445 vss.t303 vss.n692 20.82
R8446 vss.n819 vss.n818 20.82
R8447 vss.n837 vss.n836 20.82
R8448 vss.n1063 vss.n1062 20.82
R8449 vss.n1082 vss.n1081 20.82
R8450 vss.n1308 vss.n1307 20.82
R8451 vss.n23402 vss.n23401 20.82
R8452 vss.t285 vss.n23277 20.82
R8453 vss.n23177 vss.n23176 20.82
R8454 vss.n23159 vss.n23158 20.82
R8455 vss.n22933 vss.n22932 20.82
R8456 vss.n22914 vss.n22913 20.82
R8457 vss.n21772 vss.n21771 19.919
R8458 vss.n3721 vss.n3720 19.919
R8459 vss.n20493 vss.n20492 19.758
R8460 vss.n20584 vss.n20583 19.758
R8461 vss.n20722 vss.n20721 19.758
R8462 vss.n20807 vss.n20806 19.758
R8463 vss.n7103 vss.n7102 19.758
R8464 vss.n7194 vss.n7193 19.758
R8465 vss.n7332 vss.n7331 19.758
R8466 vss.n7417 vss.n7416 19.758
R8467 vss.n1716 vss.n1715 19.758
R8468 vss.n1805 vss.n1804 19.758
R8469 vss.n1947 vss.n1946 19.758
R8470 vss.n2044 vss.n2043 19.758
R8471 vss.n2192 vss.n2191 19.758
R8472 vss.n2288 vss.n2287 19.758
R8473 vss.n2436 vss.n2435 19.758
R8474 vss.n2533 vss.n2532 19.758
R8475 vss.n2680 vss.n2679 19.758
R8476 vss.n2777 vss.n2776 19.758
R8477 vss.n2919 vss.n2918 19.758
R8478 vss.n3016 vss.n3015 19.758
R8479 vss.n3163 vss.n3162 19.758
R8480 vss.n3260 vss.n3259 19.758
R8481 vss.n3403 vss.n3402 19.758
R8482 vss.n3470 vss.n3469 19.758
R8483 vss.n177 vss.n176 19.758
R8484 vss.n266 vss.n265 19.758
R8485 vss.n408 vss.n407 19.758
R8486 vss.n505 vss.n504 19.758
R8487 vss.n653 vss.n652 19.758
R8488 vss.n749 vss.n748 19.758
R8489 vss.n897 vss.n896 19.758
R8490 vss.n994 vss.n993 19.758
R8491 vss.n1141 vss.n1140 19.758
R8492 vss.n1238 vss.n1237 19.758
R8493 vss.n23333 vss.n23332 19.758
R8494 vss.n23236 vss.n23235 19.758
R8495 vss.n23089 vss.n23088 19.758
R8496 vss.n22992 vss.n22991 19.758
R8497 vss.n22850 vss.n22849 19.758
R8498 vss.n1445 vss.n1444 19.758
R8499 vss.n18976 vss.n17662 19.7
R8500 vss.n18920 vss.n17703 19.7
R8501 vss.n18853 vss.n17767 19.7
R8502 vss.n18803 vss.n17809 19.7
R8503 vss.n18736 vss.n17871 19.7
R8504 vss.n18679 vss.n17916 19.7
R8505 vss.n18612 vss.n17980 19.7
R8506 vss.n18562 vss.n18022 19.7
R8507 vss.n18495 vss.n18084 19.7
R8508 vss.n18438 vss.n18129 19.7
R8509 vss.n18371 vss.n18193 19.7
R8510 vss.n18321 vss.n18235 19.7
R8511 vss.n20246 vss.n19067 19.7
R8512 vss.n20196 vss.n19109 19.7
R8513 vss.n20122 vss.n19169 19.7
R8514 vss.n20066 vss.n19210 19.7
R8515 vss.n19999 vss.n19274 19.7
R8516 vss.n19949 vss.n19316 19.7
R8517 vss.n19875 vss.n19376 19.7
R8518 vss.n19819 vss.n19417 19.7
R8519 vss.n19752 vss.n19481 19.7
R8520 vss.n19702 vss.n19523 19.7
R8521 vss.n19628 vss.n19583 19.7
R8522 vss.n20337 vss.n20336 19.7
R8523 vss.n5586 vss.n4272 19.7
R8524 vss.n5530 vss.n4313 19.7
R8525 vss.n5463 vss.n4377 19.7
R8526 vss.n5413 vss.n4419 19.7
R8527 vss.n5346 vss.n4481 19.7
R8528 vss.n5289 vss.n4526 19.7
R8529 vss.n5222 vss.n4590 19.7
R8530 vss.n5172 vss.n4632 19.7
R8531 vss.n5105 vss.n4694 19.7
R8532 vss.n5048 vss.n4739 19.7
R8533 vss.n4981 vss.n4803 19.7
R8534 vss.n4931 vss.n4845 19.7
R8535 vss.n6856 vss.n5677 19.7
R8536 vss.n6806 vss.n5719 19.7
R8537 vss.n6732 vss.n5779 19.7
R8538 vss.n6676 vss.n5820 19.7
R8539 vss.n6609 vss.n5884 19.7
R8540 vss.n6559 vss.n5926 19.7
R8541 vss.n6485 vss.n5986 19.7
R8542 vss.n6429 vss.n6027 19.7
R8543 vss.n6362 vss.n6091 19.7
R8544 vss.n6312 vss.n6133 19.7
R8545 vss.n6238 vss.n6193 19.7
R8546 vss.n6947 vss.n6946 19.7
R8547 vss.n16736 vss.n16732 19.7
R8548 vss.n16833 vss.n16829 19.7
R8549 vss.n16966 vss.n16962 19.7
R8550 vss.n17067 vss.n17063 19.7
R8551 vss.n17202 vss.n17198 19.7
R8552 vss.n17323 vss.n17319 19.7
R8553 vss.n16013 vss.n16009 19.7
R8554 vss.n16113 vss.n16109 19.7
R8555 vss.n15285 vss.n15281 19.7
R8556 vss.n15352 vss.n15348 19.7
R8557 vss.n15486 vss.n15482 19.7
R8558 vss.n15589 vss.n15585 19.7
R8559 vss.n15722 vss.n15718 19.7
R8560 vss.n15813 vss.n15809 19.7
R8561 vss.n16433 vss.n16429 19.7
R8562 vss.n16536 vss.n16532 19.7
R8563 vss.n21763 vss.n21692 19.412
R8564 vss.n3712 vss.n3641 19.412
R8565 vss.n22625 vss.n22624 19.313
R8566 vss.n22550 vss.n22549 19.313
R8567 vss.n22417 vss.n22416 19.313
R8568 vss.n22342 vss.n22341 19.313
R8569 vss.n22209 vss.n22208 19.313
R8570 vss.n22134 vss.n22133 19.313
R8571 vss.n21553 vss.n21552 19.313
R8572 vss.n21478 vss.n21477 19.313
R8573 vss.n21345 vss.n21344 19.313
R8574 vss.n21270 vss.n21269 19.313
R8575 vss.n21137 vss.n21136 19.313
R8576 vss.n21062 vss.n21061 19.313
R8577 vss.n20929 vss.n20928 19.313
R8578 vss.n8788 vss.n8787 19.313
R8579 vss.n8713 vss.n8712 19.313
R8580 vss.n8580 vss.n8579 19.313
R8581 vss.n8505 vss.n8504 19.313
R8582 vss.n8372 vss.n8371 19.313
R8583 vss.n8297 vss.n8296 19.313
R8584 vss.n8164 vss.n8163 19.313
R8585 vss.n8089 vss.n8088 19.313
R8586 vss.n7956 vss.n7955 19.313
R8587 vss.n7881 vss.n7880 19.313
R8588 vss.n7747 vss.n7746 19.313
R8589 vss.n7672 vss.n7671 19.313
R8590 vss.n7539 vss.n7538 19.313
R8591 vss.n21695 vss.n21694 19.274
R8592 vss.n3644 vss.n3643 19.274
R8593 vss.n21780 vss.n21693 19.219
R8594 vss.n3729 vss.n3642 19.219
R8595 vss.n21787 vss.n21786 19.158
R8596 vss.n3736 vss.n3735 19.158
R8597 vss.n21721 vss.n21719 18.731
R8598 vss.n3670 vss.n3668 18.731
R8599 vss.n18988 vss.n17652 17.73
R8600 vss.n17718 vss.n17709 17.73
R8601 vss.n18864 vss.n17759 17.73
R8602 vss.n18792 vss.n17819 17.73
R8603 vss.n17867 vss.n17861 17.73
R8604 vss.n17931 vss.n17922 17.73
R8605 vss.n18623 vss.n17972 17.73
R8606 vss.n18551 vss.n18032 17.73
R8607 vss.n18080 vss.n18074 17.73
R8608 vss.n18144 vss.n18135 17.73
R8609 vss.n18382 vss.n18185 17.73
R8610 vss.n18310 vss.n18245 17.73
R8611 vss.n20257 vss.n19059 17.73
R8612 vss.n20185 vss.n19119 17.73
R8613 vss.n20134 vss.n19159 17.73
R8614 vss.n19225 vss.n19216 17.73
R8615 vss.n20010 vss.n19266 17.73
R8616 vss.n19938 vss.n19326 17.73
R8617 vss.n19887 vss.n19366 17.73
R8618 vss.n19432 vss.n19423 17.73
R8619 vss.n19763 vss.n19473 17.73
R8620 vss.n19691 vss.n19533 17.73
R8621 vss.n19640 vss.n19573 17.73
R8622 vss.n20330 vss.n17602 17.73
R8623 vss.n5598 vss.n4262 17.73
R8624 vss.n4328 vss.n4319 17.73
R8625 vss.n5474 vss.n4369 17.73
R8626 vss.n5402 vss.n4429 17.73
R8627 vss.n4477 vss.n4471 17.73
R8628 vss.n4541 vss.n4532 17.73
R8629 vss.n5233 vss.n4582 17.73
R8630 vss.n5161 vss.n4642 17.73
R8631 vss.n4690 vss.n4684 17.73
R8632 vss.n4754 vss.n4745 17.73
R8633 vss.n4992 vss.n4795 17.73
R8634 vss.n4920 vss.n4855 17.73
R8635 vss.n6867 vss.n5669 17.73
R8636 vss.n6795 vss.n5729 17.73
R8637 vss.n6744 vss.n5769 17.73
R8638 vss.n5835 vss.n5826 17.73
R8639 vss.n6620 vss.n5876 17.73
R8640 vss.n6548 vss.n5936 17.73
R8641 vss.n6497 vss.n5976 17.73
R8642 vss.n6042 vss.n6033 17.73
R8643 vss.n6373 vss.n6083 17.73
R8644 vss.n6301 vss.n6143 17.73
R8645 vss.n6250 vss.n6183 17.73
R8646 vss.n6940 vss.n4212 17.73
R8647 vss.n16718 vss.n16717 17.73
R8648 vss.n16843 vss.n16842 17.73
R8649 vss.n16948 vss.n16947 17.73
R8650 vss.n17077 vss.n17076 17.73
R8651 vss.n17184 vss.n17183 17.73
R8652 vss.n17279 vss.n17278 17.73
R8653 vss.n15887 vss.n15886 17.73
R8654 vss.n15995 vss.n15994 17.73
R8655 vss.n16123 vss.n16122 17.73
R8656 vss.n16231 vss.n16230 17.73
R8657 vss.n15267 vss.n15266 17.73
R8658 vss.n15363 vss.n15362 17.73
R8659 vss.n15468 vss.n15467 17.73
R8660 vss.n15599 vss.n15598 17.73
R8661 vss.n15704 vss.n15703 17.73
R8662 vss.n15827 vss.n15826 17.73
R8663 vss.n16310 vss.n16309 17.73
R8664 vss.n16415 vss.n16414 17.73
R8665 vss.n16546 vss.n16545 17.73
R8666 vss.n16651 vss.n16650 17.73
R8667 vss.n21883 vss.n21882 17.689
R8668 vss.n3832 vss.n3831 17.689
R8669 vss.n22748 vss.n22744 17.382
R8670 vss.n22643 vss.n22639 17.382
R8671 vss.n22540 vss.n22536 17.382
R8672 vss.n22435 vss.n22431 17.382
R8673 vss.n22332 vss.n22328 17.382
R8674 vss.n22227 vss.n22223 17.382
R8675 vss.n22124 vss.n22120 17.382
R8676 vss.n21571 vss.n21567 17.382
R8677 vss.n21468 vss.n21464 17.382
R8678 vss.n21363 vss.n21359 17.382
R8679 vss.n21260 vss.n21256 17.382
R8680 vss.n21155 vss.n21151 17.382
R8681 vss.n21052 vss.n21048 17.382
R8682 vss.n20947 vss.n20943 17.382
R8683 vss.n12071 vss.n12068 17.382
R8684 vss.n10800 vss.n10797 17.382
R8685 vss.n10963 vss.n10960 17.382
R8686 vss.n11003 vss.n11000 17.382
R8687 vss.n13853 vss.n13850 17.382
R8688 vss.n14074 vss.n14071 17.382
R8689 vss.n11720 vss.n11717 17.382
R8690 vss.n11064 vss.n11061 17.382
R8691 vss.n13351 vss.n13348 17.382
R8692 vss.n14696 vss.n14693 17.382
R8693 vss.n14189 vss.n14186 17.382
R8694 vss.n14231 vss.n14228 17.382
R8695 vss.n12871 vss.n12868 17.382
R8696 vss.n12920 vss.n12911 17.382
R8697 vss.n12466 vss.n12463 17.382
R8698 vss.n12507 vss.n12498 17.382
R8699 vss.n8911 vss.n8907 17.382
R8700 vss.n8806 vss.n8802 17.382
R8701 vss.n8703 vss.n8699 17.382
R8702 vss.n8598 vss.n8594 17.382
R8703 vss.n8495 vss.n8491 17.382
R8704 vss.n8390 vss.n8386 17.382
R8705 vss.n8287 vss.n8283 17.382
R8706 vss.n8182 vss.n8178 17.382
R8707 vss.n8079 vss.n8075 17.382
R8708 vss.n7974 vss.n7970 17.382
R8709 vss.n7871 vss.n7867 17.382
R8710 vss.n7765 vss.n7761 17.382
R8711 vss.n7662 vss.n7658 17.382
R8712 vss.n7557 vss.n7553 17.382
R8713 vss.n11687 vss.n11686 17.322
R8714 vss.n12261 vss.n12260 17.322
R8715 vss.n11937 vss.n11936 17.322
R8716 vss.n13944 vss.n13943 17.322
R8717 vss.n11528 vss.n11527 17.14
R8718 vss.n12367 vss.n12366 17.14
R8719 vss.n13168 vss.n13167 17.14
R8720 vss.n12926 vss.n12925 17.14
R8721 vss.n10709 vss.n10708 17.14
R8722 vss.n12998 vss.n12997 17.14
R8723 vss.n10562 vss.n10561 17.14
R8724 vss.n12347 vss.n12346 17.14
R8725 vss.n11507 vss.n11506 17.14
R8726 vss.n9163 vss.t315 16.877
R8727 vss.n9171 vss.t10 16.788
R8728 vss.n17530 vss.n17529 16.53
R8729 vss.n17530 vss.t280 16.53
R8730 vss.n17516 vss.t236 16.53
R8731 vss.n17516 vss.t234 16.53
R8732 vss.n17504 vss.t302 16.53
R8733 vss.n17504 vss.n17503 16.53
R8734 vss.n17498 vss.t164 16.53
R8735 vss.n4140 vss.n4139 16.53
R8736 vss.n4140 vss.t58 16.53
R8737 vss.n4126 vss.t46 16.53
R8738 vss.n4126 vss.t48 16.53
R8739 vss.n4114 vss.t28 16.53
R8740 vss.n4114 vss.n4113 16.53
R8741 vss.n4108 vss.t209 16.53
R8742 vss.n1786 vss.n1785 16.53
R8743 vss.n1786 vss.t62 16.53
R8744 vss.n1626 vss.t68 16.53
R8745 vss.n1626 vss.t54 16.53
R8746 vss.n1625 vss.t76 16.53
R8747 vss.n1625 vss.t22 16.53
R8748 vss.n1624 vss.t26 16.53
R8749 vss.n1624 vss.t34 16.53
R8750 vss.n1599 vss.t18 16.53
R8751 vss.n1599 vss.t14 16.53
R8752 vss.n2297 vss.t66 16.53
R8753 vss.n2297 vss.t74 16.53
R8754 vss.n2398 vss.t56 16.53
R8755 vss.n2398 vss.t20 16.53
R8756 vss.n1574 vss.t52 16.53
R8757 vss.n1574 vss.t36 16.53
R8758 vss.n1561 vss.t82 16.53
R8759 vss.n1561 vss.t60 16.53
R8760 vss.n1548 vss.t64 16.53
R8761 vss.n1548 vss.t72 16.53
R8762 vss.n1547 vss.t40 16.53
R8763 vss.n1547 vss.t44 16.53
R8764 vss.n2913 vss.t24 16.53
R8765 vss.n2913 vss.t32 16.53
R8766 vss.n1516 vss.t80 16.53
R8767 vss.n1516 vss.t84 16.53
R8768 vss.n1491 vss.t16 16.53
R8769 vss.n1491 vss.t70 16.53
R8770 vss.n1490 vss.t38 16.53
R8771 vss.n1490 vss.t42 16.53
R8772 vss.n1489 vss.t50 16.53
R8773 vss.n1489 vss.t30 16.53
R8774 vss.n3447 vss.t78 16.53
R8775 vss.n3453 vss.n3452 16.53
R8776 vss.n3453 vss.t89 16.53
R8777 vss.n247 vss.n246 16.53
R8778 vss.n247 vss.t244 16.53
R8779 vss.n87 vss.t278 16.53
R8780 vss.n87 vss.t264 16.53
R8781 vss.n86 vss.t262 16.53
R8782 vss.n86 vss.t276 16.53
R8783 vss.n85 vss.t294 16.53
R8784 vss.n85 vss.t238 16.53
R8785 vss.n60 vss.t282 16.53
R8786 vss.n60 vss.t304 16.53
R8787 vss.n758 vss.t256 16.53
R8788 vss.n758 vss.t250 16.53
R8789 vss.n859 vss.t266 16.53
R8790 vss.n859 vss.t272 16.53
R8791 vss.n35 vss.t296 16.53
R8792 vss.n35 vss.t290 16.53
R8793 vss.n22 vss.t284 16.53
R8794 vss.n22 vss.t260 16.53
R8795 vss.n9 vss.t240 16.53
R8796 vss.n9 vss.t252 16.53
R8797 vss.n8 vss.t248 16.53
R8798 vss.n8 vss.t300 16.53
R8799 vss.n1336 vss.t298 16.53
R8800 vss.n1336 vss.t268 16.53
R8801 vss.n1337 vss.t286 16.53
R8802 vss.n1337 vss.t242 16.53
R8803 vss.n1362 vss.t258 16.53
R8804 vss.n1362 vss.t254 16.53
R8805 vss.n1363 vss.t246 16.53
R8806 vss.n1363 vss.t274 16.53
R8807 vss.n1364 vss.t270 16.53
R8808 vss.n1364 vss.t292 16.53
R8809 vss.n1422 vss.t288 16.53
R8810 vss.n1428 vss.n1427 16.53
R8811 vss.n1428 vss.t98 16.53
R8812 vss.n20452 vss.n20447 16.465
R8813 vss.n20634 vss.n20629 16.465
R8814 vss.n20682 vss.n20677 16.465
R8815 vss.n20858 vss.n20853 16.465
R8816 vss.n7062 vss.n7057 16.465
R8817 vss.n7244 vss.n7239 16.465
R8818 vss.n7292 vss.n7287 16.465
R8819 vss.n7468 vss.n7463 16.465
R8820 vss.n1855 vss.n1850 16.465
R8821 vss.n1905 vss.n1899 16.465
R8822 vss.n2098 vss.n2092 16.465
R8823 vss.n2149 vss.n2143 16.465
R8824 vss.n2343 vss.n2337 16.465
R8825 vss.n2393 vss.n2387 16.465
R8826 vss.n2587 vss.n2581 16.465
R8827 vss.n2638 vss.n2632 16.465
R8828 vss.n2829 vss.n2824 16.465
R8829 vss.n2876 vss.n2870 16.465
R8830 vss.n3070 vss.n3064 16.465
R8831 vss.n3121 vss.n3115 16.465
R8832 vss.n3314 vss.n3308 16.465
R8833 vss.n3363 vss.n3358 16.465
R8834 vss.n316 vss.n311 16.465
R8835 vss.n366 vss.n360 16.465
R8836 vss.n559 vss.n553 16.465
R8837 vss.n610 vss.n604 16.465
R8838 vss.n804 vss.n798 16.465
R8839 vss.n854 vss.n848 16.465
R8840 vss.n1048 vss.n1042 16.465
R8841 vss.n1099 vss.n1093 16.465
R8842 vss.n1293 vss.n1287 16.465
R8843 vss.n23387 vss.n23381 16.465
R8844 vss.n23194 vss.n23188 16.465
R8845 vss.n23143 vss.n23137 16.465
R8846 vss.n22950 vss.n22944 16.465
R8847 vss.n22900 vss.n22895 16.465
R8848 vss.n14134 vss.n14133 16.219
R8849 vss.n12274 vss.n12273 16.219
R8850 vss.n10464 vss.n10463 16.219
R8851 vss.n10605 vss.n10604 16.219
R8852 vss.n18988 vss.n17654 15.76
R8853 vss.n18916 vss.n17709 15.76
R8854 vss.n18860 vss.n17759 15.76
R8855 vss.n18796 vss.n17819 15.76
R8856 vss.n18740 vss.n17867 15.76
R8857 vss.n18675 vss.n17922 15.76
R8858 vss.n18619 vss.n17972 15.76
R8859 vss.n18555 vss.n18032 15.76
R8860 vss.n18499 vss.n18080 15.76
R8861 vss.n18434 vss.n18135 15.76
R8862 vss.n18378 vss.n18185 15.76
R8863 vss.n18314 vss.n18245 15.76
R8864 vss.n20253 vss.n19059 15.76
R8865 vss.n20189 vss.n19119 15.76
R8866 vss.n20134 vss.n19161 15.76
R8867 vss.n20062 vss.n19216 15.76
R8868 vss.n20006 vss.n19266 15.76
R8869 vss.n19942 vss.n19326 15.76
R8870 vss.n19887 vss.n19368 15.76
R8871 vss.n19815 vss.n19423 15.76
R8872 vss.n19759 vss.n19473 15.76
R8873 vss.n19695 vss.n19533 15.76
R8874 vss.n19640 vss.n19575 15.76
R8875 vss.n5598 vss.n4264 15.76
R8876 vss.n5526 vss.n4319 15.76
R8877 vss.n5470 vss.n4369 15.76
R8878 vss.n5406 vss.n4429 15.76
R8879 vss.n5350 vss.n4477 15.76
R8880 vss.n5285 vss.n4532 15.76
R8881 vss.n5229 vss.n4582 15.76
R8882 vss.n5165 vss.n4642 15.76
R8883 vss.n5109 vss.n4690 15.76
R8884 vss.n5044 vss.n4745 15.76
R8885 vss.n4988 vss.n4795 15.76
R8886 vss.n4924 vss.n4855 15.76
R8887 vss.n6863 vss.n5669 15.76
R8888 vss.n6799 vss.n5729 15.76
R8889 vss.n6744 vss.n5771 15.76
R8890 vss.n6672 vss.n5826 15.76
R8891 vss.n6616 vss.n5876 15.76
R8892 vss.n6552 vss.n5936 15.76
R8893 vss.n6497 vss.n5978 15.76
R8894 vss.n6425 vss.n6033 15.76
R8895 vss.n6369 vss.n6083 15.76
R8896 vss.n6305 vss.n6143 15.76
R8897 vss.n6250 vss.n6185 15.76
R8898 vss.n16722 vss.n16718 15.76
R8899 vss.n16847 vss.n16843 15.76
R8900 vss.n16952 vss.n16948 15.76
R8901 vss.n17081 vss.n17077 15.76
R8902 vss.n17188 vss.n17184 15.76
R8903 vss.n17283 vss.n17279 15.76
R8904 vss.n15891 vss.n15887 15.76
R8905 vss.n15999 vss.n15995 15.76
R8906 vss.n16127 vss.n16123 15.76
R8907 vss.n16235 vss.n16231 15.76
R8908 vss.n15271 vss.n15267 15.76
R8909 vss.n15367 vss.n15363 15.76
R8910 vss.n15472 vss.n15468 15.76
R8911 vss.n15603 vss.n15599 15.76
R8912 vss.n15708 vss.n15704 15.76
R8913 vss.n15831 vss.n15827 15.76
R8914 vss.n16314 vss.n16310 15.76
R8915 vss.n16419 vss.n16415 15.76
R8916 vss.n16550 vss.n16546 15.76
R8917 vss.n16655 vss.n16651 15.76
R8918 vss.n21882 vss.n21881 15.724
R8919 vss.n3831 vss.n3830 15.724
R8920 vss.n22744 vss.n22743 15.45
R8921 vss.n22639 vss.n22638 15.45
R8922 vss.n22536 vss.n22535 15.45
R8923 vss.n22431 vss.n22430 15.45
R8924 vss.n22328 vss.n22327 15.45
R8925 vss.n22223 vss.n22222 15.45
R8926 vss.n22120 vss.n22119 15.45
R8927 vss.n21567 vss.n21566 15.45
R8928 vss.n21464 vss.n21463 15.45
R8929 vss.n21359 vss.n21358 15.45
R8930 vss.n21256 vss.n21255 15.45
R8931 vss.n21151 vss.n21150 15.45
R8932 vss.n21048 vss.n21047 15.45
R8933 vss.n20943 vss.n20942 15.45
R8934 vss.n8907 vss.n8906 15.45
R8935 vss.n8802 vss.n8801 15.45
R8936 vss.n8699 vss.n8698 15.45
R8937 vss.n8594 vss.n8593 15.45
R8938 vss.n8491 vss.n8490 15.45
R8939 vss.n8386 vss.n8385 15.45
R8940 vss.n8283 vss.n8282 15.45
R8941 vss.n8178 vss.n8177 15.45
R8942 vss.n8075 vss.n8074 15.45
R8943 vss.n7970 vss.n7969 15.45
R8944 vss.n7867 vss.n7866 15.45
R8945 vss.n7761 vss.n7760 15.45
R8946 vss.n7658 vss.n7657 15.45
R8947 vss.n7553 vss.n7552 15.45
R8948 vss.n13708 vss.n13707 15.29
R8949 vss.n13031 vss.n13030 15.29
R8950 vss.n14347 vss.n14346 15.29
R8951 vss.n14480 vss.n14479 15.29
R8952 vss.n10756 vss.n10755 15.29
R8953 vss.n12793 vss.n12792 15.29
R8954 vss.n13042 vss.n13041 15.29
R8955 vss.n13695 vss.n13694 15.29
R8956 vss.n12135 vss.n12134 15.272
R8957 vss.n13263 vss.n13262 15.272
R8958 vss.n12122 vss.n12112 15.272
R8959 vss.n13276 vss.n13266 15.272
R8960 vss.n20331 vss.n20330 15.113
R8961 vss.n6941 vss.n6940 15.113
R8962 vss.n14999 vss.n14998 14.628
R8963 vss.n13957 vss.n13956 14.628
R8964 vss.n11810 vss.n11809 14.628
R8965 vss.n14571 vss.n14570 14.628
R8966 vss.n13631 vss.n13630 14.628
R8967 vss.n13683 vss.n13682 14.628
R8968 vss.n11380 vss.n11379 14.628
R8969 vss.n11366 vss.n11365 14.628
R8970 vss.n11309 vss.n11308 14.628
R8971 vss.n12397 vss.n12396 14.628
R8972 vss.n14707 vss.n14706 14.628
R8973 vss.n13444 vss.n13443 14.628
R8974 vss.n13019 vss.n13018 14.628
R8975 vss.n10576 vss.n10575 14.628
R8976 vss.n10733 vss.n10732 14.628
R8977 vss.n12029 vss.n12028 14.628
R8978 vss.n13922 vss.n13921 14.35
R8979 vss.n11268 vss.n11267 14.35
R8980 vss.n13424 vss.n13423 14.35
R8981 vss.n13609 vss.n13608 14.349
R8982 vss.n11021 vss.n11020 14.349
R8983 vss.n12234 vss.n12233 14.349
R8984 vss.n12515 vss.n12514 14.349
R8985 vss.n13195 vss.n13194 14.349
R8986 vss.n13619 vss.n13618 14.349
R8987 vss.n13433 vss.n13432 14.349
R8988 vss.n11391 vss.n11390 14.349
R8989 vss.n11648 vss.n11647 14.349
R8990 vss.n14583 vss.n14582 14.272
R8991 vss.n14719 vss.n14718 14.272
R8992 vss.n14989 vss.n14988 14.272
R8993 vss.n14717 vss.n14716 14.272
R8994 vss.n14581 vss.n14580 14.272
R8995 vss.n11682 vss.n11681 14.272
R8996 vss.n11684 vss.n11683 14.272
R8997 vss.n12257 vss.n12256 14.272
R8998 vss.n11934 vss.n11933 14.272
R8999 vss.n10533 vss.n10532 14.272
R9000 vss.n21670 vss.n21660 14.085
R9001 vss.n3619 vss.n3609 14.085
R9002 vss.n20529 vss.n20526 13.88
R9003 vss.n20557 vss.n20554 13.88
R9004 vss.n20588 vss.t279 13.88
R9005 vss.n20726 vss.t301 13.88
R9006 vss.n20758 vss.n20755 13.88
R9007 vss.n20779 vss.n20776 13.88
R9008 vss.n7139 vss.n7136 13.88
R9009 vss.n7167 vss.n7164 13.88
R9010 vss.n7198 vss.t57 13.88
R9011 vss.n7336 vss.t27 13.88
R9012 vss.n7368 vss.n7365 13.88
R9013 vss.n7389 vss.n7386 13.88
R9014 vss.n1755 vss.n1752 13.88
R9015 vss.n1776 vss.n1773 13.88
R9016 vss.n1986 vss.n1981 13.88
R9017 vss.n2016 vss.n2011 13.88
R9018 vss.n2231 vss.n2226 13.88
R9019 vss.n2260 vss.n2255 13.88
R9020 vss.n2277 vss.t65 13.88
R9021 vss.n2475 vss.n2470 13.88
R9022 vss.n2504 vss.n2499 13.88
R9023 vss.n2538 vss.t35 13.88
R9024 vss.n2685 vss.t63 13.88
R9025 vss.n2720 vss.n2715 13.88
R9026 vss.n2749 vss.n2744 13.88
R9027 vss.n2940 vss.t31 13.88
R9028 vss.n2958 vss.n2953 13.88
R9029 vss.n2987 vss.n2982 13.88
R9030 vss.n3202 vss.n3197 13.88
R9031 vss.n3232 vss.n3227 13.88
R9032 vss.n15204 vss.n15201 13.88
R9033 vss.n15185 vss.n15182 13.88
R9034 vss.n216 vss.n213 13.88
R9035 vss.n237 vss.n234 13.88
R9036 vss.n447 vss.n442 13.88
R9037 vss.n477 vss.n472 13.88
R9038 vss.n692 vss.n687 13.88
R9039 vss.n721 vss.n716 13.88
R9040 vss.n738 vss.t255 13.88
R9041 vss.n936 vss.n931 13.88
R9042 vss.n965 vss.n960 13.88
R9043 vss.n999 vss.t289 13.88
R9044 vss.n1146 vss.t239 13.88
R9045 vss.n1181 vss.n1176 13.88
R9046 vss.n1210 vss.n1205 13.88
R9047 vss.n23322 vss.t267 13.88
R9048 vss.n23304 vss.n23299 13.88
R9049 vss.n23277 vss.n23272 13.88
R9050 vss.n23060 vss.n23055 13.88
R9051 vss.n23032 vss.n23027 13.88
R9052 vss.n1397 vss.n1394 13.88
R9053 vss.n22819 vss.n22816 13.88
R9054 vss.n18980 vss.n17662 13.79
R9055 vss.n18920 vss.n17707 13.79
R9056 vss.n17767 vss.n17761 13.79
R9057 vss.n17818 vss.n17809 13.79
R9058 vss.n18736 vss.n17868 13.79
R9059 vss.n18679 vss.n17920 13.79
R9060 vss.n17980 vss.n17974 13.79
R9061 vss.n18031 vss.n18022 13.79
R9062 vss.n18495 vss.n18081 13.79
R9063 vss.n18438 vss.n18133 13.79
R9064 vss.n18193 vss.n18187 13.79
R9065 vss.n18244 vss.n18235 13.79
R9066 vss.n19067 vss.n19061 13.79
R9067 vss.n19118 vss.n19109 13.79
R9068 vss.n20126 vss.n19169 13.79
R9069 vss.n20066 vss.n19214 13.79
R9070 vss.n19274 vss.n19268 13.79
R9071 vss.n19325 vss.n19316 13.79
R9072 vss.n19879 vss.n19376 13.79
R9073 vss.n19819 vss.n19421 13.79
R9074 vss.n19481 vss.n19475 13.79
R9075 vss.n19532 vss.n19523 13.79
R9076 vss.n19632 vss.n19583 13.79
R9077 vss.n5590 vss.n4272 13.79
R9078 vss.n5530 vss.n4317 13.79
R9079 vss.n4377 vss.n4371 13.79
R9080 vss.n4428 vss.n4419 13.79
R9081 vss.n5346 vss.n4478 13.79
R9082 vss.n5289 vss.n4530 13.79
R9083 vss.n4590 vss.n4584 13.79
R9084 vss.n4641 vss.n4632 13.79
R9085 vss.n5105 vss.n4691 13.79
R9086 vss.n5048 vss.n4743 13.79
R9087 vss.n4803 vss.n4797 13.79
R9088 vss.n4854 vss.n4845 13.79
R9089 vss.n5677 vss.n5671 13.79
R9090 vss.n5728 vss.n5719 13.79
R9091 vss.n6736 vss.n5779 13.79
R9092 vss.n6676 vss.n5824 13.79
R9093 vss.n5884 vss.n5878 13.79
R9094 vss.n5935 vss.n5926 13.79
R9095 vss.n6489 vss.n5986 13.79
R9096 vss.n6429 vss.n6031 13.79
R9097 vss.n6091 vss.n6085 13.79
R9098 vss.n6142 vss.n6133 13.79
R9099 vss.n6242 vss.n6193 13.79
R9100 vss.n16732 vss.n16731 13.79
R9101 vss.n16829 vss.n16828 13.79
R9102 vss.n16962 vss.n16961 13.79
R9103 vss.n17063 vss.n17062 13.79
R9104 vss.n17198 vss.n17197 13.79
R9105 vss.n17319 vss.n17318 13.79
R9106 vss.n16009 vss.n16008 13.79
R9107 vss.n16109 vss.n16108 13.79
R9108 vss.n15281 vss.n15280 13.79
R9109 vss.n15348 vss.n15347 13.79
R9110 vss.n15482 vss.n15481 13.79
R9111 vss.n15585 vss.n15584 13.79
R9112 vss.n15718 vss.n15717 13.79
R9113 vss.n15809 vss.n15808 13.79
R9114 vss.n16429 vss.n16428 13.79
R9115 vss.n16532 vss.n16531 13.79
R9116 vss.n20659 vss.n20658 13.552
R9117 vss.n21745 vss.n21712 13.552
R9118 vss.n21730 vss.n21729 13.552
R9119 vss.n21737 vss.n21714 13.552
R9120 vss.n21676 vss.n21662 13.552
R9121 vss.n21798 vss.n21797 13.552
R9122 vss.n14809 vss.n14808 13.552
R9123 vss.n3694 vss.n3661 13.552
R9124 vss.n3679 vss.n3678 13.552
R9125 vss.n3686 vss.n3663 13.552
R9126 vss.n3625 vss.n3611 13.552
R9127 vss.n3747 vss.n3746 13.552
R9128 vss.n7269 vss.n7268 13.552
R9129 vss.n1545 vss.n1544 13.552
R9130 vss.n2845 vss.n2844 13.552
R9131 vss.n22629 vss.n22625 13.519
R9132 vss.n22554 vss.n22550 13.519
R9133 vss.n22421 vss.n22417 13.519
R9134 vss.n22346 vss.n22342 13.519
R9135 vss.n22213 vss.n22209 13.519
R9136 vss.n22138 vss.n22134 13.519
R9137 vss.n21557 vss.n21553 13.519
R9138 vss.n21482 vss.n21478 13.519
R9139 vss.n21349 vss.n21345 13.519
R9140 vss.n21274 vss.n21270 13.519
R9141 vss.n21141 vss.n21137 13.519
R9142 vss.n21066 vss.n21062 13.519
R9143 vss.n20933 vss.n20929 13.519
R9144 vss.n8792 vss.n8788 13.519
R9145 vss.n8717 vss.n8713 13.519
R9146 vss.n8584 vss.n8580 13.519
R9147 vss.n8509 vss.n8505 13.519
R9148 vss.n8376 vss.n8372 13.519
R9149 vss.n8301 vss.n8297 13.519
R9150 vss.n8168 vss.n8164 13.519
R9151 vss.n8093 vss.n8089 13.519
R9152 vss.n7960 vss.n7956 13.519
R9153 vss.n7885 vss.n7881 13.519
R9154 vss.n7751 vss.n7747 13.519
R9155 vss.n7676 vss.n7672 13.519
R9156 vss.n7543 vss.n7539 13.519
R9157 vss.n17539 vss.n17538 13.176
R9158 vss.n17494 vss.n17493 13.176
R9159 vss.n4149 vss.n4148 13.176
R9160 vss.n4104 vss.n4103 13.176
R9161 vss.n3443 vss.n3442 13.176
R9162 vss.n1418 vss.n1417 13.176
R9163 vss.n20509 vss.n20508 13.172
R9164 vss.n20569 vss.n20568 13.172
R9165 vss.n20737 vss.n20736 13.172
R9166 vss.n20791 vss.n20790 13.172
R9167 vss.n7119 vss.n7118 13.172
R9168 vss.n7179 vss.n7178 13.172
R9169 vss.n7347 vss.n7346 13.172
R9170 vss.n7401 vss.n7400 13.172
R9171 vss.n1731 vss.n1730 13.172
R9172 vss.n1790 vss.n1789 13.172
R9173 vss.n1963 vss.n1962 13.172
R9174 vss.n2028 vss.n2027 13.172
R9175 vss.n2208 vss.n2207 13.172
R9176 vss.n2272 vss.n2271 13.172
R9177 vss.n2452 vss.n2451 13.172
R9178 vss.n2517 vss.n2516 13.172
R9179 vss.n2696 vss.n2695 13.172
R9180 vss.n2761 vss.n2760 13.172
R9181 vss.n2935 vss.n2934 13.172
R9182 vss.n2999 vss.n2998 13.172
R9183 vss.n3179 vss.n3178 13.172
R9184 vss.n3244 vss.n3243 13.172
R9185 vss.n3418 vss.n3417 13.172
R9186 vss.n3459 vss.n3458 13.172
R9187 vss.n192 vss.n191 13.172
R9188 vss.n251 vss.n250 13.172
R9189 vss.n424 vss.n423 13.172
R9190 vss.n489 vss.n488 13.172
R9191 vss.n669 vss.n668 13.172
R9192 vss.n733 vss.n732 13.172
R9193 vss.n913 vss.n912 13.172
R9194 vss.n978 vss.n977 13.172
R9195 vss.n1157 vss.n1156 13.172
R9196 vss.n1222 vss.n1221 13.172
R9197 vss.n23317 vss.n23316 13.172
R9198 vss.n23253 vss.n23252 13.172
R9199 vss.n23073 vss.n23072 13.172
R9200 vss.n23008 vss.n23007 13.172
R9201 vss.n22833 vss.n22832 13.172
R9202 vss.n1434 vss.n1433 13.172
R9203 vss.n9128 vss.n9127 12.805
R9204 vss.n20541 vss.n20539 12.8
R9205 vss.n20541 vss.n20540 12.8
R9206 vss.n20767 vss.n20765 12.8
R9207 vss.n20767 vss.n20766 12.8
R9208 vss.n10910 vss.n10906 12.8
R9209 vss.n10910 vss.n10909 12.8
R9210 vss.n14384 vss.n14380 12.8
R9211 vss.n14384 vss.n14383 12.8
R9212 vss.n11584 vss.n11580 12.8
R9213 vss.n11584 vss.n11583 12.8
R9214 vss.n13591 vss.n13587 12.8
R9215 vss.n13591 vss.n13590 12.8
R9216 vss.n14849 vss.n14845 12.8
R9217 vss.n14849 vss.n14848 12.8
R9218 vss.n12726 vss.n12722 12.8
R9219 vss.n12726 vss.n12725 12.8
R9220 vss.n7151 vss.n7149 12.8
R9221 vss.n7151 vss.n7150 12.8
R9222 vss.n7377 vss.n7375 12.8
R9223 vss.n7377 vss.n7376 12.8
R9224 vss.n1764 vss.n1762 12.8
R9225 vss.n1764 vss.n1763 12.8
R9226 vss.n1999 vss.n1997 12.8
R9227 vss.n1999 vss.n1998 12.8
R9228 vss.n2243 vss.n2241 12.8
R9229 vss.n2243 vss.n2242 12.8
R9230 vss.n2487 vss.n2485 12.8
R9231 vss.n2487 vss.n2486 12.8
R9232 vss.n2732 vss.n2730 12.8
R9233 vss.n2732 vss.n2731 12.8
R9234 vss.n2970 vss.n2968 12.8
R9235 vss.n2970 vss.n2969 12.8
R9236 vss.n3214 vss.n3212 12.8
R9237 vss.n3214 vss.n3213 12.8
R9238 vss.n15193 vss.n15191 12.8
R9239 vss.n15193 vss.n15192 12.8
R9240 vss.n225 vss.n223 12.8
R9241 vss.n225 vss.n224 12.8
R9242 vss.n460 vss.n458 12.8
R9243 vss.n460 vss.n459 12.8
R9244 vss.n704 vss.n702 12.8
R9245 vss.n704 vss.n703 12.8
R9246 vss.n948 vss.n946 12.8
R9247 vss.n948 vss.n947 12.8
R9248 vss.n1193 vss.n1191 12.8
R9249 vss.n1193 vss.n1192 12.8
R9250 vss.n23288 vss.n23286 12.8
R9251 vss.n23288 vss.n23287 12.8
R9252 vss.n23044 vss.n23042 12.8
R9253 vss.n23044 vss.n23043 12.8
R9254 vss.n22827 vss.n22825 12.8
R9255 vss.n22827 vss.n22826 12.8
R9256 vss.n13115 vss.n13114 12.678
R9257 vss.n13664 vss.n13663 12.678
R9258 vss.n14980 vss.n14979 12.678
R9259 vss.n13142 vss.n13141 12.678
R9260 vss.n13651 vss.n13650 12.678
R9261 vss.n14060 vss.n14059 12.678
R9262 vss.n11475 vss.n11474 12.678
R9263 vss.n11693 vss.n11692 12.678
R9264 vss.n14561 vss.n14560 12.678
R9265 vss.n14098 vss.n14097 12.678
R9266 vss.n13748 vss.n13747 12.678
R9267 vss.n11445 vss.n11444 12.678
R9268 vss.n11854 vss.n11853 12.678
R9269 vss.n10931 vss.n10930 12.678
R9270 vss.n12407 vss.n12406 12.678
R9271 vss.n10670 vss.n10669 12.678
R9272 vss.n12324 vss.n12323 12.678
R9273 vss.n11485 vss.n11484 12.678
R9274 vss.n13373 vss.n13372 12.678
R9275 vss.n13456 vss.n13455 12.678
R9276 vss.n13087 vss.n13086 12.678
R9277 vss.n10640 vss.n10639 12.678
R9278 vss.n12309 vss.n12308 12.678
R9279 vss.n10806 vss.n10805 12.678
R9280 vss.n20296 vss.n17616 12.531
R9281 vss.n20297 vss.n20296 12.531
R9282 vss.n6906 vss.n4226 12.531
R9283 vss.n6907 vss.n6906 12.531
R9284 vss.n13762 vss.n13761 12.437
R9285 vss.n13763 vss.n13762 12.437
R9286 vss.n10991 vss.n10990 12.437
R9287 vss.n10990 vss.n10989 12.437
R9288 vss.n11536 vss.n11535 12.437
R9289 vss.n11535 vss.n11534 12.437
R9290 vss.n10717 vss.n10716 12.437
R9291 vss.n12090 vss.n12089 12.437
R9292 vss.n12089 vss.n12088 12.437
R9293 vss.n12376 vss.n12375 12.437
R9294 vss.n12375 vss.n12374 12.437
R9295 vss.n12338 vss.n12337 12.437
R9296 vss.n13178 vss.n13177 12.437
R9297 vss.n13177 vss.n13176 12.437
R9298 vss.n12937 vss.n12936 12.437
R9299 vss.n12968 vss.n12967 12.437
R9300 vss.n12967 vss.n12966 12.437
R9301 vss.n13549 vss.n13548 12.437
R9302 vss.n13550 vss.n13549 12.437
R9303 vss.n12936 vss.n12935 12.437
R9304 vss.n10716 vss.n10715 12.437
R9305 vss.n13007 vss.n13006 12.437
R9306 vss.n13006 vss.n13005 12.437
R9307 vss.n10554 vss.n10553 12.437
R9308 vss.n10555 vss.n10554 12.437
R9309 vss.n12339 vss.n12338 12.437
R9310 vss.n11499 vss.n11498 12.437
R9311 vss.n11500 vss.n11499 12.437
R9312 vss.n18992 vss.n17645 11.82
R9313 vss.n18909 vss.n17719 11.82
R9314 vss.n18872 vss.n17752 11.82
R9315 vss.n18784 vss.n17822 11.82
R9316 vss.n18747 vss.n17859 11.82
R9317 vss.n18668 vss.n17932 11.82
R9318 vss.n18631 vss.n17965 11.82
R9319 vss.n18543 vss.n18035 11.82
R9320 vss.n18506 vss.n18072 11.82
R9321 vss.n18427 vss.n18145 11.82
R9322 vss.n18390 vss.n18178 11.82
R9323 vss.n18302 vss.n18248 11.82
R9324 vss.n20265 vss.n19051 11.82
R9325 vss.n20177 vss.n19122 11.82
R9326 vss.n20138 vss.n19152 11.82
R9327 vss.n20055 vss.n19226 11.82
R9328 vss.n20018 vss.n19259 11.82
R9329 vss.n19930 vss.n19329 11.82
R9330 vss.n19891 vss.n19359 11.82
R9331 vss.n19808 vss.n19433 11.82
R9332 vss.n19771 vss.n19466 11.82
R9333 vss.n19683 vss.n19536 11.82
R9334 vss.n19644 vss.n19566 11.82
R9335 vss.n20326 vss.n20325 11.82
R9336 vss.n5602 vss.n4255 11.82
R9337 vss.n5519 vss.n4329 11.82
R9338 vss.n5482 vss.n4362 11.82
R9339 vss.n5394 vss.n4432 11.82
R9340 vss.n5357 vss.n4469 11.82
R9341 vss.n5278 vss.n4542 11.82
R9342 vss.n5241 vss.n4575 11.82
R9343 vss.n5153 vss.n4645 11.82
R9344 vss.n5116 vss.n4682 11.82
R9345 vss.n5037 vss.n4755 11.82
R9346 vss.n5000 vss.n4788 11.82
R9347 vss.n4912 vss.n4858 11.82
R9348 vss.n6875 vss.n5661 11.82
R9349 vss.n6787 vss.n5732 11.82
R9350 vss.n6748 vss.n5762 11.82
R9351 vss.n6665 vss.n5836 11.82
R9352 vss.n6628 vss.n5869 11.82
R9353 vss.n6540 vss.n5939 11.82
R9354 vss.n6501 vss.n5969 11.82
R9355 vss.n6418 vss.n6043 11.82
R9356 vss.n6381 vss.n6076 11.82
R9357 vss.n6293 vss.n6146 11.82
R9358 vss.n6254 vss.n6176 11.82
R9359 vss.n6936 vss.n6935 11.82
R9360 vss.n16708 vss.n16704 11.82
R9361 vss.n16859 vss.n16855 11.82
R9362 vss.n16938 vss.n16934 11.82
R9363 vss.n17095 vss.n17091 11.82
R9364 vss.n17174 vss.n17170 11.82
R9365 vss.n17312 vss.n17308 11.82
R9366 vss.n15905 vss.n15901 11.82
R9367 vss.n15985 vss.n15981 11.82
R9368 vss.n16141 vss.n16137 11.82
R9369 vss.n16221 vss.n16217 11.82
R9370 vss.n15257 vss.n15253 11.82
R9371 vss.n15381 vss.n15377 11.82
R9372 vss.n15458 vss.n15454 11.82
R9373 vss.n15617 vss.n15613 11.82
R9374 vss.n15694 vss.n15690 11.82
R9375 vss.n15845 vss.n15841 11.82
R9376 vss.n16328 vss.n16324 11.82
R9377 vss.n16405 vss.n16401 11.82
R9378 vss.n16564 vss.n16560 11.82
R9379 vss.n16641 vss.n16637 11.82
R9380 vss.n21871 vss.n21870 11.793
R9381 vss.n3820 vss.n3819 11.793
R9382 vss.n12455 vss.n12451 11.702
R9383 vss.n12617 vss.n12613 11.702
R9384 vss.n14458 vss.n14454 11.702
R9385 vss.n14428 vss.n14424 11.702
R9386 vss.n14640 vss.n14636 11.702
R9387 vss.n13562 vss.n13558 11.702
R9388 vss.n15033 vss.n15029 11.702
R9389 vss.n10478 vss.n10474 11.702
R9390 vss.n13316 vss.n13312 11.702
R9391 vss.n14753 vss.n14749 11.702
R9392 vss.n14920 vss.n14916 11.702
R9393 vss.n14948 vss.n14944 11.702
R9394 vss.n14327 vss.n14323 11.702
R9395 vss.n13900 vss.n13896 11.702
R9396 vss.n14001 vss.n13997 11.702
R9397 vss.n11593 vss.n11589 11.702
R9398 vss.n11736 vss.n11732 11.702
R9399 vss.n11144 vss.n11140 11.702
R9400 vss.n10846 vss.n10842 11.702
R9401 vss.n10890 vss.n10886 11.702
R9402 vss.n11246 vss.n11242 11.702
R9403 vss.n11211 vss.n11207 11.702
R9404 vss.n12156 vss.n12152 11.702
R9405 vss.n12213 vss.n12209 11.702
R9406 vss.n22732 vss.n22729 11.588
R9407 vss.n22655 vss.n22652 11.588
R9408 vss.n22524 vss.n22521 11.588
R9409 vss.n22447 vss.n22444 11.588
R9410 vss.n22316 vss.n22313 11.588
R9411 vss.n22239 vss.n22236 11.588
R9412 vss.n22108 vss.n22105 11.588
R9413 vss.n17404 vss.n17401 11.588
R9414 vss.n21452 vss.n21449 11.588
R9415 vss.n21375 vss.n21372 11.588
R9416 vss.n21244 vss.n21241 11.588
R9417 vss.n21167 vss.n21164 11.588
R9418 vss.n21036 vss.n21033 11.588
R9419 vss.n20959 vss.n20956 11.588
R9420 vss.n12118 vss.n12116 11.588
R9421 vss.n12128 vss.n12126 11.588
R9422 vss.n10878 vss.n10876 11.588
R9423 vss.n11946 vss.n11944 11.588
R9424 vss.n14417 vss.n14415 11.588
R9425 vss.n14371 vss.n14369 11.588
R9426 vss.n11635 vss.n11633 11.588
R9427 vss.n11662 vss.n11660 11.588
R9428 vss.n13272 vss.n13270 11.588
R9429 vss.n13256 vss.n13254 11.588
R9430 vss.n13541 vss.n13539 11.588
R9431 vss.n14593 vss.n14591 11.588
R9432 vss.n14833 vss.n14831 11.588
R9433 vss.n14861 vss.n14859 11.588
R9434 vss.n10486 vss.n10484 11.588
R9435 vss.n10516 vss.n10514 11.588
R9436 vss.n8895 vss.n8892 11.588
R9437 vss.n8818 vss.n8815 11.588
R9438 vss.n8687 vss.n8684 11.588
R9439 vss.n8610 vss.n8607 11.588
R9440 vss.n8479 vss.n8476 11.588
R9441 vss.n8402 vss.n8399 11.588
R9442 vss.n8271 vss.n8268 11.588
R9443 vss.n8194 vss.n8191 11.588
R9444 vss.n8063 vss.n8060 11.588
R9445 vss.n7986 vss.n7983 11.588
R9446 vss.n7855 vss.n7852 11.588
R9447 vss.n7777 vss.n7774 11.588
R9448 vss.n7646 vss.n7643 11.588
R9449 vss.n7569 vss.n7566 11.588
R9450 vss.n12986 vss.n12985 10.727
R9451 vss.n12976 vss.n12975 10.727
R9452 vss.n12945 vss.n12944 10.727
R9453 vss.n13156 vss.n13155 10.727
R9454 vss.n13780 vss.n13779 10.727
R9455 vss.n13791 vss.n13790 10.727
R9456 vss.n11547 vss.n11546 10.727
R9457 vss.n11516 vss.n11515 10.727
R9458 vss.n14157 vss.n14156 10.727
R9459 vss.n14114 vss.n14113 10.727
R9460 vss.n13733 vss.n13732 10.727
R9461 vss.n11430 vss.n11429 10.727
R9462 vss.n11870 vss.n11869 10.727
R9463 vss.n11906 vss.n11905 10.727
R9464 vss.n12386 vss.n12385 10.727
R9465 vss.n12359 vss.n12358 10.727
R9466 vss.n10690 vss.n10689 10.727
R9467 vss.n10700 vss.n10699 10.727
R9468 vss.n13413 vss.n13412 10.727
R9469 vss.n13492 vss.n13491 10.727
R9470 vss.n13072 vss.n13071 10.727
R9471 vss.n10625 vss.n10624 10.727
R9472 vss.n10785 vss.n10784 10.727
R9473 vss.n12293 vss.n12292 10.727
R9474 vss.n21669 vss.n21666 10.264
R9475 vss.n3618 vss.n3615 10.264
R9476 vss.n8998 vss.n8997 10.093
R9477 vss.n20649 vss.n20644 9.879
R9478 vss.n20667 vss.n20662 9.879
R9479 vss.n7259 vss.n7254 9.879
R9480 vss.n7277 vss.n7272 9.879
R9481 vss.n1870 vss.n1865 9.879
R9482 vss.n1889 vss.n1883 9.879
R9483 vss.n2115 vss.n2109 9.879
R9484 vss.n2133 vss.n2127 9.879
R9485 vss.n2359 vss.n2353 9.879
R9486 vss.n2377 vss.n2371 9.879
R9487 vss.n2603 vss.n2597 9.879
R9488 vss.n2622 vss.n2616 9.879
R9489 vss.n2841 vss.n2836 9.879
R9490 vss.n2860 vss.n2854 9.879
R9491 vss.n3086 vss.n3080 9.879
R9492 vss.n3104 vss.n3098 9.879
R9493 vss.n3330 vss.n3324 9.879
R9494 vss.n3348 vss.n3343 9.879
R9495 vss.n331 vss.n326 9.879
R9496 vss.n350 vss.n344 9.879
R9497 vss.n576 vss.n570 9.879
R9498 vss.n594 vss.n588 9.879
R9499 vss.n820 vss.n814 9.879
R9500 vss.n838 vss.n832 9.879
R9501 vss.n1064 vss.n1058 9.879
R9502 vss.n1083 vss.n1077 9.879
R9503 vss.n1309 vss.n1303 9.879
R9504 vss.n23403 vss.n23397 9.879
R9505 vss.n23178 vss.n23172 9.879
R9506 vss.n23160 vss.n23154 9.879
R9507 vss.n22934 vss.n22928 9.879
R9508 vss.n22915 vss.n22910 9.879
R9509 vss.n17670 vss.n17664 9.85
R9510 vss.n18928 vss.n17697 9.85
R9511 vss.n18849 vss.n17768 9.85
R9512 vss.n18807 vss.n17807 9.85
R9513 vss.n18728 vss.n17878 9.85
R9514 vss.n18687 vss.n17910 9.85
R9515 vss.n18608 vss.n17981 9.85
R9516 vss.n18566 vss.n18020 9.85
R9517 vss.n18487 vss.n18091 9.85
R9518 vss.n18446 vss.n18123 9.85
R9519 vss.n18367 vss.n18194 9.85
R9520 vss.n18325 vss.n18233 9.85
R9521 vss.n20242 vss.n19068 9.85
R9522 vss.n20200 vss.n19107 9.85
R9523 vss.n19177 vss.n19171 9.85
R9524 vss.n20074 vss.n19204 9.85
R9525 vss.n19995 vss.n19275 9.85
R9526 vss.n19953 vss.n19314 9.85
R9527 vss.n19384 vss.n19378 9.85
R9528 vss.n19827 vss.n19411 9.85
R9529 vss.n19748 vss.n19482 9.85
R9530 vss.n19706 vss.n19521 9.85
R9531 vss.n19599 vss.n19585 9.85
R9532 vss.n4280 vss.n4274 9.85
R9533 vss.n5538 vss.n4307 9.85
R9534 vss.n5459 vss.n4378 9.85
R9535 vss.n5417 vss.n4417 9.85
R9536 vss.n5338 vss.n4488 9.85
R9537 vss.n5297 vss.n4520 9.85
R9538 vss.n5218 vss.n4591 9.85
R9539 vss.n5176 vss.n4630 9.85
R9540 vss.n5097 vss.n4701 9.85
R9541 vss.n5056 vss.n4733 9.85
R9542 vss.n4977 vss.n4804 9.85
R9543 vss.n4935 vss.n4843 9.85
R9544 vss.n6852 vss.n5678 9.85
R9545 vss.n6810 vss.n5717 9.85
R9546 vss.n5787 vss.n5781 9.85
R9547 vss.n6684 vss.n5814 9.85
R9548 vss.n6605 vss.n5885 9.85
R9549 vss.n6563 vss.n5924 9.85
R9550 vss.n5994 vss.n5988 9.85
R9551 vss.n6437 vss.n6021 9.85
R9552 vss.n6358 vss.n6092 9.85
R9553 vss.n6316 vss.n6131 9.85
R9554 vss.n6209 vss.n6195 9.85
R9555 vss.n16746 vss.n16745 9.85
R9556 vss.n16815 vss.n16814 9.85
R9557 vss.n16976 vss.n16975 9.85
R9558 vss.n17049 vss.n17048 9.85
R9559 vss.n17212 vss.n17211 9.85
R9560 vss.n17300 vss.n17299 9.85
R9561 vss.n16025 vss.n16022 9.85
R9562 vss.n16097 vss.n16094 9.85
R9563 vss.n15295 vss.n15294 9.85
R9564 vss.n15334 vss.n15333 9.85
R9565 vss.n15496 vss.n15495 9.85
R9566 vss.n15571 vss.n15570 9.85
R9567 vss.n15732 vss.n15731 9.85
R9568 vss.n15799 vss.n15798 9.85
R9569 vss.n16443 vss.n16442 9.85
R9570 vss.n16518 vss.n16517 9.85
R9571 vss.n9188 vss.n9181 9.777
R9572 vss.n22615 vss.n22611 9.656
R9573 vss.n22568 vss.n22564 9.656
R9574 vss.n22407 vss.n22403 9.656
R9575 vss.n22360 vss.n22356 9.656
R9576 vss.n22199 vss.n22195 9.656
R9577 vss.n22152 vss.n22148 9.656
R9578 vss.n21543 vss.n21539 9.656
R9579 vss.n21496 vss.n21492 9.656
R9580 vss.n21335 vss.n21331 9.656
R9581 vss.n21288 vss.n21284 9.656
R9582 vss.n21127 vss.n21123 9.656
R9583 vss.n21080 vss.n21076 9.656
R9584 vss.n20919 vss.n20915 9.656
R9585 vss.n8778 vss.n8774 9.656
R9586 vss.n8731 vss.n8727 9.656
R9587 vss.n8570 vss.n8566 9.656
R9588 vss.n8523 vss.n8519 9.656
R9589 vss.n8362 vss.n8358 9.656
R9590 vss.n8315 vss.n8311 9.656
R9591 vss.n8154 vss.n8150 9.656
R9592 vss.n8107 vss.n8103 9.656
R9593 vss.n7946 vss.n7942 9.656
R9594 vss.n7899 vss.n7895 9.656
R9595 vss.n7737 vss.n7733 9.656
R9596 vss.n7690 vss.n7686 9.656
R9597 vss.n7529 vss.n7525 9.656
R9598 vss.n16251 vss.n16249 9.527
R9599 vss.n16673 vss.n16672 9.527
R9600 vss.n8950 vss.n8949 9.33
R9601 vss.n3437 vss.n3436 9.319
R9602 vss.n1412 vss.n1411 9.319
R9603 vss.n21636 vss.n21609 9.307
R9604 vss.n3585 vss.n3558 9.307
R9605 vss.n19023 vss.n17630 9.3
R9606 vss.n19005 vss.n17640 9.3
R9607 vss.n17649 vss.n17648 9.3
R9608 vss.n17657 vss.n17647 9.3
R9609 vss.n18984 vss.n17656 9.3
R9610 vss.n18974 vss.n18973 9.3
R9611 vss.n17669 vss.n17666 9.3
R9612 vss.n18961 vss.n17676 9.3
R9613 vss.n18939 vss.n18938 9.3
R9614 vss.n18934 vss.n17692 9.3
R9615 vss.n18924 vss.n17704 9.3
R9616 vss.n17713 vss.n17711 9.3
R9617 vss.n18911 vss.n17714 9.3
R9618 vss.n18901 vss.n17723 9.3
R9619 vss.n17732 vss.n17730 9.3
R9620 vss.n18881 vss.n18880 9.3
R9621 vss.n17744 vss.n17742 9.3
R9622 vss.n18868 vss.n17754 9.3
R9623 vss.n18858 vss.n18857 9.3
R9624 vss.n17766 vss.n17763 9.3
R9625 vss.n18845 vss.n17773 9.3
R9626 vss.n18835 vss.n18834 9.3
R9627 vss.n18821 vss.n17795 9.3
R9628 vss.n18811 vss.n17804 9.3
R9629 vss.n17813 vss.n17811 9.3
R9630 vss.n18798 vss.n17814 9.3
R9631 vss.n18788 vss.n17823 9.3
R9632 vss.n17832 vss.n17830 9.3
R9633 vss.n18775 vss.n17833 9.3
R9634 vss.n17845 vss.n17843 9.3
R9635 vss.n18755 vss.n17854 9.3
R9636 vss.n18745 vss.n18744 9.3
R9637 vss.n17866 vss.n17863 9.3
R9638 vss.n18732 vss.n17873 9.3
R9639 vss.n18722 vss.n18721 9.3
R9640 vss.n17885 vss.n17882 9.3
R9641 vss.n18698 vss.n18697 9.3
R9642 vss.n18693 vss.n17905 9.3
R9643 vss.n18683 vss.n17917 9.3
R9644 vss.n17926 vss.n17924 9.3
R9645 vss.n18670 vss.n17927 9.3
R9646 vss.n18660 vss.n17936 9.3
R9647 vss.n17945 vss.n17943 9.3
R9648 vss.n18640 vss.n18639 9.3
R9649 vss.n17957 vss.n17955 9.3
R9650 vss.n18627 vss.n17967 9.3
R9651 vss.n18617 vss.n18616 9.3
R9652 vss.n17979 vss.n17976 9.3
R9653 vss.n18604 vss.n17986 9.3
R9654 vss.n18594 vss.n18593 9.3
R9655 vss.n18580 vss.n18008 9.3
R9656 vss.n18570 vss.n18017 9.3
R9657 vss.n18026 vss.n18024 9.3
R9658 vss.n18557 vss.n18027 9.3
R9659 vss.n18547 vss.n18036 9.3
R9660 vss.n18045 vss.n18043 9.3
R9661 vss.n18534 vss.n18046 9.3
R9662 vss.n18058 vss.n18056 9.3
R9663 vss.n18514 vss.n18067 9.3
R9664 vss.n18504 vss.n18503 9.3
R9665 vss.n18079 vss.n18076 9.3
R9666 vss.n18491 vss.n18086 9.3
R9667 vss.n18481 vss.n18480 9.3
R9668 vss.n18098 vss.n18095 9.3
R9669 vss.n18457 vss.n18456 9.3
R9670 vss.n18452 vss.n18118 9.3
R9671 vss.n18442 vss.n18130 9.3
R9672 vss.n18139 vss.n18137 9.3
R9673 vss.n18429 vss.n18140 9.3
R9674 vss.n18419 vss.n18149 9.3
R9675 vss.n18158 vss.n18156 9.3
R9676 vss.n18399 vss.n18398 9.3
R9677 vss.n18170 vss.n18168 9.3
R9678 vss.n18386 vss.n18180 9.3
R9679 vss.n18376 vss.n18375 9.3
R9680 vss.n18192 vss.n18189 9.3
R9681 vss.n18363 vss.n18199 9.3
R9682 vss.n18353 vss.n18352 9.3
R9683 vss.n18339 vss.n18221 9.3
R9684 vss.n18329 vss.n18230 9.3
R9685 vss.n18239 vss.n18237 9.3
R9686 vss.n18316 vss.n18240 9.3
R9687 vss.n18306 vss.n18249 9.3
R9688 vss.n18258 vss.n18256 9.3
R9689 vss.n18293 vss.n18259 9.3
R9690 vss.n18297 vss.n18296 9.3
R9691 vss.n18298 vss.n18297 9.3
R9692 vss.n18299 vss.n18298 9.3
R9693 vss.n18255 vss.n18250 9.3
R9694 vss.n18315 vss.n18243 9.3
R9695 vss.n18315 vss.n18314 9.3
R9696 vss.n18314 vss.n18313 9.3
R9697 vss.n18318 vss.n18317 9.3
R9698 vss.n18328 vss.n18327 9.3
R9699 vss.n18327 vss.n18229 9.3
R9700 vss.n18229 vss.n18228 9.3
R9701 vss.n18331 vss.n18330 9.3
R9702 vss.n18343 vss.n18342 9.3
R9703 vss.n18344 vss.n18343 9.3
R9704 vss.n18345 vss.n18344 9.3
R9705 vss.n18351 vss.n18207 9.3
R9706 vss.n18201 vss.n18200 9.3
R9707 vss.n18385 vss.n18384 9.3
R9708 vss.n18397 vss.n18167 9.3
R9709 vss.n18418 vss.n18417 9.3
R9710 vss.n18417 vss.n18148 9.3
R9711 vss.n18148 vss.n18147 9.3
R9712 vss.n18421 vss.n18420 9.3
R9713 vss.n18433 vss.n18432 9.3
R9714 vss.n18434 vss.n18433 9.3
R9715 vss.n18435 vss.n18434 9.3
R9716 vss.n18136 vss.n18131 9.3
R9717 vss.n18451 vss.n18121 9.3
R9718 vss.n18451 vss.n18450 9.3
R9719 vss.n18450 vss.n18449 9.3
R9720 vss.n18454 vss.n18453 9.3
R9721 vss.n18466 vss.n18465 9.3
R9722 vss.n18465 vss.n18464 9.3
R9723 vss.n18464 vss.n18463 9.3
R9724 vss.n18107 vss.n18106 9.3
R9725 vss.n18490 vss.n18489 9.3
R9726 vss.n18502 vss.n18075 9.3
R9727 vss.n18069 vss.n18068 9.3
R9728 vss.n18538 vss.n18537 9.3
R9729 vss.n18539 vss.n18538 9.3
R9730 vss.n18540 vss.n18539 9.3
R9731 vss.n18042 vss.n18037 9.3
R9732 vss.n18556 vss.n18030 9.3
R9733 vss.n18556 vss.n18555 9.3
R9734 vss.n18555 vss.n18554 9.3
R9735 vss.n18559 vss.n18558 9.3
R9736 vss.n18569 vss.n18568 9.3
R9737 vss.n18568 vss.n18016 9.3
R9738 vss.n18016 vss.n18015 9.3
R9739 vss.n18572 vss.n18571 9.3
R9740 vss.n18584 vss.n18583 9.3
R9741 vss.n18585 vss.n18584 9.3
R9742 vss.n18586 vss.n18585 9.3
R9743 vss.n18592 vss.n17994 9.3
R9744 vss.n17988 vss.n17987 9.3
R9745 vss.n18626 vss.n18625 9.3
R9746 vss.n18638 vss.n17954 9.3
R9747 vss.n18659 vss.n18658 9.3
R9748 vss.n18658 vss.n17935 9.3
R9749 vss.n17935 vss.n17934 9.3
R9750 vss.n18662 vss.n18661 9.3
R9751 vss.n18674 vss.n18673 9.3
R9752 vss.n18675 vss.n18674 9.3
R9753 vss.n18676 vss.n18675 9.3
R9754 vss.n17923 vss.n17918 9.3
R9755 vss.n18692 vss.n17908 9.3
R9756 vss.n18692 vss.n18691 9.3
R9757 vss.n18691 vss.n18690 9.3
R9758 vss.n18695 vss.n18694 9.3
R9759 vss.n18707 vss.n18706 9.3
R9760 vss.n18706 vss.n18705 9.3
R9761 vss.n18705 vss.n18704 9.3
R9762 vss.n17894 vss.n17893 9.3
R9763 vss.n18731 vss.n18730 9.3
R9764 vss.n18743 vss.n17862 9.3
R9765 vss.n17856 vss.n17855 9.3
R9766 vss.n18779 vss.n18778 9.3
R9767 vss.n18780 vss.n18779 9.3
R9768 vss.n18781 vss.n18780 9.3
R9769 vss.n17829 vss.n17824 9.3
R9770 vss.n18797 vss.n17817 9.3
R9771 vss.n18797 vss.n18796 9.3
R9772 vss.n18796 vss.n18795 9.3
R9773 vss.n18800 vss.n18799 9.3
R9774 vss.n18810 vss.n18809 9.3
R9775 vss.n18809 vss.n17803 9.3
R9776 vss.n17803 vss.n17802 9.3
R9777 vss.n18813 vss.n18812 9.3
R9778 vss.n18825 vss.n18824 9.3
R9779 vss.n18826 vss.n18825 9.3
R9780 vss.n18827 vss.n18826 9.3
R9781 vss.n18833 vss.n17781 9.3
R9782 vss.n17775 vss.n17774 9.3
R9783 vss.n18867 vss.n18866 9.3
R9784 vss.n18879 vss.n17741 9.3
R9785 vss.n18900 vss.n18899 9.3
R9786 vss.n18899 vss.n17722 9.3
R9787 vss.n17722 vss.n17721 9.3
R9788 vss.n18903 vss.n18902 9.3
R9789 vss.n18915 vss.n18914 9.3
R9790 vss.n18916 vss.n18915 9.3
R9791 vss.n18917 vss.n18916 9.3
R9792 vss.n17710 vss.n17705 9.3
R9793 vss.n18933 vss.n17695 9.3
R9794 vss.n18933 vss.n18932 9.3
R9795 vss.n18932 vss.n18931 9.3
R9796 vss.n18936 vss.n18935 9.3
R9797 vss.n18948 vss.n18947 9.3
R9798 vss.n18947 vss.n18946 9.3
R9799 vss.n18946 vss.n18945 9.3
R9800 vss.n18960 vss.n18959 9.3
R9801 vss.n18972 vss.n17665 9.3
R9802 vss.n17659 vss.n17658 9.3
R9803 vss.n19004 vss.n19003 9.3
R9804 vss.n17629 vss.n17626 9.3
R9805 vss.n19025 vss.n19024 9.3
R9806 vss.n19022 vss.n19021 9.3
R9807 vss.n19021 vss.n19020 9.3
R9808 vss.n19020 vss.n19019 9.3
R9809 vss.n19007 vss.n19006 9.3
R9810 vss.n19008 vss.n19007 9.3
R9811 vss.n19009 vss.n19008 9.3
R9812 vss.n17642 vss.n17641 9.3
R9813 vss.n17643 vss.n17642 9.3
R9814 vss.n18998 vss.n17643 9.3
R9815 vss.n17650 vss.n17646 9.3
R9816 vss.n18993 vss.n17651 9.3
R9817 vss.n18993 vss.n18992 9.3
R9818 vss.n18992 vss.n18991 9.3
R9819 vss.n18986 vss.n18985 9.3
R9820 vss.n18986 vss.n17654 9.3
R9821 vss.n17654 vss.n17653 9.3
R9822 vss.n18983 vss.n18982 9.3
R9823 vss.n18975 vss.n17660 9.3
R9824 vss.n18976 vss.n18975 9.3
R9825 vss.n18977 vss.n18976 9.3
R9826 vss.n18971 vss.n18970 9.3
R9827 vss.n18970 vss.n18969 9.3
R9828 vss.n18969 vss.n18968 9.3
R9829 vss.n17678 vss.n17677 9.3
R9830 vss.n18963 vss.n18962 9.3
R9831 vss.n18963 vss.n17674 9.3
R9832 vss.n17674 vss.n17673 9.3
R9833 vss.n18952 vss.n17679 9.3
R9834 vss.n18953 vss.n18952 9.3
R9835 vss.n18954 vss.n18953 9.3
R9836 vss.n18940 vss.n17686 9.3
R9837 vss.n18937 vss.n17691 9.3
R9838 vss.n17691 vss.n17690 9.3
R9839 vss.n17690 vss.n17689 9.3
R9840 vss.n18926 vss.n18925 9.3
R9841 vss.n18923 vss.n18922 9.3
R9842 vss.n18922 vss.n17703 9.3
R9843 vss.n17703 vss.n17702 9.3
R9844 vss.n18913 vss.n18912 9.3
R9845 vss.n18910 vss.n17717 9.3
R9846 vss.n18910 vss.n18909 9.3
R9847 vss.n18909 vss.n18908 9.3
R9848 vss.n17729 vss.n17724 9.3
R9849 vss.n18892 vss.n18891 9.3
R9850 vss.n18893 vss.n18892 9.3
R9851 vss.n18894 vss.n18893 9.3
R9852 vss.n18882 vss.n17733 9.3
R9853 vss.n18882 vss.n17740 9.3
R9854 vss.n17740 vss.n17739 9.3
R9855 vss.n18878 vss.n18877 9.3
R9856 vss.n18877 vss.n18876 9.3
R9857 vss.n18876 vss.n18875 9.3
R9858 vss.n17756 vss.n17755 9.3
R9859 vss.n18870 vss.n18869 9.3
R9860 vss.n18870 vss.n17752 9.3
R9861 vss.n17752 vss.n17751 9.3
R9862 vss.n18859 vss.n17757 9.3
R9863 vss.n18860 vss.n18859 9.3
R9864 vss.n18861 vss.n18860 9.3
R9865 vss.n18856 vss.n17762 9.3
R9866 vss.n18855 vss.n18854 9.3
R9867 vss.n18854 vss.n18853 9.3
R9868 vss.n18853 vss.n18852 9.3
R9869 vss.n18847 vss.n18846 9.3
R9870 vss.n18847 vss.n17771 9.3
R9871 vss.n17771 vss.n17770 9.3
R9872 vss.n18844 vss.n18843 9.3
R9873 vss.n18836 vss.n17776 9.3
R9874 vss.n18837 vss.n18836 9.3
R9875 vss.n18838 vss.n18837 9.3
R9876 vss.n18832 vss.n18831 9.3
R9877 vss.n18831 vss.n18830 9.3
R9878 vss.n18830 vss.n18829 9.3
R9879 vss.n18823 vss.n18822 9.3
R9880 vss.n18820 vss.n17798 9.3
R9881 vss.n18820 vss.n18819 9.3
R9882 vss.n18819 vss.n18818 9.3
R9883 vss.n17810 vss.n17805 9.3
R9884 vss.n18802 vss.n18801 9.3
R9885 vss.n18803 vss.n18802 9.3
R9886 vss.n18804 vss.n18803 9.3
R9887 vss.n18790 vss.n18789 9.3
R9888 vss.n18787 vss.n18786 9.3
R9889 vss.n18786 vss.n17822 9.3
R9890 vss.n17822 vss.n17821 9.3
R9891 vss.n18777 vss.n18776 9.3
R9892 vss.n18774 vss.n17836 9.3
R9893 vss.n18774 vss.n18773 9.3
R9894 vss.n18773 vss.n18772 9.3
R9895 vss.n18765 vss.n18764 9.3
R9896 vss.n18764 vss.n18763 9.3
R9897 vss.n18763 vss.n18762 9.3
R9898 vss.n18757 vss.n18756 9.3
R9899 vss.n18757 vss.n17852 9.3
R9900 vss.n17852 vss.n17851 9.3
R9901 vss.n18754 vss.n18753 9.3
R9902 vss.n18746 vss.n17857 9.3
R9903 vss.n18747 vss.n18746 9.3
R9904 vss.n18748 vss.n18747 9.3
R9905 vss.n18742 vss.n18741 9.3
R9906 vss.n18741 vss.n18740 9.3
R9907 vss.n18740 vss.n18739 9.3
R9908 vss.n17875 vss.n17874 9.3
R9909 vss.n18734 vss.n18733 9.3
R9910 vss.n18734 vss.n17871 9.3
R9911 vss.n17871 vss.n17870 9.3
R9912 vss.n18723 vss.n17876 9.3
R9913 vss.n18724 vss.n18723 9.3
R9914 vss.n18725 vss.n18724 9.3
R9915 vss.n18720 vss.n17881 9.3
R9916 vss.n18719 vss.n18718 9.3
R9917 vss.n18718 vss.n18717 9.3
R9918 vss.n18717 vss.n18716 9.3
R9919 vss.n18711 vss.n18710 9.3
R9920 vss.n18711 vss.n17890 9.3
R9921 vss.n17890 vss.n17889 9.3
R9922 vss.n18699 vss.n17896 9.3
R9923 vss.n18696 vss.n17904 9.3
R9924 vss.n17904 vss.n17903 9.3
R9925 vss.n17903 vss.n17902 9.3
R9926 vss.n18685 vss.n18684 9.3
R9927 vss.n18682 vss.n18681 9.3
R9928 vss.n18681 vss.n17916 9.3
R9929 vss.n17916 vss.n17915 9.3
R9930 vss.n18672 vss.n18671 9.3
R9931 vss.n18669 vss.n17930 9.3
R9932 vss.n18669 vss.n18668 9.3
R9933 vss.n18668 vss.n18667 9.3
R9934 vss.n17942 vss.n17937 9.3
R9935 vss.n18651 vss.n18650 9.3
R9936 vss.n18652 vss.n18651 9.3
R9937 vss.n18653 vss.n18652 9.3
R9938 vss.n18641 vss.n17946 9.3
R9939 vss.n18641 vss.n17953 9.3
R9940 vss.n17953 vss.n17952 9.3
R9941 vss.n18637 vss.n18636 9.3
R9942 vss.n18636 vss.n18635 9.3
R9943 vss.n18635 vss.n18634 9.3
R9944 vss.n17969 vss.n17968 9.3
R9945 vss.n18629 vss.n18628 9.3
R9946 vss.n18629 vss.n17965 9.3
R9947 vss.n17965 vss.n17964 9.3
R9948 vss.n18618 vss.n17970 9.3
R9949 vss.n18619 vss.n18618 9.3
R9950 vss.n18620 vss.n18619 9.3
R9951 vss.n18615 vss.n17975 9.3
R9952 vss.n18614 vss.n18613 9.3
R9953 vss.n18613 vss.n18612 9.3
R9954 vss.n18612 vss.n18611 9.3
R9955 vss.n18606 vss.n18605 9.3
R9956 vss.n18606 vss.n17984 9.3
R9957 vss.n17984 vss.n17983 9.3
R9958 vss.n18603 vss.n18602 9.3
R9959 vss.n18595 vss.n17989 9.3
R9960 vss.n18596 vss.n18595 9.3
R9961 vss.n18597 vss.n18596 9.3
R9962 vss.n18591 vss.n18590 9.3
R9963 vss.n18590 vss.n18589 9.3
R9964 vss.n18589 vss.n18588 9.3
R9965 vss.n18582 vss.n18581 9.3
R9966 vss.n18579 vss.n18011 9.3
R9967 vss.n18579 vss.n18578 9.3
R9968 vss.n18578 vss.n18577 9.3
R9969 vss.n18023 vss.n18018 9.3
R9970 vss.n18561 vss.n18560 9.3
R9971 vss.n18562 vss.n18561 9.3
R9972 vss.n18563 vss.n18562 9.3
R9973 vss.n18549 vss.n18548 9.3
R9974 vss.n18546 vss.n18545 9.3
R9975 vss.n18545 vss.n18035 9.3
R9976 vss.n18035 vss.n18034 9.3
R9977 vss.n18536 vss.n18535 9.3
R9978 vss.n18533 vss.n18049 9.3
R9979 vss.n18533 vss.n18532 9.3
R9980 vss.n18532 vss.n18531 9.3
R9981 vss.n18524 vss.n18523 9.3
R9982 vss.n18523 vss.n18522 9.3
R9983 vss.n18522 vss.n18521 9.3
R9984 vss.n18516 vss.n18515 9.3
R9985 vss.n18516 vss.n18065 9.3
R9986 vss.n18065 vss.n18064 9.3
R9987 vss.n18513 vss.n18512 9.3
R9988 vss.n18505 vss.n18070 9.3
R9989 vss.n18506 vss.n18505 9.3
R9990 vss.n18507 vss.n18506 9.3
R9991 vss.n18501 vss.n18500 9.3
R9992 vss.n18500 vss.n18499 9.3
R9993 vss.n18499 vss.n18498 9.3
R9994 vss.n18088 vss.n18087 9.3
R9995 vss.n18493 vss.n18492 9.3
R9996 vss.n18493 vss.n18084 9.3
R9997 vss.n18084 vss.n18083 9.3
R9998 vss.n18482 vss.n18089 9.3
R9999 vss.n18483 vss.n18482 9.3
R10000 vss.n18484 vss.n18483 9.3
R10001 vss.n18479 vss.n18094 9.3
R10002 vss.n18478 vss.n18477 9.3
R10003 vss.n18477 vss.n18476 9.3
R10004 vss.n18476 vss.n18475 9.3
R10005 vss.n18470 vss.n18469 9.3
R10006 vss.n18470 vss.n18103 9.3
R10007 vss.n18103 vss.n18102 9.3
R10008 vss.n18458 vss.n18109 9.3
R10009 vss.n18455 vss.n18117 9.3
R10010 vss.n18117 vss.n18116 9.3
R10011 vss.n18116 vss.n18115 9.3
R10012 vss.n18444 vss.n18443 9.3
R10013 vss.n18441 vss.n18440 9.3
R10014 vss.n18440 vss.n18129 9.3
R10015 vss.n18129 vss.n18128 9.3
R10016 vss.n18431 vss.n18430 9.3
R10017 vss.n18428 vss.n18143 9.3
R10018 vss.n18428 vss.n18427 9.3
R10019 vss.n18427 vss.n18426 9.3
R10020 vss.n18155 vss.n18150 9.3
R10021 vss.n18410 vss.n18409 9.3
R10022 vss.n18411 vss.n18410 9.3
R10023 vss.n18412 vss.n18411 9.3
R10024 vss.n18400 vss.n18159 9.3
R10025 vss.n18400 vss.n18166 9.3
R10026 vss.n18166 vss.n18165 9.3
R10027 vss.n18396 vss.n18395 9.3
R10028 vss.n18395 vss.n18394 9.3
R10029 vss.n18394 vss.n18393 9.3
R10030 vss.n18182 vss.n18181 9.3
R10031 vss.n18388 vss.n18387 9.3
R10032 vss.n18388 vss.n18178 9.3
R10033 vss.n18178 vss.n18177 9.3
R10034 vss.n18377 vss.n18183 9.3
R10035 vss.n18378 vss.n18377 9.3
R10036 vss.n18379 vss.n18378 9.3
R10037 vss.n18374 vss.n18188 9.3
R10038 vss.n18373 vss.n18372 9.3
R10039 vss.n18372 vss.n18371 9.3
R10040 vss.n18371 vss.n18370 9.3
R10041 vss.n18365 vss.n18364 9.3
R10042 vss.n18365 vss.n18197 9.3
R10043 vss.n18197 vss.n18196 9.3
R10044 vss.n18362 vss.n18361 9.3
R10045 vss.n18354 vss.n18202 9.3
R10046 vss.n18355 vss.n18354 9.3
R10047 vss.n18356 vss.n18355 9.3
R10048 vss.n18350 vss.n18349 9.3
R10049 vss.n18349 vss.n18348 9.3
R10050 vss.n18348 vss.n18347 9.3
R10051 vss.n18341 vss.n18340 9.3
R10052 vss.n18338 vss.n18224 9.3
R10053 vss.n18338 vss.n18337 9.3
R10054 vss.n18337 vss.n18336 9.3
R10055 vss.n18236 vss.n18231 9.3
R10056 vss.n18320 vss.n18319 9.3
R10057 vss.n18321 vss.n18320 9.3
R10058 vss.n18322 vss.n18321 9.3
R10059 vss.n18308 vss.n18307 9.3
R10060 vss.n18305 vss.n18304 9.3
R10061 vss.n18304 vss.n18248 9.3
R10062 vss.n18248 vss.n18247 9.3
R10063 vss.n18295 vss.n18294 9.3
R10064 vss.n18292 vss.n18262 9.3
R10065 vss.n18292 vss.n18291 9.3
R10066 vss.n18291 vss.n18290 9.3
R10067 vss.n18271 vss.n18269 9.3
R10068 vss.n18273 vss.n17623 9.3
R10069 vss.n18283 vss.n18282 9.3
R10070 vss.n18282 vss.n18281 9.3
R10071 vss.n18281 vss.n18280 9.3
R10072 vss.n19030 vss.n2 9.3
R10073 vss.n17591 vss.n17586 9.3
R10074 vss.n20367 vss.n20366 9.3
R10075 vss.n17590 vss.n17589 9.3
R10076 vss.n20368 vss.n17581 9.3
R10077 vss.n19594 vss.n19593 9.3
R10078 vss.n19604 vss.n19592 9.3
R10079 vss.n20289 vss.n17622 9.3
R10080 vss.n19046 vss.n19045 9.3
R10081 vss.n19054 vss.n19043 9.3
R10082 vss.n20261 vss.n19053 9.3
R10083 vss.n20251 vss.n20250 9.3
R10084 vss.n19066 vss.n19063 9.3
R10085 vss.n20238 vss.n19073 9.3
R10086 vss.n20228 vss.n20227 9.3
R10087 vss.n20214 vss.n19095 9.3
R10088 vss.n20204 vss.n19104 9.3
R10089 vss.n19113 vss.n19111 9.3
R10090 vss.n20191 vss.n19114 9.3
R10091 vss.n20181 vss.n19123 9.3
R10092 vss.n19132 vss.n19130 9.3
R10093 vss.n20168 vss.n19133 9.3
R10094 vss.n20151 vss.n19147 9.3
R10095 vss.n19156 vss.n19155 9.3
R10096 vss.n19164 vss.n19154 9.3
R10097 vss.n20130 vss.n19163 9.3
R10098 vss.n20120 vss.n20119 9.3
R10099 vss.n19176 vss.n19173 9.3
R10100 vss.n20107 vss.n19183 9.3
R10101 vss.n20085 vss.n20084 9.3
R10102 vss.n20080 vss.n19199 9.3
R10103 vss.n20070 vss.n19211 9.3
R10104 vss.n19220 vss.n19218 9.3
R10105 vss.n20057 vss.n19221 9.3
R10106 vss.n20047 vss.n19230 9.3
R10107 vss.n19239 vss.n19237 9.3
R10108 vss.n20027 vss.n20026 9.3
R10109 vss.n19251 vss.n19249 9.3
R10110 vss.n20014 vss.n19261 9.3
R10111 vss.n20004 vss.n20003 9.3
R10112 vss.n19273 vss.n19270 9.3
R10113 vss.n19991 vss.n19280 9.3
R10114 vss.n19981 vss.n19980 9.3
R10115 vss.n19967 vss.n19302 9.3
R10116 vss.n19957 vss.n19311 9.3
R10117 vss.n19320 vss.n19318 9.3
R10118 vss.n19944 vss.n19321 9.3
R10119 vss.n19934 vss.n19330 9.3
R10120 vss.n19339 vss.n19337 9.3
R10121 vss.n19921 vss.n19340 9.3
R10122 vss.n19904 vss.n19354 9.3
R10123 vss.n19363 vss.n19362 9.3
R10124 vss.n19371 vss.n19361 9.3
R10125 vss.n19883 vss.n19370 9.3
R10126 vss.n19873 vss.n19872 9.3
R10127 vss.n19383 vss.n19380 9.3
R10128 vss.n19860 vss.n19390 9.3
R10129 vss.n19838 vss.n19837 9.3
R10130 vss.n19833 vss.n19406 9.3
R10131 vss.n19823 vss.n19418 9.3
R10132 vss.n19427 vss.n19425 9.3
R10133 vss.n19810 vss.n19428 9.3
R10134 vss.n19800 vss.n19437 9.3
R10135 vss.n19446 vss.n19444 9.3
R10136 vss.n19780 vss.n19779 9.3
R10137 vss.n19458 vss.n19456 9.3
R10138 vss.n19767 vss.n19468 9.3
R10139 vss.n19757 vss.n19756 9.3
R10140 vss.n19480 vss.n19477 9.3
R10141 vss.n19744 vss.n19487 9.3
R10142 vss.n19734 vss.n19733 9.3
R10143 vss.n19720 vss.n19509 9.3
R10144 vss.n19710 vss.n19518 9.3
R10145 vss.n19527 vss.n19525 9.3
R10146 vss.n19697 vss.n19528 9.3
R10147 vss.n19687 vss.n19537 9.3
R10148 vss.n19546 vss.n19544 9.3
R10149 vss.n19674 vss.n19547 9.3
R10150 vss.n19657 vss.n19561 9.3
R10151 vss.n19570 vss.n19569 9.3
R10152 vss.n19578 vss.n19568 9.3
R10153 vss.n19636 vss.n19577 9.3
R10154 vss.n19626 vss.n19625 9.3
R10155 vss.n19635 vss.n19634 9.3
R10156 vss.n19571 vss.n19567 9.3
R10157 vss.n19676 vss.n19675 9.3
R10158 vss.n19689 vss.n19688 9.3
R10159 vss.n19524 vss.n19519 9.3
R10160 vss.n19722 vss.n19721 9.3
R10161 vss.n19743 vss.n19742 9.3
R10162 vss.n19755 vss.n19476 9.3
R10163 vss.n19470 vss.n19469 9.3
R10164 vss.n19443 vss.n19438 9.3
R10165 vss.n19812 vss.n19811 9.3
R10166 vss.n19825 vss.n19824 9.3
R10167 vss.n19839 vss.n19399 9.3
R10168 vss.n19392 vss.n19391 9.3
R10169 vss.n19882 vss.n19881 9.3
R10170 vss.n19364 vss.n19360 9.3
R10171 vss.n19923 vss.n19922 9.3
R10172 vss.n19936 vss.n19935 9.3
R10173 vss.n19317 vss.n19312 9.3
R10174 vss.n19969 vss.n19968 9.3
R10175 vss.n19990 vss.n19989 9.3
R10176 vss.n20002 vss.n19269 9.3
R10177 vss.n19263 vss.n19262 9.3
R10178 vss.n19236 vss.n19231 9.3
R10179 vss.n20059 vss.n20058 9.3
R10180 vss.n20072 vss.n20071 9.3
R10181 vss.n20086 vss.n19193 9.3
R10182 vss.n19185 vss.n19184 9.3
R10183 vss.n20129 vss.n20128 9.3
R10184 vss.n19157 vss.n19153 9.3
R10185 vss.n20170 vss.n20169 9.3
R10186 vss.n20183 vss.n20182 9.3
R10187 vss.n19110 vss.n19105 9.3
R10188 vss.n20216 vss.n20215 9.3
R10189 vss.n20237 vss.n20236 9.3
R10190 vss.n20249 vss.n19062 9.3
R10191 vss.n19056 vss.n19055 9.3
R10192 vss.n20291 vss.n20290 9.3
R10193 vss.n19047 vss.n19042 9.3
R10194 vss.n20260 vss.n20259 9.3
R10195 vss.n19075 vss.n19074 9.3
R10196 vss.n20226 vss.n19081 9.3
R10197 vss.n20206 vss.n20205 9.3
R10198 vss.n20193 vss.n20192 9.3
R10199 vss.n19129 vss.n19124 9.3
R10200 vss.n20150 vss.n20149 9.3
R10201 vss.n19166 vss.n19165 9.3
R10202 vss.n20118 vss.n19172 9.3
R10203 vss.n20106 vss.n20105 9.3
R10204 vss.n20082 vss.n20081 9.3
R10205 vss.n19217 vss.n19212 9.3
R10206 vss.n20049 vss.n20048 9.3
R10207 vss.n20025 vss.n19248 9.3
R10208 vss.n20013 vss.n20012 9.3
R10209 vss.n19282 vss.n19281 9.3
R10210 vss.n19979 vss.n19288 9.3
R10211 vss.n19959 vss.n19958 9.3
R10212 vss.n19946 vss.n19945 9.3
R10213 vss.n19336 vss.n19331 9.3
R10214 vss.n19903 vss.n19902 9.3
R10215 vss.n19373 vss.n19372 9.3
R10216 vss.n19871 vss.n19379 9.3
R10217 vss.n19859 vss.n19858 9.3
R10218 vss.n19835 vss.n19834 9.3
R10219 vss.n19424 vss.n19419 9.3
R10220 vss.n19802 vss.n19801 9.3
R10221 vss.n19778 vss.n19455 9.3
R10222 vss.n19766 vss.n19765 9.3
R10223 vss.n19489 vss.n19488 9.3
R10224 vss.n19732 vss.n19495 9.3
R10225 vss.n19712 vss.n19711 9.3
R10226 vss.n19699 vss.n19698 9.3
R10227 vss.n19543 vss.n19538 9.3
R10228 vss.n19656 vss.n19655 9.3
R10229 vss.n19580 vss.n19579 9.3
R10230 vss.n19624 vss.n19586 9.3
R10231 vss.n20322 vss.n17605 9.3
R10232 vss.n20327 vss.n20326 9.3
R10233 vss.n20332 vss.n17601 9.3
R10234 vss.n20359 vss.n20358 9.3
R10235 vss.n20358 vss.n20357 9.3
R10236 vss.n20357 vss.n20356 9.3
R10237 vss.n20354 vss.n20353 9.3
R10238 vss.n20348 vss.n17596 9.3
R10239 vss.n20343 vss.n20342 9.3
R10240 vss.n20337 vss.n17599 9.3
R10241 vss.n17613 vss.n17607 9.3
R10242 vss.n20301 vss.n20300 9.3
R10243 vss.n19673 vss.n19550 9.3
R10244 vss.n19673 vss.n19672 9.3
R10245 vss.n19672 vss.n19671 9.3
R10246 vss.n19686 vss.n19685 9.3
R10247 vss.n19685 vss.n19536 9.3
R10248 vss.n19536 vss.n19535 9.3
R10249 vss.n19701 vss.n19700 9.3
R10250 vss.n19702 vss.n19701 9.3
R10251 vss.n19703 vss.n19702 9.3
R10252 vss.n19719 vss.n19512 9.3
R10253 vss.n19719 vss.n19718 9.3
R10254 vss.n19718 vss.n19717 9.3
R10255 vss.n19791 vss.n19790 9.3
R10256 vss.n19792 vss.n19791 9.3
R10257 vss.n19793 vss.n19792 9.3
R10258 vss.n19809 vss.n19431 9.3
R10259 vss.n19809 vss.n19808 9.3
R10260 vss.n19808 vss.n19807 9.3
R10261 vss.n19822 vss.n19821 9.3
R10262 vss.n19821 vss.n19417 9.3
R10263 vss.n19417 vss.n19416 9.3
R10264 vss.n19836 vss.n19405 9.3
R10265 vss.n19405 vss.n19404 9.3
R10266 vss.n19404 vss.n19403 9.3
R10267 vss.n19920 vss.n19343 9.3
R10268 vss.n19920 vss.n19919 9.3
R10269 vss.n19919 vss.n19918 9.3
R10270 vss.n19933 vss.n19932 9.3
R10271 vss.n19932 vss.n19329 9.3
R10272 vss.n19329 vss.n19328 9.3
R10273 vss.n19948 vss.n19947 9.3
R10274 vss.n19949 vss.n19948 9.3
R10275 vss.n19950 vss.n19949 9.3
R10276 vss.n19966 vss.n19305 9.3
R10277 vss.n19966 vss.n19965 9.3
R10278 vss.n19965 vss.n19964 9.3
R10279 vss.n20038 vss.n20037 9.3
R10280 vss.n20039 vss.n20038 9.3
R10281 vss.n20040 vss.n20039 9.3
R10282 vss.n20056 vss.n19224 9.3
R10283 vss.n20056 vss.n20055 9.3
R10284 vss.n20055 vss.n20054 9.3
R10285 vss.n20069 vss.n20068 9.3
R10286 vss.n20068 vss.n19210 9.3
R10287 vss.n19210 vss.n19209 9.3
R10288 vss.n20083 vss.n19198 9.3
R10289 vss.n19198 vss.n19197 9.3
R10290 vss.n19197 vss.n19196 9.3
R10291 vss.n20167 vss.n19136 9.3
R10292 vss.n20167 vss.n20166 9.3
R10293 vss.n20166 vss.n20165 9.3
R10294 vss.n20180 vss.n20179 9.3
R10295 vss.n20179 vss.n19122 9.3
R10296 vss.n19122 vss.n19121 9.3
R10297 vss.n20195 vss.n20194 9.3
R10298 vss.n20196 vss.n20195 9.3
R10299 vss.n20197 vss.n20196 9.3
R10300 vss.n20213 vss.n19098 9.3
R10301 vss.n20213 vss.n20212 9.3
R10302 vss.n20212 vss.n20211 9.3
R10303 vss.n20288 vss.n20287 9.3
R10304 vss.n20287 vss.n17620 9.3
R10305 vss.n17620 vss.n17619 9.3
R10306 vss.n0 vss.n17618 9.3
R10307 vss.n19044 vss.n19038 9.3
R10308 vss.n19039 vss.n19038 9.3
R10309 vss.n20275 vss.n19039 9.3
R10310 vss.n20270 vss.n19048 9.3
R10311 vss.n20270 vss.n20269 9.3
R10312 vss.n20269 vss.n20268 9.3
R10313 vss.n20263 vss.n20262 9.3
R10314 vss.n20263 vss.n19051 9.3
R10315 vss.n19051 vss.n19050 9.3
R10316 vss.n20252 vss.n19057 9.3
R10317 vss.n20253 vss.n20252 9.3
R10318 vss.n20254 vss.n20253 9.3
R10319 vss.n20248 vss.n20247 9.3
R10320 vss.n20247 vss.n20246 9.3
R10321 vss.n20246 vss.n20245 9.3
R10322 vss.n20240 vss.n20239 9.3
R10323 vss.n20240 vss.n19071 9.3
R10324 vss.n19071 vss.n19070 9.3
R10325 vss.n20229 vss.n19076 9.3
R10326 vss.n20230 vss.n20229 9.3
R10327 vss.n20231 vss.n20230 9.3
R10328 vss.n20225 vss.n20224 9.3
R10329 vss.n20224 vss.n20223 9.3
R10330 vss.n20223 vss.n20222 9.3
R10331 vss.n20218 vss.n20217 9.3
R10332 vss.n20219 vss.n20218 9.3
R10333 vss.n20220 vss.n20219 9.3
R10334 vss.n20203 vss.n20202 9.3
R10335 vss.n20202 vss.n19103 9.3
R10336 vss.n19103 vss.n19102 9.3
R10337 vss.n20190 vss.n19117 9.3
R10338 vss.n20190 vss.n20189 9.3
R10339 vss.n20189 vss.n20188 9.3
R10340 vss.n20172 vss.n20171 9.3
R10341 vss.n20173 vss.n20172 9.3
R10342 vss.n20174 vss.n20173 9.3
R10343 vss.n20153 vss.n20152 9.3
R10344 vss.n20154 vss.n20153 9.3
R10345 vss.n20155 vss.n20154 9.3
R10346 vss.n19149 vss.n19148 9.3
R10347 vss.n19150 vss.n19149 9.3
R10348 vss.n20144 vss.n19150 9.3
R10349 vss.n20139 vss.n19158 9.3
R10350 vss.n20139 vss.n20138 9.3
R10351 vss.n20138 vss.n20137 9.3
R10352 vss.n20132 vss.n20131 9.3
R10353 vss.n20132 vss.n19161 9.3
R10354 vss.n19161 vss.n19160 9.3
R10355 vss.n20121 vss.n19167 9.3
R10356 vss.n20122 vss.n20121 9.3
R10357 vss.n20123 vss.n20122 9.3
R10358 vss.n20117 vss.n20116 9.3
R10359 vss.n20116 vss.n20115 9.3
R10360 vss.n20115 vss.n20114 9.3
R10361 vss.n20109 vss.n20108 9.3
R10362 vss.n20109 vss.n19181 9.3
R10363 vss.n19181 vss.n19180 9.3
R10364 vss.n20098 vss.n19186 9.3
R10365 vss.n20099 vss.n20098 9.3
R10366 vss.n20100 vss.n20099 9.3
R10367 vss.n20094 vss.n20093 9.3
R10368 vss.n20093 vss.n20092 9.3
R10369 vss.n20092 vss.n20091 9.3
R10370 vss.n20079 vss.n19202 9.3
R10371 vss.n20079 vss.n20078 9.3
R10372 vss.n20078 vss.n20077 9.3
R10373 vss.n20061 vss.n20060 9.3
R10374 vss.n20062 vss.n20061 9.3
R10375 vss.n20063 vss.n20062 9.3
R10376 vss.n20046 vss.n20045 9.3
R10377 vss.n20045 vss.n19229 9.3
R10378 vss.n19229 vss.n19228 9.3
R10379 vss.n20028 vss.n19240 9.3
R10380 vss.n20028 vss.n19247 9.3
R10381 vss.n19247 vss.n19246 9.3
R10382 vss.n20024 vss.n20023 9.3
R10383 vss.n20023 vss.n20022 9.3
R10384 vss.n20022 vss.n20021 9.3
R10385 vss.n20016 vss.n20015 9.3
R10386 vss.n20016 vss.n19259 9.3
R10387 vss.n19259 vss.n19258 9.3
R10388 vss.n20005 vss.n19264 9.3
R10389 vss.n20006 vss.n20005 9.3
R10390 vss.n20007 vss.n20006 9.3
R10391 vss.n20001 vss.n20000 9.3
R10392 vss.n20000 vss.n19999 9.3
R10393 vss.n19999 vss.n19998 9.3
R10394 vss.n19993 vss.n19992 9.3
R10395 vss.n19993 vss.n19278 9.3
R10396 vss.n19278 vss.n19277 9.3
R10397 vss.n19982 vss.n19283 9.3
R10398 vss.n19983 vss.n19982 9.3
R10399 vss.n19984 vss.n19983 9.3
R10400 vss.n19978 vss.n19977 9.3
R10401 vss.n19977 vss.n19976 9.3
R10402 vss.n19976 vss.n19975 9.3
R10403 vss.n19971 vss.n19970 9.3
R10404 vss.n19972 vss.n19971 9.3
R10405 vss.n19973 vss.n19972 9.3
R10406 vss.n19956 vss.n19955 9.3
R10407 vss.n19955 vss.n19310 9.3
R10408 vss.n19310 vss.n19309 9.3
R10409 vss.n19943 vss.n19324 9.3
R10410 vss.n19943 vss.n19942 9.3
R10411 vss.n19942 vss.n19941 9.3
R10412 vss.n19925 vss.n19924 9.3
R10413 vss.n19926 vss.n19925 9.3
R10414 vss.n19927 vss.n19926 9.3
R10415 vss.n19906 vss.n19905 9.3
R10416 vss.n19907 vss.n19906 9.3
R10417 vss.n19908 vss.n19907 9.3
R10418 vss.n19356 vss.n19355 9.3
R10419 vss.n19357 vss.n19356 9.3
R10420 vss.n19897 vss.n19357 9.3
R10421 vss.n19892 vss.n19365 9.3
R10422 vss.n19892 vss.n19891 9.3
R10423 vss.n19891 vss.n19890 9.3
R10424 vss.n19885 vss.n19884 9.3
R10425 vss.n19885 vss.n19368 9.3
R10426 vss.n19368 vss.n19367 9.3
R10427 vss.n19874 vss.n19374 9.3
R10428 vss.n19875 vss.n19874 9.3
R10429 vss.n19876 vss.n19875 9.3
R10430 vss.n19870 vss.n19869 9.3
R10431 vss.n19869 vss.n19868 9.3
R10432 vss.n19868 vss.n19867 9.3
R10433 vss.n19862 vss.n19861 9.3
R10434 vss.n19862 vss.n19388 9.3
R10435 vss.n19388 vss.n19387 9.3
R10436 vss.n19851 vss.n19393 9.3
R10437 vss.n19852 vss.n19851 9.3
R10438 vss.n19853 vss.n19852 9.3
R10439 vss.n19847 vss.n19846 9.3
R10440 vss.n19846 vss.n19845 9.3
R10441 vss.n19845 vss.n19844 9.3
R10442 vss.n19832 vss.n19409 9.3
R10443 vss.n19832 vss.n19831 9.3
R10444 vss.n19831 vss.n19830 9.3
R10445 vss.n19814 vss.n19813 9.3
R10446 vss.n19815 vss.n19814 9.3
R10447 vss.n19816 vss.n19815 9.3
R10448 vss.n19799 vss.n19798 9.3
R10449 vss.n19798 vss.n19436 9.3
R10450 vss.n19436 vss.n19435 9.3
R10451 vss.n19781 vss.n19447 9.3
R10452 vss.n19781 vss.n19454 9.3
R10453 vss.n19454 vss.n19453 9.3
R10454 vss.n19777 vss.n19776 9.3
R10455 vss.n19776 vss.n19775 9.3
R10456 vss.n19775 vss.n19774 9.3
R10457 vss.n19769 vss.n19768 9.3
R10458 vss.n19769 vss.n19466 9.3
R10459 vss.n19466 vss.n19465 9.3
R10460 vss.n19758 vss.n19471 9.3
R10461 vss.n19759 vss.n19758 9.3
R10462 vss.n19760 vss.n19759 9.3
R10463 vss.n19754 vss.n19753 9.3
R10464 vss.n19753 vss.n19752 9.3
R10465 vss.n19752 vss.n19751 9.3
R10466 vss.n19746 vss.n19745 9.3
R10467 vss.n19746 vss.n19485 9.3
R10468 vss.n19485 vss.n19484 9.3
R10469 vss.n19735 vss.n19490 9.3
R10470 vss.n19736 vss.n19735 9.3
R10471 vss.n19737 vss.n19736 9.3
R10472 vss.n19731 vss.n19730 9.3
R10473 vss.n19730 vss.n19729 9.3
R10474 vss.n19729 vss.n19728 9.3
R10475 vss.n19724 vss.n19723 9.3
R10476 vss.n19725 vss.n19724 9.3
R10477 vss.n19726 vss.n19725 9.3
R10478 vss.n19709 vss.n19708 9.3
R10479 vss.n19708 vss.n19517 9.3
R10480 vss.n19517 vss.n19516 9.3
R10481 vss.n19696 vss.n19531 9.3
R10482 vss.n19696 vss.n19695 9.3
R10483 vss.n19695 vss.n19694 9.3
R10484 vss.n19678 vss.n19677 9.3
R10485 vss.n19679 vss.n19678 9.3
R10486 vss.n19680 vss.n19679 9.3
R10487 vss.n19659 vss.n19658 9.3
R10488 vss.n19660 vss.n19659 9.3
R10489 vss.n19661 vss.n19660 9.3
R10490 vss.n19563 vss.n19562 9.3
R10491 vss.n19564 vss.n19563 9.3
R10492 vss.n19650 vss.n19564 9.3
R10493 vss.n19645 vss.n19572 9.3
R10494 vss.n19645 vss.n19644 9.3
R10495 vss.n19644 vss.n19643 9.3
R10496 vss.n19638 vss.n19637 9.3
R10497 vss.n19638 vss.n19575 9.3
R10498 vss.n19575 vss.n19574 9.3
R10499 vss.n19627 vss.n19581 9.3
R10500 vss.n19628 vss.n19627 9.3
R10501 vss.n19629 vss.n19628 9.3
R10502 vss.n19590 vss.n19587 9.3
R10503 vss.n19602 vss.n19590 9.3
R10504 vss.n19602 vss.n19601 9.3
R10505 vss.n19608 vss.n19595 9.3
R10506 vss.n20304 vss.n17558 9.3
R10507 vss.n20295 vss.n17556 9.3
R10508 vss.n17535 vss.n17534 9.3
R10509 vss.n17537 vss.n17536 9.3
R10510 vss.n17533 vss.n17532 9.3
R10511 vss.n17540 vss.n17539 9.3
R10512 vss.n17545 vss.n17544 9.3
R10513 vss.n17542 vss.n17541 9.3
R10514 vss.n20456 vss.n20455 9.3
R10515 vss.n20472 vss.n20471 9.3
R10516 vss.n20487 vss.n20486 9.3
R10517 vss.n20502 vss.n20501 9.3
R10518 vss.n20518 vss.n20517 9.3
R10519 vss.n20536 vss.n20535 9.3
R10520 vss.n20546 vss.n20545 9.3
R10521 vss.n20565 vss.n20564 9.3
R10522 vss.n20580 vss.n20579 9.3
R10523 vss.n20576 vss.n20575 9.3
R10524 vss.n20575 vss.n20574 9.3
R10525 vss.n20574 vss.n20573 9.3
R10526 vss.n20563 vss.n20562 9.3
R10527 vss.n20520 vss.n20519 9.3
R10528 vss.n20489 vss.n20488 9.3
R10529 vss.n20459 vss.n20458 9.3
R10530 vss.n20454 vss.n20453 9.3
R10531 vss.n20453 vss.n20452 9.3
R10532 vss.n20452 vss.n20451 9.3
R10533 vss.n20470 vss.n20469 9.3
R10534 vss.n20469 vss.n20468 9.3
R10535 vss.n20468 vss.n20467 9.3
R10536 vss.n20474 vss.n20473 9.3
R10537 vss.n20485 vss.n20484 9.3
R10538 vss.n20484 vss.n20483 9.3
R10539 vss.n20483 vss.n20482 9.3
R10540 vss.n20500 vss.n20499 9.3
R10541 vss.n20499 vss.n20498 9.3
R10542 vss.n20498 vss.n20497 9.3
R10543 vss.n20504 vss.n20503 9.3
R10544 vss.n20516 vss.n20515 9.3
R10545 vss.n20515 vss.n20514 9.3
R10546 vss.n20514 vss.n20513 9.3
R10547 vss.n20534 vss.n20533 9.3
R10548 vss.n20533 vss.n20532 9.3
R10549 vss.n20532 vss.n20531 9.3
R10550 vss.n20538 vss.n20537 9.3
R10551 vss.n20544 vss.n20543 9.3
R10552 vss.n20561 vss.n20560 9.3
R10553 vss.n20560 vss.n20559 9.3
R10554 vss.n20559 vss.n20558 9.3
R10555 vss.n20578 vss.n20577 9.3
R10556 vss.n17490 vss.n17489 9.3
R10557 vss.n17492 vss.n17491 9.3
R10558 vss.n17488 vss.n17487 9.3
R10559 vss.n17495 vss.n17494 9.3
R10560 vss.n17500 vss.n17499 9.3
R10561 vss.n17497 vss.n17496 9.3
R10562 vss.n20595 vss.n20594 9.3
R10563 vss.n20610 vss.n20609 9.3
R10564 vss.n20625 vss.n20624 9.3
R10565 vss.n20640 vss.n20639 9.3
R10566 vss.n20671 vss.n20670 9.3
R10567 vss.n20686 vss.n20685 9.3
R10568 vss.n20701 vss.n20700 9.3
R10569 vss.n20716 vss.n20715 9.3
R10570 vss.n20731 vss.n20730 9.3
R10571 vss.n20746 vss.n20745 9.3
R10572 vss.n20787 vss.n20786 9.3
R10573 vss.n20803 vss.n20802 9.3
R10574 vss.n20818 vss.n20817 9.3
R10575 vss.n20833 vss.n20832 9.3
R10576 vss.n20849 vss.n20848 9.3
R10577 vss.n20860 vss.n20859 9.3
R10578 vss.n20859 vss.n20858 9.3
R10579 vss.n20858 vss.n20857 9.3
R10580 vss.n20847 vss.n20846 9.3
R10581 vss.n20829 vss.n20828 9.3
R10582 vss.n20828 vss.n20827 9.3
R10583 vss.n20827 vss.n20826 9.3
R10584 vss.n20816 vss.n20815 9.3
R10585 vss.n20798 vss.n20797 9.3
R10586 vss.n20797 vss.n20796 9.3
R10587 vss.n20796 vss.n20795 9.3
R10588 vss.n20785 vss.n20784 9.3
R10589 vss.n20748 vss.n20747 9.3
R10590 vss.n20718 vss.n20717 9.3
R10591 vss.n20688 vss.n20687 9.3
R10592 vss.n20658 vss.n20657 9.3
R10593 vss.n17527 vss.n17526 9.3
R10594 vss.n17526 vss.n17525 9.3
R10595 vss.n20653 vss.n20652 9.3
R10596 vss.n20636 vss.n20635 9.3
R10597 vss.n20635 vss.n20634 9.3
R10598 vss.n20634 vss.n20633 9.3
R10599 vss.n20623 vss.n20622 9.3
R10600 vss.n20606 vss.n20605 9.3
R10601 vss.n20605 vss.n20604 9.3
R10602 vss.n20604 vss.n20603 9.3
R10603 vss.n20593 vss.n20592 9.3
R10604 vss.n20591 vss.n20590 9.3
R10605 vss.n20590 vss.n20589 9.3
R10606 vss.n20589 vss.n20588 9.3
R10607 vss.n20608 vss.n20607 9.3
R10608 vss.n20621 vss.n20620 9.3
R10609 vss.n20620 vss.n20619 9.3
R10610 vss.n20619 vss.n20618 9.3
R10611 vss.n20638 vss.n20637 9.3
R10612 vss.n20651 vss.n20650 9.3
R10613 vss.n20650 vss.n20649 9.3
R10614 vss.n20649 vss.n20648 9.3
R10615 vss.n17514 vss.n17513 9.3
R10616 vss.n17513 vss.n17512 9.3
R10617 vss.n20669 vss.n20668 9.3
R10618 vss.n20668 vss.n20667 9.3
R10619 vss.n20667 vss.n20666 9.3
R10620 vss.n20673 vss.n20672 9.3
R10621 vss.n20684 vss.n20683 9.3
R10622 vss.n20683 vss.n20682 9.3
R10623 vss.n20682 vss.n20681 9.3
R10624 vss.n20699 vss.n20698 9.3
R10625 vss.n20698 vss.n20697 9.3
R10626 vss.n20697 vss.n20696 9.3
R10627 vss.n20703 vss.n20702 9.3
R10628 vss.n20714 vss.n20713 9.3
R10629 vss.n20713 vss.n20712 9.3
R10630 vss.n20712 vss.n20711 9.3
R10631 vss.n20729 vss.n20728 9.3
R10632 vss.n20728 vss.n20727 9.3
R10633 vss.n20727 vss.n20726 9.3
R10634 vss.n20733 vss.n20732 9.3
R10635 vss.n20744 vss.n20743 9.3
R10636 vss.n20743 vss.n20742 9.3
R10637 vss.n20742 vss.n20741 9.3
R10638 vss.n20763 vss.n20762 9.3
R10639 vss.n20762 vss.n20761 9.3
R10640 vss.n20761 vss.n20760 9.3
R10641 vss.n20783 vss.n20782 9.3
R10642 vss.n20782 vss.n20781 9.3
R10643 vss.n20781 vss.n20780 9.3
R10644 vss.n20801 vss.n20800 9.3
R10645 vss.n20814 vss.n20813 9.3
R10646 vss.n20813 vss.n20812 9.3
R10647 vss.n20812 vss.n20811 9.3
R10648 vss.n20831 vss.n20830 9.3
R10649 vss.n20844 vss.n20843 9.3
R10650 vss.n20843 vss.n20842 9.3
R10651 vss.n20842 vss.n20841 9.3
R10652 vss.n17483 vss.n17482 9.3
R10653 vss.n17482 vss.n17481 9.3
R10654 vss.n20906 vss.n20905 9.3
R10655 vss.n20905 vss.n20904 9.3
R10656 vss.n20920 vss.n20919 9.3
R10657 vss.n20919 vss.n20918 9.3
R10658 vss.n20934 vss.n20933 9.3
R10659 vss.n20933 vss.n20932 9.3
R10660 vss.n20948 vss.n20947 9.3
R10661 vss.n20947 vss.n20946 9.3
R10662 vss.n20962 vss.n20961 9.3
R10663 vss.n20961 vss.n20960 9.3
R10664 vss.n20976 vss.n20975 9.3
R10665 vss.n20975 vss.n20974 9.3
R10666 vss.n20992 vss.n20991 9.3
R10667 vss.n20991 vss.n20990 9.3
R10668 vss.n21011 vss.n21010 9.3
R10669 vss.n21010 vss.n21009 9.3
R10670 vss.n21025 vss.n21024 9.3
R10671 vss.n21024 vss.n21023 9.3
R10672 vss.n21039 vss.n21038 9.3
R10673 vss.n21038 vss.n21037 9.3
R10674 vss.n21053 vss.n21052 9.3
R10675 vss.n21052 vss.n21051 9.3
R10676 vss.n21067 vss.n21066 9.3
R10677 vss.n21066 vss.n21065 9.3
R10678 vss.n21081 vss.n21080 9.3
R10679 vss.n21080 vss.n21079 9.3
R10680 vss.n21095 vss.n21094 9.3
R10681 vss.n21094 vss.n21093 9.3
R10682 vss.n17472 vss.n17471 9.3
R10683 vss.n17471 vss.n17470 9.3
R10684 vss.n17461 vss.n17460 9.3
R10685 vss.n17460 vss.n17459 9.3
R10686 vss.n21114 vss.n21113 9.3
R10687 vss.n21113 vss.n21112 9.3
R10688 vss.n21128 vss.n21127 9.3
R10689 vss.n21127 vss.n21126 9.3
R10690 vss.n21142 vss.n21141 9.3
R10691 vss.n21141 vss.n21140 9.3
R10692 vss.n21156 vss.n21155 9.3
R10693 vss.n21155 vss.n21154 9.3
R10694 vss.n21170 vss.n21169 9.3
R10695 vss.n21169 vss.n21168 9.3
R10696 vss.n21184 vss.n21183 9.3
R10697 vss.n21183 vss.n21182 9.3
R10698 vss.n21200 vss.n21199 9.3
R10699 vss.n21199 vss.n21198 9.3
R10700 vss.n21219 vss.n21218 9.3
R10701 vss.n21218 vss.n21217 9.3
R10702 vss.n21233 vss.n21232 9.3
R10703 vss.n21232 vss.n21231 9.3
R10704 vss.n21247 vss.n21246 9.3
R10705 vss.n21246 vss.n21245 9.3
R10706 vss.n21261 vss.n21260 9.3
R10707 vss.n21260 vss.n21259 9.3
R10708 vss.n21275 vss.n21274 9.3
R10709 vss.n21274 vss.n21273 9.3
R10710 vss.n21289 vss.n21288 9.3
R10711 vss.n21288 vss.n21287 9.3
R10712 vss.n21303 vss.n21302 9.3
R10713 vss.n21302 vss.n21301 9.3
R10714 vss.n17450 vss.n17449 9.3
R10715 vss.n17449 vss.n17448 9.3
R10716 vss.n17439 vss.n17438 9.3
R10717 vss.n17438 vss.n17437 9.3
R10718 vss.n21322 vss.n21321 9.3
R10719 vss.n21321 vss.n21320 9.3
R10720 vss.n21336 vss.n21335 9.3
R10721 vss.n21335 vss.n21334 9.3
R10722 vss.n21350 vss.n21349 9.3
R10723 vss.n21349 vss.n21348 9.3
R10724 vss.n21364 vss.n21363 9.3
R10725 vss.n21363 vss.n21362 9.3
R10726 vss.n21378 vss.n21377 9.3
R10727 vss.n21377 vss.n21376 9.3
R10728 vss.n21392 vss.n21391 9.3
R10729 vss.n21391 vss.n21390 9.3
R10730 vss.n21408 vss.n21407 9.3
R10731 vss.n21407 vss.n21406 9.3
R10732 vss.n21427 vss.n21426 9.3
R10733 vss.n21426 vss.n21425 9.3
R10734 vss.n21441 vss.n21440 9.3
R10735 vss.n21440 vss.n21439 9.3
R10736 vss.n21455 vss.n21454 9.3
R10737 vss.n21454 vss.n21453 9.3
R10738 vss.n21469 vss.n21468 9.3
R10739 vss.n21468 vss.n21467 9.3
R10740 vss.n21483 vss.n21482 9.3
R10741 vss.n21482 vss.n21481 9.3
R10742 vss.n21497 vss.n21496 9.3
R10743 vss.n21496 vss.n21495 9.3
R10744 vss.n21511 vss.n21510 9.3
R10745 vss.n21510 vss.n21509 9.3
R10746 vss.n17428 vss.n17427 9.3
R10747 vss.n17427 vss.n17426 9.3
R10748 vss.n17417 vss.n17416 9.3
R10749 vss.n17416 vss.n17415 9.3
R10750 vss.n21530 vss.n21529 9.3
R10751 vss.n21529 vss.n21528 9.3
R10752 vss.n21544 vss.n21543 9.3
R10753 vss.n21543 vss.n21542 9.3
R10754 vss.n21558 vss.n21557 9.3
R10755 vss.n21557 vss.n21556 9.3
R10756 vss.n21572 vss.n21571 9.3
R10757 vss.n21571 vss.n21570 9.3
R10758 vss.n17407 vss.n17406 9.3
R10759 vss.n17406 vss.n17405 9.3
R10760 vss.n21588 vss.n21587 9.3
R10761 vss.n21587 vss.n21586 9.3
R10762 vss.n21867 vss.n21866 9.3
R10763 vss.n21878 vss.n21877 9.3
R10764 vss.n21865 vss.n21864 9.3
R10765 vss.n21874 vss.n21873 9.3
R10766 vss.n21873 vss.n21872 9.3
R10767 vss.n21876 vss.n21875 9.3
R10768 vss.n21885 vss.n21884 9.3
R10769 vss.n21884 vss.n21883 9.3
R10770 vss.n21860 vss.n21859 9.3
R10771 vss.n21842 vss.n21841 9.3
R10772 vss.n21841 vss.n21840 9.3
R10773 vss.n21826 vss.n21825 9.3
R10774 vss.n21835 vss.n21834 9.3
R10775 vss.n21834 vss.n21833 9.3
R10776 vss.n21828 vss.n21827 9.3
R10777 vss.n21844 vss.n21843 9.3
R10778 vss.n21846 vss.n21845 9.3
R10779 vss.n21854 vss.n21853 9.3
R10780 vss.n21853 vss.n21852 9.3
R10781 vss.n21905 vss.n21904 9.3
R10782 vss.n21856 vss.n21855 9.3
R10783 vss.n21937 vss.n21936 9.3
R10784 vss.n21930 vss.n21929 9.3
R10785 vss.n21932 vss.n21931 9.3
R10786 vss.n21934 vss.n21933 9.3
R10787 vss.n22004 vss.n22003 9.3
R10788 vss.n22011 vss.n22010 9.3
R10789 vss.n22024 vss.n22023 9.3
R10790 vss.n22018 vss.n22017 9.3
R10791 vss.n21808 vss.n21807 9.3
R10792 vss.n22020 vss.n22019 9.3
R10793 vss.n22022 vss.n22021 9.3
R10794 vss.n22026 vss.n22025 9.3
R10795 vss.n22014 vss.n22013 9.3
R10796 vss.n22009 vss.n22008 9.3
R10797 vss.n22007 vss.n22006 9.3
R10798 vss.n22002 vss.n22001 9.3
R10799 vss.n22046 vss.n22045 9.3
R10800 vss.n22041 vss.n22040 9.3
R10801 vss.n22036 vss.n22035 9.3
R10802 vss.n22043 vss.n22042 9.3
R10803 vss.n22034 vss.n22033 9.3
R10804 vss.n22039 vss.n22038 9.3
R10805 vss.n22048 vss.n22047 9.3
R10806 vss.n21973 vss.n21972 9.3
R10807 vss.n21969 vss.n21968 9.3
R10808 vss.n21961 vss.n21960 9.3
R10809 vss.n21957 vss.n21956 9.3
R10810 vss.n21959 vss.n21958 9.3
R10811 vss.n21964 vss.n21963 9.3
R10812 vss.n22049 vss.n21985 9.3
R10813 vss.n21712 vss.n21711 9.3
R10814 vss.n21747 vss.n21746 9.3
R10815 vss.n21742 vss.n21705 9.3
R10816 vss.n21743 vss.n21742 9.3
R10817 vss.n21740 vss.n21739 9.3
R10818 vss.n21723 vss.n21720 9.3
R10819 vss.n21722 vss.n21721 9.3
R10820 vss.n21725 vss.n21724 9.3
R10821 vss.n21726 vss.n21725 9.3
R10822 vss.n21735 vss.n21717 9.3
R10823 vss.n21735 vss.n21734 9.3
R10824 vss.n21738 vss.n21737 9.3
R10825 vss.n21736 vss.n21715 9.3
R10826 vss.n21769 vss.n21761 9.3
R10827 vss.n21764 vss.n21762 9.3
R10828 vss.n21771 vss.n21770 9.3
R10829 vss.n21768 vss.n21767 9.3
R10830 vss.n21766 vss.n21765 9.3
R10831 vss.n21763 vss.n21687 9.3
R10832 vss.n21784 vss.n21775 9.3
R10833 vss.n21779 vss.n21776 9.3
R10834 vss.n21793 vss.n21686 9.3
R10835 vss.n21694 vss.n21685 9.3
R10836 vss.n21778 vss.n21777 9.3
R10837 vss.n21781 vss.n21780 9.3
R10838 vss.n21783 vss.n21782 9.3
R10839 vss.n21786 vss.n21785 9.3
R10840 vss.n21792 vss.n21791 9.3
R10841 vss.n21683 vss.n21682 9.3
R10842 vss.n21677 vss.n21665 9.3
R10843 vss.n21674 vss.n21673 9.3
R10844 vss.n21684 vss.n21664 9.3
R10845 vss.n21681 vss.n21680 9.3
R10846 vss.n21679 vss.n21678 9.3
R10847 vss.n21676 vss.n21675 9.3
R10848 vss.n21672 vss.n21671 9.3
R10849 vss.n21652 vss.n21646 9.3
R10850 vss.n21654 vss.n21653 9.3
R10851 vss.n21668 vss.n21667 9.3
R10852 vss.n21648 vss.n21642 9.3
R10853 vss.n21796 vss.n21648 9.3
R10854 vss.n21799 vss.n21798 9.3
R10855 vss.n21657 vss.n21656 9.3
R10856 vss.n21602 vss.n21601 9.3
R10857 vss.n21601 vss.n21600 9.3
R10858 vss.n22065 vss.n22064 9.3
R10859 vss.n22058 vss.n22057 9.3
R10860 vss.n21639 vss.n21638 9.3
R10861 vss.n22056 vss.n22055 9.3
R10862 vss.n22060 vss.n22059 9.3
R10863 vss.n22063 vss.n22062 9.3
R10864 vss.n22067 vss.n22066 9.3
R10865 vss.n10317 vss.n10316 9.3
R10866 vss.n10349 vss.n10340 9.3
R10867 vss.n10350 vss.n10339 9.3
R10868 vss.n10352 vss.n10324 9.3
R10869 vss.n10384 vss.n10365 9.3
R10870 vss.n10382 vss.n10366 9.3
R10871 vss.n10385 vss.n10358 9.3
R10872 vss.n10413 vss.n10398 9.3
R10873 vss.n10415 vss.n10414 9.3
R10874 vss.n10397 vss.n10396 9.3
R10875 vss.n10427 vss.n10426 9.3
R10876 vss.n8986 vss.n8985 9.3
R10877 vss.n8988 vss.n8987 9.3
R10878 vss.n8983 vss.n8982 9.3
R10879 vss.n9016 vss.n9015 9.3
R10880 vss.n9018 vss.n9017 9.3
R10881 vss.n9013 vss.n9012 9.3
R10882 vss.n9047 vss.n9046 9.3
R10883 vss.n9049 vss.n9048 9.3
R10884 vss.n9044 vss.n9043 9.3
R10885 vss.n9078 vss.n9077 9.3
R10886 vss.n9080 vss.n9079 9.3
R10887 vss.n9075 vss.n9074 9.3
R10888 vss.n9098 vss.n9097 9.3
R10889 vss.n9123 vss.n9122 9.3
R10890 vss.n9150 vss.n9149 9.3
R10891 vss.n12279 vss.n12277 9.3
R10892 vss.n10777 vss.n10776 9.3
R10893 vss.n13478 vss.n13476 9.3
R10894 vss.n13405 vss.n13404 9.3
R10895 vss.n12883 vss.n12882 9.3
R10896 vss.n12914 vss.n12913 9.3
R10897 vss.n12808 vss.n12807 9.3
R10898 vss.n15048 vss.n15047 9.3
R10899 vss.n12474 vss.n12473 9.3
R10900 vss.n12501 vss.n12500 9.3
R10901 vss.n12552 vss.n12551 9.3
R10902 vss.n12906 vss.n12905 9.3
R10903 vss.n12901 vss.n12900 9.3
R10904 vss.n12921 vss.n12920 9.3
R10905 vss.n12920 vss.n12919 9.3
R10906 vss.n12822 vss.n12821 9.3
R10907 vss.n12815 vss.n12814 9.3
R10908 vss.n12814 vss.n12813 9.3
R10909 vss.n15056 vss.n15055 9.3
R10910 vss.n15055 vss.n15054 9.3
R10911 vss.n12493 vss.n12492 9.3
R10912 vss.n12636 vss.n12635 9.3
R10913 vss.n12508 vss.n12507 9.3
R10914 vss.n12507 vss.n12506 9.3
R10915 vss.n12489 vss.n12488 9.3
R10916 vss.n12559 vss.n12558 9.3
R10917 vss.n12558 vss.n12557 9.3
R10918 vss.n12604 vss.n12603 9.3
R10919 vss.n12621 vss.n12620 9.3
R10920 vss.n12632 vss.n12631 9.3
R10921 vss.n12619 vss.n12618 9.3
R10922 vss.n12618 vss.n12617 9.3
R10923 vss.n12617 vss.n12616 9.3
R10924 vss.n12607 vss.n12606 9.3
R10925 vss.n12602 vss.n12601 9.3
R10926 vss.n12601 vss.n12600 9.3
R10927 vss.n12600 vss.n12599 9.3
R10928 vss.n12529 vss.n12528 9.3
R10929 vss.n12528 vss.n12527 9.3
R10930 vss.n12519 vss.n12518 9.3
R10931 vss.n12629 vss.n12627 9.3
R10932 vss.n12131 vss.n12130 9.3
R10933 vss.n12130 vss.n12129 9.3
R10934 vss.n12121 vss.n12120 9.3
R10935 vss.n12120 vss.n12119 9.3
R10936 vss.n12145 vss.n12144 9.3
R10937 vss.n12144 vss.n12143 9.3
R10938 vss.n12586 vss.n12585 9.3
R10939 vss.n12585 vss.n12584 9.3
R10940 vss.n12568 vss.n12567 9.3
R10941 vss.n12219 vss.n12218 9.3
R10942 vss.n12013 vss.n12012 9.3
R10943 vss.n11328 vss.n11327 9.3
R10944 vss.n11303 vss.n11302 9.3
R10945 vss.n11287 vss.n11286 9.3
R10946 vss.n11261 vss.n11260 9.3
R10947 vss.n11189 vss.n11188 9.3
R10948 vss.n11173 vss.n11172 9.3
R10949 vss.n11152 vss.n11151 9.3
R10950 vss.n11075 vss.n11074 9.3
R10951 vss.n11074 vss.n11073 9.3
R10952 vss.n11085 vss.n11084 9.3
R10953 vss.n11084 vss.n11083 9.3
R10954 vss.n11215 vss.n10995 9.3
R10955 vss.n11221 vss.n11220 9.3
R10956 vss.n11259 vss.n11258 9.3
R10957 vss.n11258 vss.n11257 9.3
R10958 vss.n11257 vss.n11256 9.3
R10959 vss.n11301 vss.n11300 9.3
R10960 vss.n11300 vss.n11299 9.3
R10961 vss.n11299 vss.n11298 9.3
R10962 vss.n11924 vss.n11923 9.3
R10963 vss.n11923 vss.n11922 9.3
R10964 vss.n11922 vss.n11921 9.3
R10965 vss.n11967 vss.n10881 9.3
R10966 vss.n10881 vss.n10880 9.3
R10967 vss.n10880 vss.n10879 9.3
R10968 vss.n11982 vss.n11981 9.3
R10969 vss.n10836 vss.n10835 9.3
R10970 vss.n10857 vss.n10856 9.3
R10971 vss.n10856 vss.n10855 9.3
R10972 vss.n11992 vss.n11991 9.3
R10973 vss.n11991 vss.n11990 9.3
R10974 vss.n11990 vss.n11989 9.3
R10975 vss.n12072 vss.n12071 9.3
R10976 vss.n12071 vss.n12070 9.3
R10977 vss.n12202 vss.n12201 9.3
R10978 vss.n12201 vss.n12200 9.3
R10979 vss.n12200 vss.n12199 9.3
R10980 vss.n12188 vss.n12187 9.3
R10981 vss.n12187 vss.n12186 9.3
R10982 vss.n12186 vss.n12185 9.3
R10983 vss.n12204 vss.n12203 9.3
R10984 vss.n12162 vss.n12095 9.3
R10985 vss.n12176 vss.n12175 9.3
R10986 vss.n12174 vss.n12173 9.3
R10987 vss.n12173 vss.n12172 9.3
R10988 vss.n12172 vss.n12171 9.3
R10989 vss.n12164 vss.n12163 9.3
R10990 vss.n12158 vss.n12157 9.3
R10991 vss.n12157 vss.n12156 9.3
R10992 vss.n12156 vss.n12155 9.3
R10993 vss.n12162 vss.n12161 9.3
R10994 vss.n12160 vss.n12159 9.3
R10995 vss.n12178 vss.n12177 9.3
R10996 vss.n12237 vss.n12236 9.3
R10997 vss.n12082 vss.n12081 9.3
R10998 vss.n12081 vss.n12080 9.3
R10999 vss.n12061 vss.n12060 9.3
R11000 vss.n12215 vss.n12214 9.3
R11001 vss.n12214 vss.n12213 9.3
R11002 vss.n12213 vss.n12212 9.3
R11003 vss.n12206 vss.n12205 9.3
R11004 vss.n12192 vss.n12191 9.3
R11005 vss.n12190 vss.n12189 9.3
R11006 vss.n12217 vss.n12216 9.3
R11007 vss.n12229 vss.n12228 9.3
R11008 vss.n12228 vss.n12227 9.3
R11009 vss.n12227 vss.n12226 9.3
R11010 vss.n12242 vss.n12241 9.3
R11011 vss.n12247 vss.n12246 9.3
R11012 vss.n12055 vss.n12054 9.3
R11013 vss.n12054 vss.n12053 9.3
R11014 vss.n12045 vss.n12044 9.3
R11015 vss.n12044 vss.n12043 9.3
R11016 vss.n12267 vss.n12266 9.3
R11017 vss.n12025 vss.n12024 9.3
R11018 vss.n10801 vss.n10800 9.3
R11019 vss.n10800 vss.n10799 9.3
R11020 vss.n12023 vss.n12022 9.3
R11021 vss.n12022 vss.n12021 9.3
R11022 vss.n12021 vss.n12020 9.3
R11023 vss.n12011 vss.n12010 9.3
R11024 vss.n12005 vss.n12004 9.3
R11025 vss.n12004 vss.n12003 9.3
R11026 vss.n11980 vss.n11979 9.3
R11027 vss.n11978 vss.n11977 9.3
R11028 vss.n11977 vss.n11976 9.3
R11029 vss.n11976 vss.n11975 9.3
R11030 vss.n11950 vss.n11949 9.3
R11031 vss.n11949 vss.n11948 9.3
R11032 vss.n11948 vss.n11947 9.3
R11033 vss.n11330 vss.n11329 9.3
R11034 vss.n11326 vss.n11325 9.3
R11035 vss.n11325 vss.n11324 9.3
R11036 vss.n11324 vss.n11323 9.3
R11037 vss.n11305 vss.n11304 9.3
R11038 vss.n11289 vss.n11288 9.3
R11039 vss.n11285 vss.n11284 9.3
R11040 vss.n11284 vss.n11283 9.3
R11041 vss.n11283 vss.n11282 9.3
R11042 vss.n11263 vss.n11262 9.3
R11043 vss.n11224 vss.n11223 9.3
R11044 vss.n10964 vss.n10963 9.3
R11045 vss.n10963 vss.n10962 9.3
R11046 vss.n10974 vss.n10973 9.3
R11047 vss.n10973 vss.n10972 9.3
R11048 vss.n11271 vss.n11270 9.3
R11049 vss.n11024 vss.n11023 9.3
R11050 vss.n11053 vss.n11052 9.3
R11051 vss.n11052 vss.n11051 9.3
R11052 vss.n11043 vss.n11042 9.3
R11053 vss.n11042 vss.n11041 9.3
R11054 vss.n10984 vss.n10983 9.3
R11055 vss.n10983 vss.n10982 9.3
R11056 vss.n11004 vss.n11003 9.3
R11057 vss.n11003 vss.n11002 9.3
R11058 vss.n11201 vss.n11027 9.3
R11059 vss.n11186 vss.n11185 9.3
R11060 vss.n11199 vss.n11198 9.3
R11061 vss.n11198 vss.n11197 9.3
R11062 vss.n11197 vss.n11196 9.3
R11063 vss.n11183 vss.n11182 9.3
R11064 vss.n11182 vss.n11181 9.3
R11065 vss.n11181 vss.n11180 9.3
R11066 vss.n11171 vss.n11170 9.3
R11067 vss.n11150 vss.n11149 9.3
R11068 vss.n11162 vss.n11161 9.3
R11069 vss.n11161 vss.n11160 9.3
R11070 vss.n11160 vss.n11159 9.3
R11071 vss.n11095 vss.n11094 9.3
R11072 vss.n11094 vss.n11093 9.3
R11073 vss.n11065 vss.n11064 9.3
R11074 vss.n11064 vss.n11063 9.3
R11075 vss.n10916 vss.n10915 9.3
R11076 vss.n11891 vss.n11890 9.3
R11077 vss.n11359 vss.n11358 9.3
R11078 vss.n11415 vss.n11414 9.3
R11079 vss.n11403 vss.n11402 9.3
R11080 vss.n13711 vss.n13710 9.3
R11081 vss.n14130 vss.n14129 9.3
R11082 vss.n13623 vss.n13622 9.3
R11083 vss.n13613 vss.n13612 9.3
R11084 vss.n14138 vss.n14136 9.3
R11085 vss.n11899 vss.n11897 9.3
R11086 vss.n11351 vss.n11350 9.3
R11087 vss.n10760 vss.n10759 9.3
R11088 vss.n10590 vss.n10589 9.3
R11089 vss.n10610 vss.n10608 9.3
R11090 vss.n13046 vss.n13045 9.3
R11091 vss.n10748 vss.n10747 9.3
R11092 vss.n13436 vss.n13435 9.3
R11093 vss.n13427 vss.n13426 9.3
R11094 vss.n10618 vss.n10617 9.3
R11095 vss.n10598 vss.n10597 9.3
R11096 vss.n13034 vss.n13033 9.3
R11097 vss.n10479 vss.n10478 9.3
R11098 vss.n10478 vss.n10477 9.3
R11099 vss.n10509 vss.n10508 9.3
R11100 vss.n10508 vss.n10507 9.3
R11101 vss.n10526 vss.n10525 9.3
R11102 vss.n12417 vss.n12416 9.3
R11103 vss.n12428 vss.n12427 9.3
R11104 vss.n12427 vss.n12426 9.3
R11105 vss.n12456 vss.n12455 9.3
R11106 vss.n12455 vss.n12454 9.3
R11107 vss.n10497 vss.n10496 9.3
R11108 vss.n12467 vss.n12466 9.3
R11109 vss.n12466 vss.n12465 9.3
R11110 vss.n12673 vss.n12672 9.3
R11111 vss.n12672 vss.n12671 9.3
R11112 vss.n12706 vss.n12705 9.3
R11113 vss.n12705 vss.n12704 9.3
R11114 vss.n10519 vss.n10518 9.3
R11115 vss.n10518 vss.n10517 9.3
R11116 vss.n10489 vss.n10488 9.3
R11117 vss.n10488 vss.n10487 9.3
R11118 vss.n10549 vss.n10548 9.3
R11119 vss.n10548 vss.n10547 9.3
R11120 vss.n12690 vss.n12689 9.3
R11121 vss.n12689 vss.n12688 9.3
R11122 vss.n12657 vss.n12656 9.3
R11123 vss.n12656 vss.n12655 9.3
R11124 vss.n12484 vss.n12483 9.3
R11125 vss.n12483 vss.n12482 9.3
R11126 vss.n12436 vss.n12435 9.3
R11127 vss.n10469 vss.n10467 9.3
R11128 vss.n10847 vss.n10846 9.3
R11129 vss.n10846 vss.n10845 9.3
R11130 vss.n10827 vss.n10826 9.3
R11131 vss.n10826 vss.n10825 9.3
R11132 vss.n10816 vss.n10815 9.3
R11133 vss.n10901 vss.n10900 9.3
R11134 vss.n10900 vss.n10899 9.3
R11135 vss.n10923 vss.n10922 9.3
R11136 vss.n10891 vss.n10890 9.3
R11137 vss.n10890 vss.n10889 9.3
R11138 vss.n11217 vss.n11216 9.3
R11139 vss.n10954 vss.n10953 9.3
R11140 vss.n10953 vss.n10952 9.3
R11141 vss.n10941 vss.n10940 9.3
R11142 vss.n11226 vss.n11225 9.3
R11143 vss.n11239 vss.n11238 9.3
R11144 vss.n11248 vss.n11247 9.3
R11145 vss.n11247 vss.n11246 9.3
R11146 vss.n11246 vss.n11245 9.3
R11147 vss.n11014 vss.n11013 9.3
R11148 vss.n11013 vss.n11012 9.3
R11149 vss.n11032 vss.n11031 9.3
R11150 vss.n11213 vss.n11212 9.3
R11151 vss.n11212 vss.n11211 9.3
R11152 vss.n11211 vss.n11210 9.3
R11153 vss.n11215 vss.n11214 9.3
R11154 vss.n11395 vss.n11394 9.3
R11155 vss.n11423 vss.n11422 9.3
R11156 vss.n13699 vss.n13698 9.3
R11157 vss.n14320 vss.n14319 9.3
R11158 vss.n13893 vss.n13868 9.3
R11159 vss.n11729 vss.n11728 9.3
R11160 vss.n11138 vss.n11110 9.3
R11161 vss.n11751 vss.n11750 9.3
R11162 vss.n11788 vss.n11787 9.3
R11163 vss.n11804 vss.n11803 9.3
R11164 vss.n11829 vss.n11828 9.3
R11165 vss.n11616 vss.n11615 9.3
R11166 vss.n14044 vss.n13964 9.3
R11167 vss.n13906 vss.n13905 9.3
R11168 vss.n13872 vss.n13871 9.3
R11169 vss.n14302 vss.n14301 9.3
R11170 vss.n14316 vss.n14315 9.3
R11171 vss.n13827 vss.n13826 9.3
R11172 vss.n13826 vss.n13825 9.3
R11173 vss.n14054 vss.n14053 9.3
R11174 vss.n14053 vss.n14052 9.3
R11175 vss.n14052 vss.n14051 9.3
R11176 vss.n14012 vss.n14011 9.3
R11177 vss.n14011 vss.n14010 9.3
R11178 vss.n11628 vss.n11627 9.3
R11179 vss.n11627 vss.n11626 9.3
R11180 vss.n11626 vss.n11625 9.3
R11181 vss.n11119 vss.n11118 9.3
R11182 vss.n11118 vss.n11117 9.3
R11183 vss.n14391 vss.n14390 9.3
R11184 vss.n14232 vss.n14231 9.3
R11185 vss.n14231 vss.n14230 9.3
R11186 vss.n14222 vss.n14221 9.3
R11187 vss.n14221 vss.n14220 9.3
R11188 vss.n14242 vss.n14241 9.3
R11189 vss.n14241 vss.n14240 9.3
R11190 vss.n14252 vss.n14251 9.3
R11191 vss.n14251 vss.n14250 9.3
R11192 vss.n11651 vss.n11650 9.3
R11193 vss.n11603 vss.n11602 9.3
R11194 vss.n14037 vss.n14036 9.3
R11195 vss.n13925 vss.n13924 9.3
R11196 vss.n13892 vss.n13891 9.3
R11197 vss.n14350 vss.n14349 9.3
R11198 vss.n11109 vss.n11107 9.3
R11199 vss.n11774 vss.n11773 9.3
R11200 vss.n14401 vss.n14400 9.3
R11201 vss.n14400 vss.n14399 9.3
R11202 vss.n14278 vss.n14277 9.3
R11203 vss.n14277 vss.n14276 9.3
R11204 vss.n14360 vss.n14359 9.3
R11205 vss.n14359 vss.n14358 9.3
R11206 vss.n14329 vss.n14328 9.3
R11207 vss.n14328 vss.n14327 9.3
R11208 vss.n14327 vss.n14326 9.3
R11209 vss.n14318 vss.n14290 9.3
R11210 vss.n13884 vss.n13883 9.3
R11211 vss.n13902 vss.n13901 9.3
R11212 vss.n13901 vss.n13900 9.3
R11213 vss.n13900 vss.n13899 9.3
R11214 vss.n13866 vss.n13865 9.3
R11215 vss.n13865 vss.n13864 9.3
R11216 vss.n13843 vss.n13842 9.3
R11217 vss.n13969 vss.n13968 9.3
R11218 vss.n13981 vss.n13980 9.3
R11219 vss.n13980 vss.n13979 9.3
R11220 vss.n14002 vss.n14001 9.3
R11221 vss.n14001 vss.n14000 9.3
R11222 vss.n11594 vss.n11593 9.3
R11223 vss.n11593 vss.n11592 9.3
R11224 vss.n11576 vss.n11575 9.3
R11225 vss.n11575 vss.n11574 9.3
R11226 vss.n11564 vss.n11563 9.3
R11227 vss.n11703 vss.n11702 9.3
R11228 vss.n11763 vss.n11762 9.3
R11229 vss.n11762 vss.n11761 9.3
R11230 vss.n11738 vss.n11737 9.3
R11231 vss.n11737 vss.n11736 9.3
R11232 vss.n11736 vss.n11735 9.3
R11233 vss.n11727 vss.n11726 9.3
R11234 vss.n11136 vss.n11135 9.3
R11235 vss.n11146 vss.n11145 9.3
R11236 vss.n11145 vss.n11144 9.3
R11237 vss.n11144 vss.n11143 9.3
R11238 vss.n11138 vss.n11137 9.3
R11239 vss.n11132 vss.n11131 9.3
R11240 vss.n11129 vss.n11128 9.3
R11241 vss.n11128 vss.n11127 9.3
R11242 vss.n11721 vss.n11720 9.3
R11243 vss.n11720 vss.n11719 9.3
R11244 vss.n11725 vss.n11724 9.3
R11245 vss.n11753 vss.n11752 9.3
R11246 vss.n11749 vss.n11748 9.3
R11247 vss.n11748 vss.n11747 9.3
R11248 vss.n11747 vss.n11746 9.3
R11249 vss.n11786 vss.n11785 9.3
R11250 vss.n11785 vss.n11784 9.3
R11251 vss.n11784 vss.n11783 9.3
R11252 vss.n11790 vss.n11789 9.3
R11253 vss.n11806 vss.n11805 9.3
R11254 vss.n11802 vss.n11801 9.3
R11255 vss.n11801 vss.n11800 9.3
R11256 vss.n11800 vss.n11799 9.3
R11257 vss.n11827 vss.n11826 9.3
R11258 vss.n11826 vss.n11825 9.3
R11259 vss.n11825 vss.n11824 9.3
R11260 vss.n11831 vss.n11830 9.3
R11261 vss.n11677 vss.n11676 9.3
R11262 vss.n11676 vss.n11675 9.3
R11263 vss.n11675 vss.n11674 9.3
R11264 vss.n11666 vss.n11665 9.3
R11265 vss.n11665 vss.n11664 9.3
R11266 vss.n11664 vss.n11663 9.3
R11267 vss.n11639 vss.n11638 9.3
R11268 vss.n11638 vss.n11637 9.3
R11269 vss.n11637 vss.n11636 9.3
R11270 vss.n11618 vss.n11617 9.3
R11271 vss.n11614 vss.n11613 9.3
R11272 vss.n11613 vss.n11612 9.3
R11273 vss.n11612 vss.n11611 9.3
R11274 vss.n14043 vss.n14042 9.3
R11275 vss.n13991 vss.n13990 9.3
R11276 vss.n13990 vss.n13989 9.3
R11277 vss.n14056 vss.n14055 9.3
R11278 vss.n13953 vss.n13952 9.3
R11279 vss.n14075 vss.n14074 9.3
R11280 vss.n14074 vss.n14073 9.3
R11281 vss.n13934 vss.n13933 9.3
R11282 vss.n13837 vss.n13836 9.3
R11283 vss.n13836 vss.n13835 9.3
R11284 vss.n13854 vss.n13853 9.3
R11285 vss.n13853 vss.n13852 9.3
R11286 vss.n13929 vss.n13928 9.3
R11287 vss.n13904 vss.n13903 9.3
R11288 vss.n13916 vss.n13915 9.3
R11289 vss.n13915 vss.n13914 9.3
R11290 vss.n13914 vss.n13913 9.3
R11291 vss.n13882 vss.n13881 9.3
R11292 vss.n13881 vss.n13880 9.3
R11293 vss.n13880 vss.n13879 9.3
R11294 vss.n13870 vss.n13869 9.3
R11295 vss.n14304 vss.n14303 9.3
R11296 vss.n14300 vss.n14299 9.3
R11297 vss.n14299 vss.n14298 9.3
R11298 vss.n14298 vss.n14297 9.3
R11299 vss.n14314 vss.n14313 9.3
R11300 vss.n14313 vss.n14312 9.3
R11301 vss.n14312 vss.n14311 9.3
R11302 vss.n14318 vss.n14317 9.3
R11303 vss.n14340 vss.n14339 9.3
R11304 vss.n14339 vss.n14338 9.3
R11305 vss.n14338 vss.n14337 9.3
R11306 vss.n14375 vss.n14374 9.3
R11307 vss.n14374 vss.n14373 9.3
R11308 vss.n14373 vss.n14372 9.3
R11309 vss.n14421 vss.n14420 9.3
R11310 vss.n14420 vss.n14419 9.3
R11311 vss.n14419 vss.n14418 9.3
R11312 vss.n14262 vss.n14261 9.3
R11313 vss.n14261 vss.n14260 9.3
R11314 vss.n13320 vss.n13319 9.3
R11315 vss.n14806 vss.n14805 9.3
R11316 vss.n14792 vss.n14791 9.3
R11317 vss.n14778 vss.n14777 9.3
R11318 vss.n14764 vss.n13321 9.3
R11319 vss.n14745 vss.n14744 9.3
R11320 vss.n14674 vss.n14673 9.3
R11321 vss.n14621 vss.n14620 9.3
R11322 vss.n14544 vss.n14543 9.3
R11323 vss.n14527 vss.n14526 9.3
R11324 vss.n14511 vss.n14510 9.3
R11325 vss.n14473 vss.n14472 9.3
R11326 vss.n14451 vss.n14181 9.3
R11327 vss.n14439 vss.n14213 9.3
R11328 vss.n14450 vss.n14449 9.3
R11329 vss.n13596 vss.n13595 9.3
R11330 vss.n13357 vss.n13356 9.3
R11331 vss.n14807 vss.n13277 9.3
R11332 vss.n14808 vss.n14807 9.3
R11333 vss.n14804 vss.n14803 9.3
R11334 vss.n14803 vss.n14802 9.3
R11335 vss.n14802 vss.n14801 9.3
R11336 vss.n14780 vss.n14779 9.3
R11337 vss.n14776 vss.n14775 9.3
R11338 vss.n14775 vss.n14774 9.3
R11339 vss.n14774 vss.n14773 9.3
R11340 vss.n14731 vss.n14730 9.3
R11341 vss.n13352 vss.n13351 9.3
R11342 vss.n13351 vss.n13350 9.3
R11343 vss.n14697 vss.n14696 9.3
R11344 vss.n14696 vss.n14695 9.3
R11345 vss.n14686 vss.n14685 9.3
R11346 vss.n13516 vss.n13515 9.3
R11347 vss.n13515 vss.n13514 9.3
R11348 vss.n14631 vss.n14630 9.3
R11349 vss.n14630 vss.n14629 9.3
R11350 vss.n14629 vss.n14628 9.3
R11351 vss.n14619 vss.n14618 9.3
R11352 vss.n14606 vss.n13544 9.3
R11353 vss.n13544 vss.n13543 9.3
R11354 vss.n13543 vss.n13542 9.3
R11355 vss.n14597 vss.n14596 9.3
R11356 vss.n14596 vss.n14595 9.3
R11357 vss.n14595 vss.n14594 9.3
R11358 vss.n14546 vss.n14545 9.3
R11359 vss.n14542 vss.n14541 9.3
R11360 vss.n14541 vss.n14540 9.3
R11361 vss.n14540 vss.n14539 9.3
R11362 vss.n14513 vss.n14512 9.3
R11363 vss.n14509 vss.n14508 9.3
R11364 vss.n14508 vss.n14507 9.3
R11365 vss.n14507 vss.n14506 9.3
R11366 vss.n14448 vss.n14447 9.3
R11367 vss.n14190 vss.n14189 9.3
R11368 vss.n14189 vss.n14188 9.3
R11369 vss.n14439 vss.n14212 9.3
R11370 vss.n14210 vss.n14209 9.3
R11371 vss.n14209 vss.n14208 9.3
R11372 vss.n14200 vss.n14199 9.3
R11373 vss.n14199 vss.n14198 9.3
R11374 vss.n14445 vss.n14444 9.3
R11375 vss.n14471 vss.n14470 9.3
R11376 vss.n14470 vss.n14469 9.3
R11377 vss.n14469 vss.n14468 9.3
R11378 vss.n14475 vss.n14474 9.3
R11379 vss.n14525 vss.n14524 9.3
R11380 vss.n14524 vss.n14523 9.3
R11381 vss.n14523 vss.n14522 9.3
R11382 vss.n14529 vss.n14528 9.3
R11383 vss.n14557 vss.n14556 9.3
R11384 vss.n14556 vss.n14555 9.3
R11385 vss.n14555 vss.n14554 9.3
R11386 vss.n14617 vss.n14616 9.3
R11387 vss.n14616 vss.n14615 9.3
R11388 vss.n14615 vss.n14614 9.3
R11389 vss.n13533 vss.n13532 9.3
R11390 vss.n13532 vss.n13531 9.3
R11391 vss.n14672 vss.n14671 9.3
R11392 vss.n14684 vss.n14683 9.3
R11393 vss.n14683 vss.n14682 9.3
R11394 vss.n14682 vss.n14681 9.3
R11395 vss.n14702 vss.n14701 9.3
R11396 vss.n13388 vss.n13387 9.3
R11397 vss.n13387 vss.n13386 9.3
R11398 vss.n13368 vss.n13367 9.3
R11399 vss.n13367 vss.n13366 9.3
R11400 vss.n14726 vss.n14725 9.3
R11401 vss.n14743 vss.n14742 9.3
R11402 vss.n14742 vss.n14741 9.3
R11403 vss.n14741 vss.n14740 9.3
R11404 vss.n14746 vss.n13322 9.3
R11405 vss.n14790 vss.n14789 9.3
R11406 vss.n14789 vss.n14788 9.3
R11407 vss.n14788 vss.n14787 9.3
R11408 vss.n14794 vss.n14793 9.3
R11409 vss.n13330 vss.n13329 9.3
R11410 vss.n13318 vss.n13317 9.3
R11411 vss.n13317 vss.n13316 9.3
R11412 vss.n13316 vss.n13315 9.3
R11413 vss.n14766 vss.n14765 9.3
R11414 vss.n14755 vss.n14754 9.3
R11415 vss.n14754 vss.n14753 9.3
R11416 vss.n14753 vss.n14752 9.3
R11417 vss.n13342 vss.n13341 9.3
R11418 vss.n13341 vss.n13340 9.3
R11419 vss.n14653 vss.n14652 9.3
R11420 vss.n13572 vss.n13571 9.3
R11421 vss.n13505 vss.n13504 9.3
R11422 vss.n14664 vss.n14663 9.3
R11423 vss.n14663 vss.n14662 9.3
R11424 vss.n14641 vss.n14640 9.3
R11425 vss.n14640 vss.n14639 9.3
R11426 vss.n13563 vss.n13562 9.3
R11427 vss.n13562 vss.n13561 9.3
R11428 vss.n13583 vss.n13582 9.3
R11429 vss.n13582 vss.n13581 9.3
R11430 vss.n14483 vss.n14482 9.3
R11431 vss.n14170 vss.n14169 9.3
R11432 vss.n14494 vss.n14493 9.3
R11433 vss.n14493 vss.n14492 9.3
R11434 vss.n14460 vss.n14459 9.3
R11435 vss.n14459 vss.n14458 9.3
R11436 vss.n14458 vss.n14457 9.3
R11437 vss.n14441 vss.n14440 9.3
R11438 vss.n14430 vss.n14429 9.3
R11439 vss.n14429 vss.n14428 9.3
R11440 vss.n14428 vss.n14427 9.3
R11441 vss.n15037 vss.n15036 9.3
R11442 vss.n15021 vss.n15020 9.3
R11443 vss.n14956 vss.n14955 9.3
R11444 vss.n14940 vss.n14939 9.3
R11445 vss.n14924 vss.n14923 9.3
R11446 vss.n13246 vss.n13245 9.3
R11447 vss.n13229 vss.n13228 9.3
R11448 vss.n13228 vss.n13227 9.3
R11449 vss.n13244 vss.n13243 9.3
R11450 vss.n13243 vss.n13242 9.3
R11451 vss.n13242 vss.n13241 9.3
R11452 vss.n13249 vss.n13248 9.3
R11453 vss.n14922 vss.n14921 9.3
R11454 vss.n14921 vss.n14920 9.3
R11455 vss.n14920 vss.n14919 9.3
R11456 vss.n14927 vss.n14926 9.3
R11457 vss.n14929 vss.n14928 9.3
R11458 vss.n14950 vss.n14949 9.3
R11459 vss.n14949 vss.n14948 9.3
R11460 vss.n14948 vss.n14947 9.3
R11461 vss.n14953 vss.n14952 9.3
R11462 vss.n14965 vss.n14964 9.3
R11463 vss.n14964 vss.n14963 9.3
R11464 vss.n14963 vss.n14962 9.3
R11465 vss.n13188 vss.n13187 9.3
R11466 vss.n12828 vss.n12827 9.3
R11467 vss.n15019 vss.n15018 9.3
R11468 vss.n15018 vss.n15017 9.3
R11469 vss.n15017 vss.n15016 9.3
R11470 vss.n15024 vss.n15023 9.3
R11471 vss.n15035 vss.n15034 9.3
R11472 vss.n15034 vss.n15033 9.3
R11473 vss.n15033 vss.n15032 9.3
R11474 vss.n15040 vss.n15039 9.3
R11475 vss.n13198 vss.n13197 9.3
R11476 vss.n13275 vss.n13274 9.3
R11477 vss.n13274 vss.n13273 9.3
R11478 vss.n13259 vss.n13258 9.3
R11479 vss.n13258 vss.n13257 9.3
R11480 vss.n14817 vss.n14816 9.3
R11481 vss.n14816 vss.n14815 9.3
R11482 vss.n12797 vss.n12796 9.3
R11483 vss.n13219 vss.n13218 9.3
R11484 vss.n14937 vss.n14935 9.3
R11485 vss.n13289 vss.n13288 9.3
R11486 vss.n13301 vss.n13300 9.3
R11487 vss.n13300 vss.n13299 9.3
R11488 vss.n12872 vss.n12871 9.3
R11489 vss.n12871 vss.n12870 9.3
R11490 vss.n12863 vss.n12862 9.3
R11491 vss.n12842 vss.n12841 9.3
R11492 vss.n12841 vss.n12840 9.3
R11493 vss.n14894 vss.n14893 9.3
R11494 vss.n14893 vss.n14892 9.3
R11495 vss.n14865 vss.n14864 9.3
R11496 vss.n14864 vss.n14863 9.3
R11497 vss.n14863 vss.n14862 9.3
R11498 vss.n14837 vss.n14836 9.3
R11499 vss.n14836 vss.n14835 9.3
R11500 vss.n14835 vss.n14834 9.3
R11501 vss.n14908 vss.n14907 9.3
R11502 vss.n14907 vss.n14906 9.3
R11503 vss.n14906 vss.n14905 9.3
R11504 vss.n14879 vss.n14878 9.3
R11505 vss.n14878 vss.n14877 9.3
R11506 vss.n12857 vss.n12856 9.3
R11507 vss.n12856 vss.n12855 9.3
R11508 vss.n12878 vss.n12877 9.3
R11509 vss.n12893 vss.n12892 9.3
R11510 vss.n12892 vss.n12891 9.3
R11511 vss.n3816 vss.n3815 9.3
R11512 vss.n3827 vss.n3826 9.3
R11513 vss.n3814 vss.n3813 9.3
R11514 vss.n3823 vss.n3822 9.3
R11515 vss.n3822 vss.n3821 9.3
R11516 vss.n3825 vss.n3824 9.3
R11517 vss.n3834 vss.n3833 9.3
R11518 vss.n3833 vss.n3832 9.3
R11519 vss.n3809 vss.n3808 9.3
R11520 vss.n3791 vss.n3790 9.3
R11521 vss.n3790 vss.n3789 9.3
R11522 vss.n3775 vss.n3774 9.3
R11523 vss.n3784 vss.n3783 9.3
R11524 vss.n3783 vss.n3782 9.3
R11525 vss.n3777 vss.n3776 9.3
R11526 vss.n3793 vss.n3792 9.3
R11527 vss.n3795 vss.n3794 9.3
R11528 vss.n3803 vss.n3802 9.3
R11529 vss.n3802 vss.n3801 9.3
R11530 vss.n3854 vss.n3853 9.3
R11531 vss.n3805 vss.n3804 9.3
R11532 vss.n3886 vss.n3885 9.3
R11533 vss.n3879 vss.n3878 9.3
R11534 vss.n3881 vss.n3880 9.3
R11535 vss.n3883 vss.n3882 9.3
R11536 vss.n3953 vss.n3952 9.3
R11537 vss.n3960 vss.n3959 9.3
R11538 vss.n3973 vss.n3972 9.3
R11539 vss.n3967 vss.n3966 9.3
R11540 vss.n3757 vss.n3756 9.3
R11541 vss.n3969 vss.n3968 9.3
R11542 vss.n3971 vss.n3970 9.3
R11543 vss.n3975 vss.n3974 9.3
R11544 vss.n3963 vss.n3962 9.3
R11545 vss.n3958 vss.n3957 9.3
R11546 vss.n3956 vss.n3955 9.3
R11547 vss.n3951 vss.n3950 9.3
R11548 vss.n3995 vss.n3994 9.3
R11549 vss.n3990 vss.n3989 9.3
R11550 vss.n3985 vss.n3984 9.3
R11551 vss.n3992 vss.n3991 9.3
R11552 vss.n3983 vss.n3982 9.3
R11553 vss.n3988 vss.n3987 9.3
R11554 vss.n3997 vss.n3996 9.3
R11555 vss.n3922 vss.n3921 9.3
R11556 vss.n3918 vss.n3917 9.3
R11557 vss.n3910 vss.n3909 9.3
R11558 vss.n3906 vss.n3905 9.3
R11559 vss.n3908 vss.n3907 9.3
R11560 vss.n3913 vss.n3912 9.3
R11561 vss.n3998 vss.n3934 9.3
R11562 vss.n3661 vss.n3660 9.3
R11563 vss.n3696 vss.n3695 9.3
R11564 vss.n3691 vss.n3654 9.3
R11565 vss.n3692 vss.n3691 9.3
R11566 vss.n3689 vss.n3688 9.3
R11567 vss.n3672 vss.n3669 9.3
R11568 vss.n3671 vss.n3670 9.3
R11569 vss.n3674 vss.n3673 9.3
R11570 vss.n3675 vss.n3674 9.3
R11571 vss.n3684 vss.n3666 9.3
R11572 vss.n3684 vss.n3683 9.3
R11573 vss.n3687 vss.n3686 9.3
R11574 vss.n3685 vss.n3664 9.3
R11575 vss.n3718 vss.n3710 9.3
R11576 vss.n3713 vss.n3711 9.3
R11577 vss.n3720 vss.n3719 9.3
R11578 vss.n3717 vss.n3716 9.3
R11579 vss.n3715 vss.n3714 9.3
R11580 vss.n3712 vss.n3636 9.3
R11581 vss.n3733 vss.n3724 9.3
R11582 vss.n3728 vss.n3725 9.3
R11583 vss.n3742 vss.n3635 9.3
R11584 vss.n3643 vss.n3634 9.3
R11585 vss.n3727 vss.n3726 9.3
R11586 vss.n3730 vss.n3729 9.3
R11587 vss.n3732 vss.n3731 9.3
R11588 vss.n3735 vss.n3734 9.3
R11589 vss.n3741 vss.n3740 9.3
R11590 vss.n3632 vss.n3631 9.3
R11591 vss.n3626 vss.n3614 9.3
R11592 vss.n3623 vss.n3622 9.3
R11593 vss.n3633 vss.n3613 9.3
R11594 vss.n3630 vss.n3629 9.3
R11595 vss.n3628 vss.n3627 9.3
R11596 vss.n3625 vss.n3624 9.3
R11597 vss.n3621 vss.n3620 9.3
R11598 vss.n3601 vss.n3595 9.3
R11599 vss.n3603 vss.n3602 9.3
R11600 vss.n3617 vss.n3616 9.3
R11601 vss.n3597 vss.n3591 9.3
R11602 vss.n3745 vss.n3597 9.3
R11603 vss.n3748 vss.n3747 9.3
R11604 vss.n3606 vss.n3605 9.3
R11605 vss.n5633 vss.n4240 9.3
R11606 vss.n5615 vss.n4250 9.3
R11607 vss.n4259 vss.n4258 9.3
R11608 vss.n4267 vss.n4257 9.3
R11609 vss.n5594 vss.n4266 9.3
R11610 vss.n5584 vss.n5583 9.3
R11611 vss.n4279 vss.n4276 9.3
R11612 vss.n5571 vss.n4286 9.3
R11613 vss.n5549 vss.n5548 9.3
R11614 vss.n5544 vss.n4302 9.3
R11615 vss.n5534 vss.n4314 9.3
R11616 vss.n4323 vss.n4321 9.3
R11617 vss.n5521 vss.n4324 9.3
R11618 vss.n5511 vss.n4333 9.3
R11619 vss.n4342 vss.n4340 9.3
R11620 vss.n5491 vss.n5490 9.3
R11621 vss.n4354 vss.n4352 9.3
R11622 vss.n5478 vss.n4364 9.3
R11623 vss.n5468 vss.n5467 9.3
R11624 vss.n4376 vss.n4373 9.3
R11625 vss.n5455 vss.n4383 9.3
R11626 vss.n5445 vss.n5444 9.3
R11627 vss.n5431 vss.n4405 9.3
R11628 vss.n5421 vss.n4414 9.3
R11629 vss.n4423 vss.n4421 9.3
R11630 vss.n5408 vss.n4424 9.3
R11631 vss.n5398 vss.n4433 9.3
R11632 vss.n4442 vss.n4440 9.3
R11633 vss.n5385 vss.n4443 9.3
R11634 vss.n4455 vss.n4453 9.3
R11635 vss.n5365 vss.n4464 9.3
R11636 vss.n5355 vss.n5354 9.3
R11637 vss.n4476 vss.n4473 9.3
R11638 vss.n5342 vss.n4483 9.3
R11639 vss.n5332 vss.n5331 9.3
R11640 vss.n4495 vss.n4492 9.3
R11641 vss.n5308 vss.n5307 9.3
R11642 vss.n5303 vss.n4515 9.3
R11643 vss.n5293 vss.n4527 9.3
R11644 vss.n4536 vss.n4534 9.3
R11645 vss.n5280 vss.n4537 9.3
R11646 vss.n5270 vss.n4546 9.3
R11647 vss.n4555 vss.n4553 9.3
R11648 vss.n5250 vss.n5249 9.3
R11649 vss.n4567 vss.n4565 9.3
R11650 vss.n5237 vss.n4577 9.3
R11651 vss.n5227 vss.n5226 9.3
R11652 vss.n4589 vss.n4586 9.3
R11653 vss.n5214 vss.n4596 9.3
R11654 vss.n5204 vss.n5203 9.3
R11655 vss.n5190 vss.n4618 9.3
R11656 vss.n5180 vss.n4627 9.3
R11657 vss.n4636 vss.n4634 9.3
R11658 vss.n5167 vss.n4637 9.3
R11659 vss.n5157 vss.n4646 9.3
R11660 vss.n4655 vss.n4653 9.3
R11661 vss.n5144 vss.n4656 9.3
R11662 vss.n4668 vss.n4666 9.3
R11663 vss.n5124 vss.n4677 9.3
R11664 vss.n5114 vss.n5113 9.3
R11665 vss.n4689 vss.n4686 9.3
R11666 vss.n5101 vss.n4696 9.3
R11667 vss.n5091 vss.n5090 9.3
R11668 vss.n4708 vss.n4705 9.3
R11669 vss.n5067 vss.n5066 9.3
R11670 vss.n5062 vss.n4728 9.3
R11671 vss.n5052 vss.n4740 9.3
R11672 vss.n4749 vss.n4747 9.3
R11673 vss.n5039 vss.n4750 9.3
R11674 vss.n5029 vss.n4759 9.3
R11675 vss.n4768 vss.n4766 9.3
R11676 vss.n5009 vss.n5008 9.3
R11677 vss.n4780 vss.n4778 9.3
R11678 vss.n4996 vss.n4790 9.3
R11679 vss.n4986 vss.n4985 9.3
R11680 vss.n4802 vss.n4799 9.3
R11681 vss.n4973 vss.n4809 9.3
R11682 vss.n4963 vss.n4962 9.3
R11683 vss.n4949 vss.n4831 9.3
R11684 vss.n4939 vss.n4840 9.3
R11685 vss.n4849 vss.n4847 9.3
R11686 vss.n4926 vss.n4850 9.3
R11687 vss.n4916 vss.n4859 9.3
R11688 vss.n4868 vss.n4866 9.3
R11689 vss.n4903 vss.n4869 9.3
R11690 vss.n4907 vss.n4906 9.3
R11691 vss.n4908 vss.n4907 9.3
R11692 vss.n4909 vss.n4908 9.3
R11693 vss.n4865 vss.n4860 9.3
R11694 vss.n4925 vss.n4853 9.3
R11695 vss.n4925 vss.n4924 9.3
R11696 vss.n4924 vss.n4923 9.3
R11697 vss.n4928 vss.n4927 9.3
R11698 vss.n4938 vss.n4937 9.3
R11699 vss.n4937 vss.n4839 9.3
R11700 vss.n4839 vss.n4838 9.3
R11701 vss.n4941 vss.n4940 9.3
R11702 vss.n4953 vss.n4952 9.3
R11703 vss.n4954 vss.n4953 9.3
R11704 vss.n4955 vss.n4954 9.3
R11705 vss.n4961 vss.n4817 9.3
R11706 vss.n4811 vss.n4810 9.3
R11707 vss.n4995 vss.n4994 9.3
R11708 vss.n5007 vss.n4777 9.3
R11709 vss.n5028 vss.n5027 9.3
R11710 vss.n5027 vss.n4758 9.3
R11711 vss.n4758 vss.n4757 9.3
R11712 vss.n5031 vss.n5030 9.3
R11713 vss.n5043 vss.n5042 9.3
R11714 vss.n5044 vss.n5043 9.3
R11715 vss.n5045 vss.n5044 9.3
R11716 vss.n4746 vss.n4741 9.3
R11717 vss.n5061 vss.n4731 9.3
R11718 vss.n5061 vss.n5060 9.3
R11719 vss.n5060 vss.n5059 9.3
R11720 vss.n5064 vss.n5063 9.3
R11721 vss.n5076 vss.n5075 9.3
R11722 vss.n5075 vss.n5074 9.3
R11723 vss.n5074 vss.n5073 9.3
R11724 vss.n4717 vss.n4716 9.3
R11725 vss.n5100 vss.n5099 9.3
R11726 vss.n5112 vss.n4685 9.3
R11727 vss.n4679 vss.n4678 9.3
R11728 vss.n5148 vss.n5147 9.3
R11729 vss.n5149 vss.n5148 9.3
R11730 vss.n5150 vss.n5149 9.3
R11731 vss.n4652 vss.n4647 9.3
R11732 vss.n5166 vss.n4640 9.3
R11733 vss.n5166 vss.n5165 9.3
R11734 vss.n5165 vss.n5164 9.3
R11735 vss.n5169 vss.n5168 9.3
R11736 vss.n5179 vss.n5178 9.3
R11737 vss.n5178 vss.n4626 9.3
R11738 vss.n4626 vss.n4625 9.3
R11739 vss.n5182 vss.n5181 9.3
R11740 vss.n5194 vss.n5193 9.3
R11741 vss.n5195 vss.n5194 9.3
R11742 vss.n5196 vss.n5195 9.3
R11743 vss.n5202 vss.n4604 9.3
R11744 vss.n4598 vss.n4597 9.3
R11745 vss.n5236 vss.n5235 9.3
R11746 vss.n5248 vss.n4564 9.3
R11747 vss.n5269 vss.n5268 9.3
R11748 vss.n5268 vss.n4545 9.3
R11749 vss.n4545 vss.n4544 9.3
R11750 vss.n5272 vss.n5271 9.3
R11751 vss.n5284 vss.n5283 9.3
R11752 vss.n5285 vss.n5284 9.3
R11753 vss.n5286 vss.n5285 9.3
R11754 vss.n4533 vss.n4528 9.3
R11755 vss.n5302 vss.n4518 9.3
R11756 vss.n5302 vss.n5301 9.3
R11757 vss.n5301 vss.n5300 9.3
R11758 vss.n5305 vss.n5304 9.3
R11759 vss.n5317 vss.n5316 9.3
R11760 vss.n5316 vss.n5315 9.3
R11761 vss.n5315 vss.n5314 9.3
R11762 vss.n4504 vss.n4503 9.3
R11763 vss.n5341 vss.n5340 9.3
R11764 vss.n5353 vss.n4472 9.3
R11765 vss.n4466 vss.n4465 9.3
R11766 vss.n5389 vss.n5388 9.3
R11767 vss.n5390 vss.n5389 9.3
R11768 vss.n5391 vss.n5390 9.3
R11769 vss.n4439 vss.n4434 9.3
R11770 vss.n5407 vss.n4427 9.3
R11771 vss.n5407 vss.n5406 9.3
R11772 vss.n5406 vss.n5405 9.3
R11773 vss.n5410 vss.n5409 9.3
R11774 vss.n5420 vss.n5419 9.3
R11775 vss.n5419 vss.n4413 9.3
R11776 vss.n4413 vss.n4412 9.3
R11777 vss.n5423 vss.n5422 9.3
R11778 vss.n5435 vss.n5434 9.3
R11779 vss.n5436 vss.n5435 9.3
R11780 vss.n5437 vss.n5436 9.3
R11781 vss.n5443 vss.n4391 9.3
R11782 vss.n4385 vss.n4384 9.3
R11783 vss.n5477 vss.n5476 9.3
R11784 vss.n5489 vss.n4351 9.3
R11785 vss.n5510 vss.n5509 9.3
R11786 vss.n5509 vss.n4332 9.3
R11787 vss.n4332 vss.n4331 9.3
R11788 vss.n5513 vss.n5512 9.3
R11789 vss.n5525 vss.n5524 9.3
R11790 vss.n5526 vss.n5525 9.3
R11791 vss.n5527 vss.n5526 9.3
R11792 vss.n4320 vss.n4315 9.3
R11793 vss.n5543 vss.n4305 9.3
R11794 vss.n5543 vss.n5542 9.3
R11795 vss.n5542 vss.n5541 9.3
R11796 vss.n5546 vss.n5545 9.3
R11797 vss.n5558 vss.n5557 9.3
R11798 vss.n5557 vss.n5556 9.3
R11799 vss.n5556 vss.n5555 9.3
R11800 vss.n5570 vss.n5569 9.3
R11801 vss.n5582 vss.n4275 9.3
R11802 vss.n4269 vss.n4268 9.3
R11803 vss.n5614 vss.n5613 9.3
R11804 vss.n4239 vss.n4236 9.3
R11805 vss.n5635 vss.n5634 9.3
R11806 vss.n5632 vss.n5631 9.3
R11807 vss.n5631 vss.n5630 9.3
R11808 vss.n5630 vss.n5629 9.3
R11809 vss.n5617 vss.n5616 9.3
R11810 vss.n5618 vss.n5617 9.3
R11811 vss.n5619 vss.n5618 9.3
R11812 vss.n4252 vss.n4251 9.3
R11813 vss.n4253 vss.n4252 9.3
R11814 vss.n5608 vss.n4253 9.3
R11815 vss.n4260 vss.n4256 9.3
R11816 vss.n5603 vss.n4261 9.3
R11817 vss.n5603 vss.n5602 9.3
R11818 vss.n5602 vss.n5601 9.3
R11819 vss.n5596 vss.n5595 9.3
R11820 vss.n5596 vss.n4264 9.3
R11821 vss.n4264 vss.n4263 9.3
R11822 vss.n5593 vss.n5592 9.3
R11823 vss.n5585 vss.n4270 9.3
R11824 vss.n5586 vss.n5585 9.3
R11825 vss.n5587 vss.n5586 9.3
R11826 vss.n5581 vss.n5580 9.3
R11827 vss.n5580 vss.n5579 9.3
R11828 vss.n5579 vss.n5578 9.3
R11829 vss.n4288 vss.n4287 9.3
R11830 vss.n5573 vss.n5572 9.3
R11831 vss.n5573 vss.n4284 9.3
R11832 vss.n4284 vss.n4283 9.3
R11833 vss.n5562 vss.n4289 9.3
R11834 vss.n5563 vss.n5562 9.3
R11835 vss.n5564 vss.n5563 9.3
R11836 vss.n5550 vss.n4296 9.3
R11837 vss.n5547 vss.n4301 9.3
R11838 vss.n4301 vss.n4300 9.3
R11839 vss.n4300 vss.n4299 9.3
R11840 vss.n5536 vss.n5535 9.3
R11841 vss.n5533 vss.n5532 9.3
R11842 vss.n5532 vss.n4313 9.3
R11843 vss.n4313 vss.n4312 9.3
R11844 vss.n5523 vss.n5522 9.3
R11845 vss.n5520 vss.n4327 9.3
R11846 vss.n5520 vss.n5519 9.3
R11847 vss.n5519 vss.n5518 9.3
R11848 vss.n4339 vss.n4334 9.3
R11849 vss.n5502 vss.n5501 9.3
R11850 vss.n5503 vss.n5502 9.3
R11851 vss.n5504 vss.n5503 9.3
R11852 vss.n5492 vss.n4343 9.3
R11853 vss.n5492 vss.n4350 9.3
R11854 vss.n4350 vss.n4349 9.3
R11855 vss.n5488 vss.n5487 9.3
R11856 vss.n5487 vss.n5486 9.3
R11857 vss.n5486 vss.n5485 9.3
R11858 vss.n4366 vss.n4365 9.3
R11859 vss.n5480 vss.n5479 9.3
R11860 vss.n5480 vss.n4362 9.3
R11861 vss.n4362 vss.n4361 9.3
R11862 vss.n5469 vss.n4367 9.3
R11863 vss.n5470 vss.n5469 9.3
R11864 vss.n5471 vss.n5470 9.3
R11865 vss.n5466 vss.n4372 9.3
R11866 vss.n5465 vss.n5464 9.3
R11867 vss.n5464 vss.n5463 9.3
R11868 vss.n5463 vss.n5462 9.3
R11869 vss.n5457 vss.n5456 9.3
R11870 vss.n5457 vss.n4381 9.3
R11871 vss.n4381 vss.n4380 9.3
R11872 vss.n5454 vss.n5453 9.3
R11873 vss.n5446 vss.n4386 9.3
R11874 vss.n5447 vss.n5446 9.3
R11875 vss.n5448 vss.n5447 9.3
R11876 vss.n5442 vss.n5441 9.3
R11877 vss.n5441 vss.n5440 9.3
R11878 vss.n5440 vss.n5439 9.3
R11879 vss.n5433 vss.n5432 9.3
R11880 vss.n5430 vss.n4408 9.3
R11881 vss.n5430 vss.n5429 9.3
R11882 vss.n5429 vss.n5428 9.3
R11883 vss.n4420 vss.n4415 9.3
R11884 vss.n5412 vss.n5411 9.3
R11885 vss.n5413 vss.n5412 9.3
R11886 vss.n5414 vss.n5413 9.3
R11887 vss.n5400 vss.n5399 9.3
R11888 vss.n5397 vss.n5396 9.3
R11889 vss.n5396 vss.n4432 9.3
R11890 vss.n4432 vss.n4431 9.3
R11891 vss.n5387 vss.n5386 9.3
R11892 vss.n5384 vss.n4446 9.3
R11893 vss.n5384 vss.n5383 9.3
R11894 vss.n5383 vss.n5382 9.3
R11895 vss.n5375 vss.n5374 9.3
R11896 vss.n5374 vss.n5373 9.3
R11897 vss.n5373 vss.n5372 9.3
R11898 vss.n5367 vss.n5366 9.3
R11899 vss.n5367 vss.n4462 9.3
R11900 vss.n4462 vss.n4461 9.3
R11901 vss.n5364 vss.n5363 9.3
R11902 vss.n5356 vss.n4467 9.3
R11903 vss.n5357 vss.n5356 9.3
R11904 vss.n5358 vss.n5357 9.3
R11905 vss.n5352 vss.n5351 9.3
R11906 vss.n5351 vss.n5350 9.3
R11907 vss.n5350 vss.n5349 9.3
R11908 vss.n4485 vss.n4484 9.3
R11909 vss.n5344 vss.n5343 9.3
R11910 vss.n5344 vss.n4481 9.3
R11911 vss.n4481 vss.n4480 9.3
R11912 vss.n5333 vss.n4486 9.3
R11913 vss.n5334 vss.n5333 9.3
R11914 vss.n5335 vss.n5334 9.3
R11915 vss.n5330 vss.n4491 9.3
R11916 vss.n5329 vss.n5328 9.3
R11917 vss.n5328 vss.n5327 9.3
R11918 vss.n5327 vss.n5326 9.3
R11919 vss.n5321 vss.n5320 9.3
R11920 vss.n5321 vss.n4500 9.3
R11921 vss.n4500 vss.n4499 9.3
R11922 vss.n5309 vss.n4506 9.3
R11923 vss.n5306 vss.n4514 9.3
R11924 vss.n4514 vss.n4513 9.3
R11925 vss.n4513 vss.n4512 9.3
R11926 vss.n5295 vss.n5294 9.3
R11927 vss.n5292 vss.n5291 9.3
R11928 vss.n5291 vss.n4526 9.3
R11929 vss.n4526 vss.n4525 9.3
R11930 vss.n5282 vss.n5281 9.3
R11931 vss.n5279 vss.n4540 9.3
R11932 vss.n5279 vss.n5278 9.3
R11933 vss.n5278 vss.n5277 9.3
R11934 vss.n4552 vss.n4547 9.3
R11935 vss.n5261 vss.n5260 9.3
R11936 vss.n5262 vss.n5261 9.3
R11937 vss.n5263 vss.n5262 9.3
R11938 vss.n5251 vss.n4556 9.3
R11939 vss.n5251 vss.n4563 9.3
R11940 vss.n4563 vss.n4562 9.3
R11941 vss.n5247 vss.n5246 9.3
R11942 vss.n5246 vss.n5245 9.3
R11943 vss.n5245 vss.n5244 9.3
R11944 vss.n4579 vss.n4578 9.3
R11945 vss.n5239 vss.n5238 9.3
R11946 vss.n5239 vss.n4575 9.3
R11947 vss.n4575 vss.n4574 9.3
R11948 vss.n5228 vss.n4580 9.3
R11949 vss.n5229 vss.n5228 9.3
R11950 vss.n5230 vss.n5229 9.3
R11951 vss.n5225 vss.n4585 9.3
R11952 vss.n5224 vss.n5223 9.3
R11953 vss.n5223 vss.n5222 9.3
R11954 vss.n5222 vss.n5221 9.3
R11955 vss.n5216 vss.n5215 9.3
R11956 vss.n5216 vss.n4594 9.3
R11957 vss.n4594 vss.n4593 9.3
R11958 vss.n5213 vss.n5212 9.3
R11959 vss.n5205 vss.n4599 9.3
R11960 vss.n5206 vss.n5205 9.3
R11961 vss.n5207 vss.n5206 9.3
R11962 vss.n5201 vss.n5200 9.3
R11963 vss.n5200 vss.n5199 9.3
R11964 vss.n5199 vss.n5198 9.3
R11965 vss.n5192 vss.n5191 9.3
R11966 vss.n5189 vss.n4621 9.3
R11967 vss.n5189 vss.n5188 9.3
R11968 vss.n5188 vss.n5187 9.3
R11969 vss.n4633 vss.n4628 9.3
R11970 vss.n5171 vss.n5170 9.3
R11971 vss.n5172 vss.n5171 9.3
R11972 vss.n5173 vss.n5172 9.3
R11973 vss.n5159 vss.n5158 9.3
R11974 vss.n5156 vss.n5155 9.3
R11975 vss.n5155 vss.n4645 9.3
R11976 vss.n4645 vss.n4644 9.3
R11977 vss.n5146 vss.n5145 9.3
R11978 vss.n5143 vss.n4659 9.3
R11979 vss.n5143 vss.n5142 9.3
R11980 vss.n5142 vss.n5141 9.3
R11981 vss.n5134 vss.n5133 9.3
R11982 vss.n5133 vss.n5132 9.3
R11983 vss.n5132 vss.n5131 9.3
R11984 vss.n5126 vss.n5125 9.3
R11985 vss.n5126 vss.n4675 9.3
R11986 vss.n4675 vss.n4674 9.3
R11987 vss.n5123 vss.n5122 9.3
R11988 vss.n5115 vss.n4680 9.3
R11989 vss.n5116 vss.n5115 9.3
R11990 vss.n5117 vss.n5116 9.3
R11991 vss.n5111 vss.n5110 9.3
R11992 vss.n5110 vss.n5109 9.3
R11993 vss.n5109 vss.n5108 9.3
R11994 vss.n4698 vss.n4697 9.3
R11995 vss.n5103 vss.n5102 9.3
R11996 vss.n5103 vss.n4694 9.3
R11997 vss.n4694 vss.n4693 9.3
R11998 vss.n5092 vss.n4699 9.3
R11999 vss.n5093 vss.n5092 9.3
R12000 vss.n5094 vss.n5093 9.3
R12001 vss.n5089 vss.n4704 9.3
R12002 vss.n5088 vss.n5087 9.3
R12003 vss.n5087 vss.n5086 9.3
R12004 vss.n5086 vss.n5085 9.3
R12005 vss.n5080 vss.n5079 9.3
R12006 vss.n5080 vss.n4713 9.3
R12007 vss.n4713 vss.n4712 9.3
R12008 vss.n5068 vss.n4719 9.3
R12009 vss.n5065 vss.n4727 9.3
R12010 vss.n4727 vss.n4726 9.3
R12011 vss.n4726 vss.n4725 9.3
R12012 vss.n5054 vss.n5053 9.3
R12013 vss.n5051 vss.n5050 9.3
R12014 vss.n5050 vss.n4739 9.3
R12015 vss.n4739 vss.n4738 9.3
R12016 vss.n5041 vss.n5040 9.3
R12017 vss.n5038 vss.n4753 9.3
R12018 vss.n5038 vss.n5037 9.3
R12019 vss.n5037 vss.n5036 9.3
R12020 vss.n4765 vss.n4760 9.3
R12021 vss.n5020 vss.n5019 9.3
R12022 vss.n5021 vss.n5020 9.3
R12023 vss.n5022 vss.n5021 9.3
R12024 vss.n5010 vss.n4769 9.3
R12025 vss.n5010 vss.n4776 9.3
R12026 vss.n4776 vss.n4775 9.3
R12027 vss.n5006 vss.n5005 9.3
R12028 vss.n5005 vss.n5004 9.3
R12029 vss.n5004 vss.n5003 9.3
R12030 vss.n4792 vss.n4791 9.3
R12031 vss.n4998 vss.n4997 9.3
R12032 vss.n4998 vss.n4788 9.3
R12033 vss.n4788 vss.n4787 9.3
R12034 vss.n4987 vss.n4793 9.3
R12035 vss.n4988 vss.n4987 9.3
R12036 vss.n4989 vss.n4988 9.3
R12037 vss.n4984 vss.n4798 9.3
R12038 vss.n4983 vss.n4982 9.3
R12039 vss.n4982 vss.n4981 9.3
R12040 vss.n4981 vss.n4980 9.3
R12041 vss.n4975 vss.n4974 9.3
R12042 vss.n4975 vss.n4807 9.3
R12043 vss.n4807 vss.n4806 9.3
R12044 vss.n4972 vss.n4971 9.3
R12045 vss.n4964 vss.n4812 9.3
R12046 vss.n4965 vss.n4964 9.3
R12047 vss.n4966 vss.n4965 9.3
R12048 vss.n4960 vss.n4959 9.3
R12049 vss.n4959 vss.n4958 9.3
R12050 vss.n4958 vss.n4957 9.3
R12051 vss.n4951 vss.n4950 9.3
R12052 vss.n4948 vss.n4834 9.3
R12053 vss.n4948 vss.n4947 9.3
R12054 vss.n4947 vss.n4946 9.3
R12055 vss.n4846 vss.n4841 9.3
R12056 vss.n4930 vss.n4929 9.3
R12057 vss.n4931 vss.n4930 9.3
R12058 vss.n4932 vss.n4931 9.3
R12059 vss.n4918 vss.n4917 9.3
R12060 vss.n4915 vss.n4914 9.3
R12061 vss.n4914 vss.n4858 9.3
R12062 vss.n4858 vss.n4857 9.3
R12063 vss.n4905 vss.n4904 9.3
R12064 vss.n4902 vss.n4872 9.3
R12065 vss.n4902 vss.n4901 9.3
R12066 vss.n4901 vss.n4900 9.3
R12067 vss.n4881 vss.n4879 9.3
R12068 vss.n4883 vss.n4233 9.3
R12069 vss.n4893 vss.n4892 9.3
R12070 vss.n4892 vss.n4891 9.3
R12071 vss.n4891 vss.n4890 9.3
R12072 vss.n5640 vss.n6 9.3
R12073 vss.n4201 vss.n4196 9.3
R12074 vss.n6977 vss.n6976 9.3
R12075 vss.n4200 vss.n4199 9.3
R12076 vss.n6978 vss.n4191 9.3
R12077 vss.n6204 vss.n6203 9.3
R12078 vss.n6214 vss.n6202 9.3
R12079 vss.n6899 vss.n4232 9.3
R12080 vss.n5656 vss.n5655 9.3
R12081 vss.n5664 vss.n5653 9.3
R12082 vss.n6871 vss.n5663 9.3
R12083 vss.n6861 vss.n6860 9.3
R12084 vss.n5676 vss.n5673 9.3
R12085 vss.n6848 vss.n5683 9.3
R12086 vss.n6838 vss.n6837 9.3
R12087 vss.n6824 vss.n5705 9.3
R12088 vss.n6814 vss.n5714 9.3
R12089 vss.n5723 vss.n5721 9.3
R12090 vss.n6801 vss.n5724 9.3
R12091 vss.n6791 vss.n5733 9.3
R12092 vss.n5742 vss.n5740 9.3
R12093 vss.n6778 vss.n5743 9.3
R12094 vss.n6761 vss.n5757 9.3
R12095 vss.n5766 vss.n5765 9.3
R12096 vss.n5774 vss.n5764 9.3
R12097 vss.n6740 vss.n5773 9.3
R12098 vss.n6730 vss.n6729 9.3
R12099 vss.n5786 vss.n5783 9.3
R12100 vss.n6717 vss.n5793 9.3
R12101 vss.n6695 vss.n6694 9.3
R12102 vss.n6690 vss.n5809 9.3
R12103 vss.n6680 vss.n5821 9.3
R12104 vss.n5830 vss.n5828 9.3
R12105 vss.n6667 vss.n5831 9.3
R12106 vss.n6657 vss.n5840 9.3
R12107 vss.n5849 vss.n5847 9.3
R12108 vss.n6637 vss.n6636 9.3
R12109 vss.n5861 vss.n5859 9.3
R12110 vss.n6624 vss.n5871 9.3
R12111 vss.n6614 vss.n6613 9.3
R12112 vss.n5883 vss.n5880 9.3
R12113 vss.n6601 vss.n5890 9.3
R12114 vss.n6591 vss.n6590 9.3
R12115 vss.n6577 vss.n5912 9.3
R12116 vss.n6567 vss.n5921 9.3
R12117 vss.n5930 vss.n5928 9.3
R12118 vss.n6554 vss.n5931 9.3
R12119 vss.n6544 vss.n5940 9.3
R12120 vss.n5949 vss.n5947 9.3
R12121 vss.n6531 vss.n5950 9.3
R12122 vss.n6514 vss.n5964 9.3
R12123 vss.n5973 vss.n5972 9.3
R12124 vss.n5981 vss.n5971 9.3
R12125 vss.n6493 vss.n5980 9.3
R12126 vss.n6483 vss.n6482 9.3
R12127 vss.n5993 vss.n5990 9.3
R12128 vss.n6470 vss.n6000 9.3
R12129 vss.n6448 vss.n6447 9.3
R12130 vss.n6443 vss.n6016 9.3
R12131 vss.n6433 vss.n6028 9.3
R12132 vss.n6037 vss.n6035 9.3
R12133 vss.n6420 vss.n6038 9.3
R12134 vss.n6410 vss.n6047 9.3
R12135 vss.n6056 vss.n6054 9.3
R12136 vss.n6390 vss.n6389 9.3
R12137 vss.n6068 vss.n6066 9.3
R12138 vss.n6377 vss.n6078 9.3
R12139 vss.n6367 vss.n6366 9.3
R12140 vss.n6090 vss.n6087 9.3
R12141 vss.n6354 vss.n6097 9.3
R12142 vss.n6344 vss.n6343 9.3
R12143 vss.n6330 vss.n6119 9.3
R12144 vss.n6320 vss.n6128 9.3
R12145 vss.n6137 vss.n6135 9.3
R12146 vss.n6307 vss.n6138 9.3
R12147 vss.n6297 vss.n6147 9.3
R12148 vss.n6156 vss.n6154 9.3
R12149 vss.n6284 vss.n6157 9.3
R12150 vss.n6267 vss.n6171 9.3
R12151 vss.n6180 vss.n6179 9.3
R12152 vss.n6188 vss.n6178 9.3
R12153 vss.n6246 vss.n6187 9.3
R12154 vss.n6236 vss.n6235 9.3
R12155 vss.n6245 vss.n6244 9.3
R12156 vss.n6181 vss.n6177 9.3
R12157 vss.n6286 vss.n6285 9.3
R12158 vss.n6299 vss.n6298 9.3
R12159 vss.n6134 vss.n6129 9.3
R12160 vss.n6332 vss.n6331 9.3
R12161 vss.n6353 vss.n6352 9.3
R12162 vss.n6365 vss.n6086 9.3
R12163 vss.n6080 vss.n6079 9.3
R12164 vss.n6053 vss.n6048 9.3
R12165 vss.n6422 vss.n6421 9.3
R12166 vss.n6435 vss.n6434 9.3
R12167 vss.n6449 vss.n6009 9.3
R12168 vss.n6002 vss.n6001 9.3
R12169 vss.n6492 vss.n6491 9.3
R12170 vss.n5974 vss.n5970 9.3
R12171 vss.n6533 vss.n6532 9.3
R12172 vss.n6546 vss.n6545 9.3
R12173 vss.n5927 vss.n5922 9.3
R12174 vss.n6579 vss.n6578 9.3
R12175 vss.n6600 vss.n6599 9.3
R12176 vss.n6612 vss.n5879 9.3
R12177 vss.n5873 vss.n5872 9.3
R12178 vss.n5846 vss.n5841 9.3
R12179 vss.n6669 vss.n6668 9.3
R12180 vss.n6682 vss.n6681 9.3
R12181 vss.n6696 vss.n5803 9.3
R12182 vss.n5795 vss.n5794 9.3
R12183 vss.n6739 vss.n6738 9.3
R12184 vss.n5767 vss.n5763 9.3
R12185 vss.n6780 vss.n6779 9.3
R12186 vss.n6793 vss.n6792 9.3
R12187 vss.n5720 vss.n5715 9.3
R12188 vss.n6826 vss.n6825 9.3
R12189 vss.n6847 vss.n6846 9.3
R12190 vss.n6859 vss.n5672 9.3
R12191 vss.n5666 vss.n5665 9.3
R12192 vss.n6901 vss.n6900 9.3
R12193 vss.n5657 vss.n5652 9.3
R12194 vss.n6870 vss.n6869 9.3
R12195 vss.n5685 vss.n5684 9.3
R12196 vss.n6836 vss.n5691 9.3
R12197 vss.n6816 vss.n6815 9.3
R12198 vss.n6803 vss.n6802 9.3
R12199 vss.n5739 vss.n5734 9.3
R12200 vss.n6760 vss.n6759 9.3
R12201 vss.n5776 vss.n5775 9.3
R12202 vss.n6728 vss.n5782 9.3
R12203 vss.n6716 vss.n6715 9.3
R12204 vss.n6692 vss.n6691 9.3
R12205 vss.n5827 vss.n5822 9.3
R12206 vss.n6659 vss.n6658 9.3
R12207 vss.n6635 vss.n5858 9.3
R12208 vss.n6623 vss.n6622 9.3
R12209 vss.n5892 vss.n5891 9.3
R12210 vss.n6589 vss.n5898 9.3
R12211 vss.n6569 vss.n6568 9.3
R12212 vss.n6556 vss.n6555 9.3
R12213 vss.n5946 vss.n5941 9.3
R12214 vss.n6513 vss.n6512 9.3
R12215 vss.n5983 vss.n5982 9.3
R12216 vss.n6481 vss.n5989 9.3
R12217 vss.n6469 vss.n6468 9.3
R12218 vss.n6445 vss.n6444 9.3
R12219 vss.n6034 vss.n6029 9.3
R12220 vss.n6412 vss.n6411 9.3
R12221 vss.n6388 vss.n6065 9.3
R12222 vss.n6376 vss.n6375 9.3
R12223 vss.n6099 vss.n6098 9.3
R12224 vss.n6342 vss.n6105 9.3
R12225 vss.n6322 vss.n6321 9.3
R12226 vss.n6309 vss.n6308 9.3
R12227 vss.n6153 vss.n6148 9.3
R12228 vss.n6266 vss.n6265 9.3
R12229 vss.n6190 vss.n6189 9.3
R12230 vss.n6234 vss.n6196 9.3
R12231 vss.n6932 vss.n4215 9.3
R12232 vss.n6937 vss.n6936 9.3
R12233 vss.n6942 vss.n4211 9.3
R12234 vss.n6969 vss.n6968 9.3
R12235 vss.n6968 vss.n6967 9.3
R12236 vss.n6967 vss.n6966 9.3
R12237 vss.n6964 vss.n6963 9.3
R12238 vss.n6958 vss.n4206 9.3
R12239 vss.n6953 vss.n6952 9.3
R12240 vss.n6947 vss.n4209 9.3
R12241 vss.n4223 vss.n4217 9.3
R12242 vss.n6911 vss.n6910 9.3
R12243 vss.n6283 vss.n6160 9.3
R12244 vss.n6283 vss.n6282 9.3
R12245 vss.n6282 vss.n6281 9.3
R12246 vss.n6296 vss.n6295 9.3
R12247 vss.n6295 vss.n6146 9.3
R12248 vss.n6146 vss.n6145 9.3
R12249 vss.n6311 vss.n6310 9.3
R12250 vss.n6312 vss.n6311 9.3
R12251 vss.n6313 vss.n6312 9.3
R12252 vss.n6329 vss.n6122 9.3
R12253 vss.n6329 vss.n6328 9.3
R12254 vss.n6328 vss.n6327 9.3
R12255 vss.n6401 vss.n6400 9.3
R12256 vss.n6402 vss.n6401 9.3
R12257 vss.n6403 vss.n6402 9.3
R12258 vss.n6419 vss.n6041 9.3
R12259 vss.n6419 vss.n6418 9.3
R12260 vss.n6418 vss.n6417 9.3
R12261 vss.n6432 vss.n6431 9.3
R12262 vss.n6431 vss.n6027 9.3
R12263 vss.n6027 vss.n6026 9.3
R12264 vss.n6446 vss.n6015 9.3
R12265 vss.n6015 vss.n6014 9.3
R12266 vss.n6014 vss.n6013 9.3
R12267 vss.n6530 vss.n5953 9.3
R12268 vss.n6530 vss.n6529 9.3
R12269 vss.n6529 vss.n6528 9.3
R12270 vss.n6543 vss.n6542 9.3
R12271 vss.n6542 vss.n5939 9.3
R12272 vss.n5939 vss.n5938 9.3
R12273 vss.n6558 vss.n6557 9.3
R12274 vss.n6559 vss.n6558 9.3
R12275 vss.n6560 vss.n6559 9.3
R12276 vss.n6576 vss.n5915 9.3
R12277 vss.n6576 vss.n6575 9.3
R12278 vss.n6575 vss.n6574 9.3
R12279 vss.n6648 vss.n6647 9.3
R12280 vss.n6649 vss.n6648 9.3
R12281 vss.n6650 vss.n6649 9.3
R12282 vss.n6666 vss.n5834 9.3
R12283 vss.n6666 vss.n6665 9.3
R12284 vss.n6665 vss.n6664 9.3
R12285 vss.n6679 vss.n6678 9.3
R12286 vss.n6678 vss.n5820 9.3
R12287 vss.n5820 vss.n5819 9.3
R12288 vss.n6693 vss.n5808 9.3
R12289 vss.n5808 vss.n5807 9.3
R12290 vss.n5807 vss.n5806 9.3
R12291 vss.n6777 vss.n5746 9.3
R12292 vss.n6777 vss.n6776 9.3
R12293 vss.n6776 vss.n6775 9.3
R12294 vss.n6790 vss.n6789 9.3
R12295 vss.n6789 vss.n5732 9.3
R12296 vss.n5732 vss.n5731 9.3
R12297 vss.n6805 vss.n6804 9.3
R12298 vss.n6806 vss.n6805 9.3
R12299 vss.n6807 vss.n6806 9.3
R12300 vss.n6823 vss.n5708 9.3
R12301 vss.n6823 vss.n6822 9.3
R12302 vss.n6822 vss.n6821 9.3
R12303 vss.n6898 vss.n6897 9.3
R12304 vss.n6897 vss.n4230 9.3
R12305 vss.n4230 vss.n4229 9.3
R12306 vss.n4 vss.n4228 9.3
R12307 vss.n5654 vss.n5648 9.3
R12308 vss.n5649 vss.n5648 9.3
R12309 vss.n6885 vss.n5649 9.3
R12310 vss.n6880 vss.n5658 9.3
R12311 vss.n6880 vss.n6879 9.3
R12312 vss.n6879 vss.n6878 9.3
R12313 vss.n6873 vss.n6872 9.3
R12314 vss.n6873 vss.n5661 9.3
R12315 vss.n5661 vss.n5660 9.3
R12316 vss.n6862 vss.n5667 9.3
R12317 vss.n6863 vss.n6862 9.3
R12318 vss.n6864 vss.n6863 9.3
R12319 vss.n6858 vss.n6857 9.3
R12320 vss.n6857 vss.n6856 9.3
R12321 vss.n6856 vss.n6855 9.3
R12322 vss.n6850 vss.n6849 9.3
R12323 vss.n6850 vss.n5681 9.3
R12324 vss.n5681 vss.n5680 9.3
R12325 vss.n6839 vss.n5686 9.3
R12326 vss.n6840 vss.n6839 9.3
R12327 vss.n6841 vss.n6840 9.3
R12328 vss.n6835 vss.n6834 9.3
R12329 vss.n6834 vss.n6833 9.3
R12330 vss.n6833 vss.n6832 9.3
R12331 vss.n6828 vss.n6827 9.3
R12332 vss.n6829 vss.n6828 9.3
R12333 vss.n6830 vss.n6829 9.3
R12334 vss.n6813 vss.n6812 9.3
R12335 vss.n6812 vss.n5713 9.3
R12336 vss.n5713 vss.n5712 9.3
R12337 vss.n6800 vss.n5727 9.3
R12338 vss.n6800 vss.n6799 9.3
R12339 vss.n6799 vss.n6798 9.3
R12340 vss.n6782 vss.n6781 9.3
R12341 vss.n6783 vss.n6782 9.3
R12342 vss.n6784 vss.n6783 9.3
R12343 vss.n6763 vss.n6762 9.3
R12344 vss.n6764 vss.n6763 9.3
R12345 vss.n6765 vss.n6764 9.3
R12346 vss.n5759 vss.n5758 9.3
R12347 vss.n5760 vss.n5759 9.3
R12348 vss.n6754 vss.n5760 9.3
R12349 vss.n6749 vss.n5768 9.3
R12350 vss.n6749 vss.n6748 9.3
R12351 vss.n6748 vss.n6747 9.3
R12352 vss.n6742 vss.n6741 9.3
R12353 vss.n6742 vss.n5771 9.3
R12354 vss.n5771 vss.n5770 9.3
R12355 vss.n6731 vss.n5777 9.3
R12356 vss.n6732 vss.n6731 9.3
R12357 vss.n6733 vss.n6732 9.3
R12358 vss.n6727 vss.n6726 9.3
R12359 vss.n6726 vss.n6725 9.3
R12360 vss.n6725 vss.n6724 9.3
R12361 vss.n6719 vss.n6718 9.3
R12362 vss.n6719 vss.n5791 9.3
R12363 vss.n5791 vss.n5790 9.3
R12364 vss.n6708 vss.n5796 9.3
R12365 vss.n6709 vss.n6708 9.3
R12366 vss.n6710 vss.n6709 9.3
R12367 vss.n6704 vss.n6703 9.3
R12368 vss.n6703 vss.n6702 9.3
R12369 vss.n6702 vss.n6701 9.3
R12370 vss.n6689 vss.n5812 9.3
R12371 vss.n6689 vss.n6688 9.3
R12372 vss.n6688 vss.n6687 9.3
R12373 vss.n6671 vss.n6670 9.3
R12374 vss.n6672 vss.n6671 9.3
R12375 vss.n6673 vss.n6672 9.3
R12376 vss.n6656 vss.n6655 9.3
R12377 vss.n6655 vss.n5839 9.3
R12378 vss.n5839 vss.n5838 9.3
R12379 vss.n6638 vss.n5850 9.3
R12380 vss.n6638 vss.n5857 9.3
R12381 vss.n5857 vss.n5856 9.3
R12382 vss.n6634 vss.n6633 9.3
R12383 vss.n6633 vss.n6632 9.3
R12384 vss.n6632 vss.n6631 9.3
R12385 vss.n6626 vss.n6625 9.3
R12386 vss.n6626 vss.n5869 9.3
R12387 vss.n5869 vss.n5868 9.3
R12388 vss.n6615 vss.n5874 9.3
R12389 vss.n6616 vss.n6615 9.3
R12390 vss.n6617 vss.n6616 9.3
R12391 vss.n6611 vss.n6610 9.3
R12392 vss.n6610 vss.n6609 9.3
R12393 vss.n6609 vss.n6608 9.3
R12394 vss.n6603 vss.n6602 9.3
R12395 vss.n6603 vss.n5888 9.3
R12396 vss.n5888 vss.n5887 9.3
R12397 vss.n6592 vss.n5893 9.3
R12398 vss.n6593 vss.n6592 9.3
R12399 vss.n6594 vss.n6593 9.3
R12400 vss.n6588 vss.n6587 9.3
R12401 vss.n6587 vss.n6586 9.3
R12402 vss.n6586 vss.n6585 9.3
R12403 vss.n6581 vss.n6580 9.3
R12404 vss.n6582 vss.n6581 9.3
R12405 vss.n6583 vss.n6582 9.3
R12406 vss.n6566 vss.n6565 9.3
R12407 vss.n6565 vss.n5920 9.3
R12408 vss.n5920 vss.n5919 9.3
R12409 vss.n6553 vss.n5934 9.3
R12410 vss.n6553 vss.n6552 9.3
R12411 vss.n6552 vss.n6551 9.3
R12412 vss.n6535 vss.n6534 9.3
R12413 vss.n6536 vss.n6535 9.3
R12414 vss.n6537 vss.n6536 9.3
R12415 vss.n6516 vss.n6515 9.3
R12416 vss.n6517 vss.n6516 9.3
R12417 vss.n6518 vss.n6517 9.3
R12418 vss.n5966 vss.n5965 9.3
R12419 vss.n5967 vss.n5966 9.3
R12420 vss.n6507 vss.n5967 9.3
R12421 vss.n6502 vss.n5975 9.3
R12422 vss.n6502 vss.n6501 9.3
R12423 vss.n6501 vss.n6500 9.3
R12424 vss.n6495 vss.n6494 9.3
R12425 vss.n6495 vss.n5978 9.3
R12426 vss.n5978 vss.n5977 9.3
R12427 vss.n6484 vss.n5984 9.3
R12428 vss.n6485 vss.n6484 9.3
R12429 vss.n6486 vss.n6485 9.3
R12430 vss.n6480 vss.n6479 9.3
R12431 vss.n6479 vss.n6478 9.3
R12432 vss.n6478 vss.n6477 9.3
R12433 vss.n6472 vss.n6471 9.3
R12434 vss.n6472 vss.n5998 9.3
R12435 vss.n5998 vss.n5997 9.3
R12436 vss.n6461 vss.n6003 9.3
R12437 vss.n6462 vss.n6461 9.3
R12438 vss.n6463 vss.n6462 9.3
R12439 vss.n6457 vss.n6456 9.3
R12440 vss.n6456 vss.n6455 9.3
R12441 vss.n6455 vss.n6454 9.3
R12442 vss.n6442 vss.n6019 9.3
R12443 vss.n6442 vss.n6441 9.3
R12444 vss.n6441 vss.n6440 9.3
R12445 vss.n6424 vss.n6423 9.3
R12446 vss.n6425 vss.n6424 9.3
R12447 vss.n6426 vss.n6425 9.3
R12448 vss.n6409 vss.n6408 9.3
R12449 vss.n6408 vss.n6046 9.3
R12450 vss.n6046 vss.n6045 9.3
R12451 vss.n6391 vss.n6057 9.3
R12452 vss.n6391 vss.n6064 9.3
R12453 vss.n6064 vss.n6063 9.3
R12454 vss.n6387 vss.n6386 9.3
R12455 vss.n6386 vss.n6385 9.3
R12456 vss.n6385 vss.n6384 9.3
R12457 vss.n6379 vss.n6378 9.3
R12458 vss.n6379 vss.n6076 9.3
R12459 vss.n6076 vss.n6075 9.3
R12460 vss.n6368 vss.n6081 9.3
R12461 vss.n6369 vss.n6368 9.3
R12462 vss.n6370 vss.n6369 9.3
R12463 vss.n6364 vss.n6363 9.3
R12464 vss.n6363 vss.n6362 9.3
R12465 vss.n6362 vss.n6361 9.3
R12466 vss.n6356 vss.n6355 9.3
R12467 vss.n6356 vss.n6095 9.3
R12468 vss.n6095 vss.n6094 9.3
R12469 vss.n6345 vss.n6100 9.3
R12470 vss.n6346 vss.n6345 9.3
R12471 vss.n6347 vss.n6346 9.3
R12472 vss.n6341 vss.n6340 9.3
R12473 vss.n6340 vss.n6339 9.3
R12474 vss.n6339 vss.n6338 9.3
R12475 vss.n6334 vss.n6333 9.3
R12476 vss.n6335 vss.n6334 9.3
R12477 vss.n6336 vss.n6335 9.3
R12478 vss.n6319 vss.n6318 9.3
R12479 vss.n6318 vss.n6127 9.3
R12480 vss.n6127 vss.n6126 9.3
R12481 vss.n6306 vss.n6141 9.3
R12482 vss.n6306 vss.n6305 9.3
R12483 vss.n6305 vss.n6304 9.3
R12484 vss.n6288 vss.n6287 9.3
R12485 vss.n6289 vss.n6288 9.3
R12486 vss.n6290 vss.n6289 9.3
R12487 vss.n6269 vss.n6268 9.3
R12488 vss.n6270 vss.n6269 9.3
R12489 vss.n6271 vss.n6270 9.3
R12490 vss.n6173 vss.n6172 9.3
R12491 vss.n6174 vss.n6173 9.3
R12492 vss.n6260 vss.n6174 9.3
R12493 vss.n6255 vss.n6182 9.3
R12494 vss.n6255 vss.n6254 9.3
R12495 vss.n6254 vss.n6253 9.3
R12496 vss.n6248 vss.n6247 9.3
R12497 vss.n6248 vss.n6185 9.3
R12498 vss.n6185 vss.n6184 9.3
R12499 vss.n6237 vss.n6191 9.3
R12500 vss.n6238 vss.n6237 9.3
R12501 vss.n6239 vss.n6238 9.3
R12502 vss.n6200 vss.n6197 9.3
R12503 vss.n6212 vss.n6200 9.3
R12504 vss.n6212 vss.n6211 9.3
R12505 vss.n6218 vss.n6205 9.3
R12506 vss.n6914 vss.n4168 9.3
R12507 vss.n6905 vss.n4166 9.3
R12508 vss.n4145 vss.n4144 9.3
R12509 vss.n4147 vss.n4146 9.3
R12510 vss.n4143 vss.n4142 9.3
R12511 vss.n4150 vss.n4149 9.3
R12512 vss.n4155 vss.n4154 9.3
R12513 vss.n4152 vss.n4151 9.3
R12514 vss.n7066 vss.n7065 9.3
R12515 vss.n7082 vss.n7081 9.3
R12516 vss.n7097 vss.n7096 9.3
R12517 vss.n7112 vss.n7111 9.3
R12518 vss.n7128 vss.n7127 9.3
R12519 vss.n7146 vss.n7145 9.3
R12520 vss.n7156 vss.n7155 9.3
R12521 vss.n7175 vss.n7174 9.3
R12522 vss.n7190 vss.n7189 9.3
R12523 vss.n7186 vss.n7185 9.3
R12524 vss.n7185 vss.n7184 9.3
R12525 vss.n7184 vss.n7183 9.3
R12526 vss.n7173 vss.n7172 9.3
R12527 vss.n7130 vss.n7129 9.3
R12528 vss.n7099 vss.n7098 9.3
R12529 vss.n7069 vss.n7068 9.3
R12530 vss.n7064 vss.n7063 9.3
R12531 vss.n7063 vss.n7062 9.3
R12532 vss.n7062 vss.n7061 9.3
R12533 vss.n7080 vss.n7079 9.3
R12534 vss.n7079 vss.n7078 9.3
R12535 vss.n7078 vss.n7077 9.3
R12536 vss.n7084 vss.n7083 9.3
R12537 vss.n7095 vss.n7094 9.3
R12538 vss.n7094 vss.n7093 9.3
R12539 vss.n7093 vss.n7092 9.3
R12540 vss.n7110 vss.n7109 9.3
R12541 vss.n7109 vss.n7108 9.3
R12542 vss.n7108 vss.n7107 9.3
R12543 vss.n7114 vss.n7113 9.3
R12544 vss.n7126 vss.n7125 9.3
R12545 vss.n7125 vss.n7124 9.3
R12546 vss.n7124 vss.n7123 9.3
R12547 vss.n7144 vss.n7143 9.3
R12548 vss.n7143 vss.n7142 9.3
R12549 vss.n7142 vss.n7141 9.3
R12550 vss.n7148 vss.n7147 9.3
R12551 vss.n7154 vss.n7153 9.3
R12552 vss.n7171 vss.n7170 9.3
R12553 vss.n7170 vss.n7169 9.3
R12554 vss.n7169 vss.n7168 9.3
R12555 vss.n7188 vss.n7187 9.3
R12556 vss.n4100 vss.n4099 9.3
R12557 vss.n4102 vss.n4101 9.3
R12558 vss.n4098 vss.n4097 9.3
R12559 vss.n4105 vss.n4104 9.3
R12560 vss.n4110 vss.n4109 9.3
R12561 vss.n4107 vss.n4106 9.3
R12562 vss.n7205 vss.n7204 9.3
R12563 vss.n7220 vss.n7219 9.3
R12564 vss.n7235 vss.n7234 9.3
R12565 vss.n7250 vss.n7249 9.3
R12566 vss.n7281 vss.n7280 9.3
R12567 vss.n7296 vss.n7295 9.3
R12568 vss.n7311 vss.n7310 9.3
R12569 vss.n7326 vss.n7325 9.3
R12570 vss.n7341 vss.n7340 9.3
R12571 vss.n7356 vss.n7355 9.3
R12572 vss.n7397 vss.n7396 9.3
R12573 vss.n7413 vss.n7412 9.3
R12574 vss.n7428 vss.n7427 9.3
R12575 vss.n7443 vss.n7442 9.3
R12576 vss.n7459 vss.n7458 9.3
R12577 vss.n7470 vss.n7469 9.3
R12578 vss.n7469 vss.n7468 9.3
R12579 vss.n7468 vss.n7467 9.3
R12580 vss.n7457 vss.n7456 9.3
R12581 vss.n7439 vss.n7438 9.3
R12582 vss.n7438 vss.n7437 9.3
R12583 vss.n7437 vss.n7436 9.3
R12584 vss.n7426 vss.n7425 9.3
R12585 vss.n7408 vss.n7407 9.3
R12586 vss.n7407 vss.n7406 9.3
R12587 vss.n7406 vss.n7405 9.3
R12588 vss.n7395 vss.n7394 9.3
R12589 vss.n7358 vss.n7357 9.3
R12590 vss.n7328 vss.n7327 9.3
R12591 vss.n7298 vss.n7297 9.3
R12592 vss.n7268 vss.n7267 9.3
R12593 vss.n4137 vss.n4136 9.3
R12594 vss.n4136 vss.n4135 9.3
R12595 vss.n7263 vss.n7262 9.3
R12596 vss.n7246 vss.n7245 9.3
R12597 vss.n7245 vss.n7244 9.3
R12598 vss.n7244 vss.n7243 9.3
R12599 vss.n7233 vss.n7232 9.3
R12600 vss.n7216 vss.n7215 9.3
R12601 vss.n7215 vss.n7214 9.3
R12602 vss.n7214 vss.n7213 9.3
R12603 vss.n7203 vss.n7202 9.3
R12604 vss.n7201 vss.n7200 9.3
R12605 vss.n7200 vss.n7199 9.3
R12606 vss.n7199 vss.n7198 9.3
R12607 vss.n7218 vss.n7217 9.3
R12608 vss.n7231 vss.n7230 9.3
R12609 vss.n7230 vss.n7229 9.3
R12610 vss.n7229 vss.n7228 9.3
R12611 vss.n7248 vss.n7247 9.3
R12612 vss.n7261 vss.n7260 9.3
R12613 vss.n7260 vss.n7259 9.3
R12614 vss.n7259 vss.n7258 9.3
R12615 vss.n4124 vss.n4123 9.3
R12616 vss.n4123 vss.n4122 9.3
R12617 vss.n7279 vss.n7278 9.3
R12618 vss.n7278 vss.n7277 9.3
R12619 vss.n7277 vss.n7276 9.3
R12620 vss.n7283 vss.n7282 9.3
R12621 vss.n7294 vss.n7293 9.3
R12622 vss.n7293 vss.n7292 9.3
R12623 vss.n7292 vss.n7291 9.3
R12624 vss.n7309 vss.n7308 9.3
R12625 vss.n7308 vss.n7307 9.3
R12626 vss.n7307 vss.n7306 9.3
R12627 vss.n7313 vss.n7312 9.3
R12628 vss.n7324 vss.n7323 9.3
R12629 vss.n7323 vss.n7322 9.3
R12630 vss.n7322 vss.n7321 9.3
R12631 vss.n7339 vss.n7338 9.3
R12632 vss.n7338 vss.n7337 9.3
R12633 vss.n7337 vss.n7336 9.3
R12634 vss.n7343 vss.n7342 9.3
R12635 vss.n7354 vss.n7353 9.3
R12636 vss.n7353 vss.n7352 9.3
R12637 vss.n7352 vss.n7351 9.3
R12638 vss.n7373 vss.n7372 9.3
R12639 vss.n7372 vss.n7371 9.3
R12640 vss.n7371 vss.n7370 9.3
R12641 vss.n7393 vss.n7392 9.3
R12642 vss.n7392 vss.n7391 9.3
R12643 vss.n7391 vss.n7390 9.3
R12644 vss.n7411 vss.n7410 9.3
R12645 vss.n7424 vss.n7423 9.3
R12646 vss.n7423 vss.n7422 9.3
R12647 vss.n7422 vss.n7421 9.3
R12648 vss.n7441 vss.n7440 9.3
R12649 vss.n7454 vss.n7453 9.3
R12650 vss.n7453 vss.n7452 9.3
R12651 vss.n7452 vss.n7451 9.3
R12652 vss.n4014 vss.n4013 9.3
R12653 vss.n4007 vss.n4006 9.3
R12654 vss.n3588 vss.n3587 9.3
R12655 vss.n4005 vss.n4004 9.3
R12656 vss.n4009 vss.n4008 9.3
R12657 vss.n4012 vss.n4011 9.3
R12658 vss.n4016 vss.n4015 9.3
R12659 vss.n4093 vss.n4092 9.3
R12660 vss.n4092 vss.n4091 9.3
R12661 vss.n7516 vss.n7515 9.3
R12662 vss.n7515 vss.n7514 9.3
R12663 vss.n7530 vss.n7529 9.3
R12664 vss.n7529 vss.n7528 9.3
R12665 vss.n7544 vss.n7543 9.3
R12666 vss.n7543 vss.n7542 9.3
R12667 vss.n7558 vss.n7557 9.3
R12668 vss.n7557 vss.n7556 9.3
R12669 vss.n7572 vss.n7571 9.3
R12670 vss.n7571 vss.n7570 9.3
R12671 vss.n7586 vss.n7585 9.3
R12672 vss.n7585 vss.n7584 9.3
R12673 vss.n7602 vss.n7601 9.3
R12674 vss.n7601 vss.n7600 9.3
R12675 vss.n7621 vss.n7620 9.3
R12676 vss.n7620 vss.n7619 9.3
R12677 vss.n7635 vss.n7634 9.3
R12678 vss.n7634 vss.n7633 9.3
R12679 vss.n7649 vss.n7648 9.3
R12680 vss.n7648 vss.n7647 9.3
R12681 vss.n7663 vss.n7662 9.3
R12682 vss.n7662 vss.n7661 9.3
R12683 vss.n7677 vss.n7676 9.3
R12684 vss.n7676 vss.n7675 9.3
R12685 vss.n7691 vss.n7690 9.3
R12686 vss.n7690 vss.n7689 9.3
R12687 vss.n7705 vss.n7704 9.3
R12688 vss.n7704 vss.n7703 9.3
R12689 vss.n4082 vss.n4081 9.3
R12690 vss.n4081 vss.n4080 9.3
R12691 vss.n4071 vss.n4070 9.3
R12692 vss.n4070 vss.n4069 9.3
R12693 vss.n7724 vss.n7723 9.3
R12694 vss.n7723 vss.n7722 9.3
R12695 vss.n7738 vss.n7737 9.3
R12696 vss.n7737 vss.n7736 9.3
R12697 vss.n7752 vss.n7751 9.3
R12698 vss.n7751 vss.n7750 9.3
R12699 vss.n7766 vss.n7765 9.3
R12700 vss.n7765 vss.n7764 9.3
R12701 vss.n7780 vss.n7779 9.3
R12702 vss.n7779 vss.n7778 9.3
R12703 vss.n7794 vss.n7793 9.3
R12704 vss.n7793 vss.n7792 9.3
R12705 vss.n7810 vss.n7809 9.3
R12706 vss.n7809 vss.n7808 9.3
R12707 vss.n7829 vss.n7828 9.3
R12708 vss.n7828 vss.n7827 9.3
R12709 vss.n7843 vss.n7842 9.3
R12710 vss.n7842 vss.n7841 9.3
R12711 vss.n7858 vss.n7857 9.3
R12712 vss.n7857 vss.n7856 9.3
R12713 vss.n7872 vss.n7871 9.3
R12714 vss.n7871 vss.n7870 9.3
R12715 vss.n7886 vss.n7885 9.3
R12716 vss.n7885 vss.n7884 9.3
R12717 vss.n7900 vss.n7899 9.3
R12718 vss.n7899 vss.n7898 9.3
R12719 vss.n7914 vss.n7913 9.3
R12720 vss.n7913 vss.n7912 9.3
R12721 vss.n4060 vss.n4059 9.3
R12722 vss.n4059 vss.n4058 9.3
R12723 vss.n4049 vss.n4048 9.3
R12724 vss.n4048 vss.n4047 9.3
R12725 vss.n7933 vss.n7932 9.3
R12726 vss.n7932 vss.n7931 9.3
R12727 vss.n7947 vss.n7946 9.3
R12728 vss.n7946 vss.n7945 9.3
R12729 vss.n7961 vss.n7960 9.3
R12730 vss.n7960 vss.n7959 9.3
R12731 vss.n7975 vss.n7974 9.3
R12732 vss.n7974 vss.n7973 9.3
R12733 vss.n7989 vss.n7988 9.3
R12734 vss.n7988 vss.n7987 9.3
R12735 vss.n8003 vss.n8002 9.3
R12736 vss.n8002 vss.n8001 9.3
R12737 vss.n8019 vss.n8018 9.3
R12738 vss.n8018 vss.n8017 9.3
R12739 vss.n8038 vss.n8037 9.3
R12740 vss.n8037 vss.n8036 9.3
R12741 vss.n8052 vss.n8051 9.3
R12742 vss.n8051 vss.n8050 9.3
R12743 vss.n8066 vss.n8065 9.3
R12744 vss.n8065 vss.n8064 9.3
R12745 vss.n8080 vss.n8079 9.3
R12746 vss.n8079 vss.n8078 9.3
R12747 vss.n8094 vss.n8093 9.3
R12748 vss.n8093 vss.n8092 9.3
R12749 vss.n8108 vss.n8107 9.3
R12750 vss.n8107 vss.n8106 9.3
R12751 vss.n8122 vss.n8121 9.3
R12752 vss.n8121 vss.n8120 9.3
R12753 vss.n4038 vss.n4037 9.3
R12754 vss.n4037 vss.n4036 9.3
R12755 vss.n4027 vss.n4026 9.3
R12756 vss.n4026 vss.n4025 9.3
R12757 vss.n8141 vss.n8140 9.3
R12758 vss.n8140 vss.n8139 9.3
R12759 vss.n8155 vss.n8154 9.3
R12760 vss.n8154 vss.n8153 9.3
R12761 vss.n8169 vss.n8168 9.3
R12762 vss.n8168 vss.n8167 9.3
R12763 vss.n8183 vss.n8182 9.3
R12764 vss.n8182 vss.n8181 9.3
R12765 vss.n8197 vss.n8196 9.3
R12766 vss.n8196 vss.n8195 9.3
R12767 vss.n8211 vss.n8210 9.3
R12768 vss.n8210 vss.n8209 9.3
R12769 vss.n8228 vss.n8227 9.3
R12770 vss.n8227 vss.n8226 9.3
R12771 vss.n8241 vss.n8240 9.3
R12772 vss.n8240 vss.n8239 9.3
R12773 vss.n8260 vss.n8259 9.3
R12774 vss.n8259 vss.n8258 9.3
R12775 vss.n8274 vss.n8273 9.3
R12776 vss.n8273 vss.n8272 9.3
R12777 vss.n8288 vss.n8287 9.3
R12778 vss.n8287 vss.n8286 9.3
R12779 vss.n8302 vss.n8301 9.3
R12780 vss.n8301 vss.n8300 9.3
R12781 vss.n8316 vss.n8315 9.3
R12782 vss.n8315 vss.n8314 9.3
R12783 vss.n8330 vss.n8329 9.3
R12784 vss.n8329 vss.n8328 9.3
R12785 vss.n3553 vss.n3552 9.3
R12786 vss.n3552 vss.n3551 9.3
R12787 vss.n3542 vss.n3541 9.3
R12788 vss.n3541 vss.n3540 9.3
R12789 vss.n8349 vss.n8348 9.3
R12790 vss.n8348 vss.n8347 9.3
R12791 vss.n8363 vss.n8362 9.3
R12792 vss.n8362 vss.n8361 9.3
R12793 vss.n8377 vss.n8376 9.3
R12794 vss.n8376 vss.n8375 9.3
R12795 vss.n8391 vss.n8390 9.3
R12796 vss.n8390 vss.n8389 9.3
R12797 vss.n8405 vss.n8404 9.3
R12798 vss.n8404 vss.n8403 9.3
R12799 vss.n8419 vss.n8418 9.3
R12800 vss.n8418 vss.n8417 9.3
R12801 vss.n8435 vss.n8434 9.3
R12802 vss.n8434 vss.n8433 9.3
R12803 vss.n8454 vss.n8453 9.3
R12804 vss.n8453 vss.n8452 9.3
R12805 vss.n8468 vss.n8467 9.3
R12806 vss.n8467 vss.n8466 9.3
R12807 vss.n8482 vss.n8481 9.3
R12808 vss.n8481 vss.n8480 9.3
R12809 vss.n8496 vss.n8495 9.3
R12810 vss.n8495 vss.n8494 9.3
R12811 vss.n8510 vss.n8509 9.3
R12812 vss.n8509 vss.n8508 9.3
R12813 vss.n8524 vss.n8523 9.3
R12814 vss.n8523 vss.n8522 9.3
R12815 vss.n8538 vss.n8537 9.3
R12816 vss.n8537 vss.n8536 9.3
R12817 vss.n3531 vss.n3530 9.3
R12818 vss.n3530 vss.n3529 9.3
R12819 vss.n3520 vss.n3519 9.3
R12820 vss.n3519 vss.n3518 9.3
R12821 vss.n8557 vss.n8556 9.3
R12822 vss.n8556 vss.n8555 9.3
R12823 vss.n8571 vss.n8570 9.3
R12824 vss.n8570 vss.n8569 9.3
R12825 vss.n8585 vss.n8584 9.3
R12826 vss.n8584 vss.n8583 9.3
R12827 vss.n8599 vss.n8598 9.3
R12828 vss.n8598 vss.n8597 9.3
R12829 vss.n8613 vss.n8612 9.3
R12830 vss.n8612 vss.n8611 9.3
R12831 vss.n8627 vss.n8626 9.3
R12832 vss.n8626 vss.n8625 9.3
R12833 vss.n8643 vss.n8642 9.3
R12834 vss.n8642 vss.n8641 9.3
R12835 vss.n8662 vss.n8661 9.3
R12836 vss.n8661 vss.n8660 9.3
R12837 vss.n8676 vss.n8675 9.3
R12838 vss.n8675 vss.n8674 9.3
R12839 vss.n8690 vss.n8689 9.3
R12840 vss.n8689 vss.n8688 9.3
R12841 vss.n8704 vss.n8703 9.3
R12842 vss.n8703 vss.n8702 9.3
R12843 vss.n8718 vss.n8717 9.3
R12844 vss.n8717 vss.n8716 9.3
R12845 vss.n8732 vss.n8731 9.3
R12846 vss.n8731 vss.n8730 9.3
R12847 vss.n8746 vss.n8745 9.3
R12848 vss.n8745 vss.n8744 9.3
R12849 vss.n3509 vss.n3508 9.3
R12850 vss.n3508 vss.n3507 9.3
R12851 vss.n3498 vss.n3497 9.3
R12852 vss.n3497 vss.n3496 9.3
R12853 vss.n8765 vss.n8764 9.3
R12854 vss.n8764 vss.n8763 9.3
R12855 vss.n8779 vss.n8778 9.3
R12856 vss.n8778 vss.n8777 9.3
R12857 vss.n8793 vss.n8792 9.3
R12858 vss.n8792 vss.n8791 9.3
R12859 vss.n8807 vss.n8806 9.3
R12860 vss.n8806 vss.n8805 9.3
R12861 vss.n8821 vss.n8820 9.3
R12862 vss.n8820 vss.n8819 9.3
R12863 vss.n8835 vss.n8834 9.3
R12864 vss.n8834 vss.n8833 9.3
R12865 vss.n8851 vss.n8850 9.3
R12866 vss.n8850 vss.n8849 9.3
R12867 vss.n8870 vss.n8869 9.3
R12868 vss.n8869 vss.n8868 9.3
R12869 vss.n8884 vss.n8883 9.3
R12870 vss.n8883 vss.n8882 9.3
R12871 vss.n8898 vss.n8897 9.3
R12872 vss.n8897 vss.n8896 9.3
R12873 vss.n8912 vss.n8911 9.3
R12874 vss.n8911 vss.n8910 9.3
R12875 vss.n1782 vss.n1781 9.3
R12876 vss.n1727 vss.n1726 9.3
R12877 vss.n1697 vss.n1696 9.3
R12878 vss.n1695 vss.n1694 9.3
R12879 vss.n1693 vss.n1692 9.3
R12880 vss.n1692 vss.n1691 9.3
R12881 vss.n1691 vss.n1690 9.3
R12882 vss.n1708 vss.n1707 9.3
R12883 vss.n1707 vss.n1706 9.3
R12884 vss.n1706 vss.n1705 9.3
R12885 vss.n1712 vss.n1711 9.3
R12886 vss.n1710 vss.n1709 9.3
R12887 vss.n1725 vss.n1724 9.3
R12888 vss.n1723 vss.n1722 9.3
R12889 vss.n1722 vss.n1721 9.3
R12890 vss.n1721 vss.n1720 9.3
R12891 vss.n1738 vss.n1737 9.3
R12892 vss.n1737 vss.n1736 9.3
R12893 vss.n1736 vss.n1735 9.3
R12894 vss.n1742 vss.n1741 9.3
R12895 vss.n1740 vss.n1739 9.3
R12896 vss.n1760 vss.n1759 9.3
R12897 vss.n1759 vss.n1758 9.3
R12898 vss.n1758 vss.n1757 9.3
R12899 vss.n1780 vss.n1779 9.3
R12900 vss.n1779 vss.n1778 9.3
R12901 vss.n1778 vss.n1777 9.3
R12902 vss.n1797 vss.n1796 9.3
R12903 vss.n1796 vss.n1795 9.3
R12904 vss.n1795 vss.n1794 9.3
R12905 vss.n1784 vss.n1783 9.3
R12906 vss.n3399 vss.n3398 9.3
R12907 vss.n3369 vss.n3368 9.3
R12908 vss.n3339 vss.n3338 9.3
R12909 vss.n3335 vss.n3334 9.3
R12910 vss.n3318 vss.n3317 9.3
R12911 vss.n3302 vss.n3301 9.3
R12912 vss.n3286 vss.n3285 9.3
R12913 vss.n3270 vss.n3269 9.3
R12914 vss.n3254 vss.n3253 9.3
R12915 vss.n3238 vss.n3237 9.3
R12916 vss.n3218 vss.n3217 9.3
R12917 vss.n3211 vss.n3210 9.3
R12918 vss.n3175 vss.n3174 9.3
R12919 vss.n3143 vss.n3142 9.3
R12920 vss.n3110 vss.n3109 9.3
R12921 vss.n3090 vss.n3089 9.3
R12922 vss.n3074 vss.n3073 9.3
R12923 vss.n3058 vss.n3057 9.3
R12924 vss.n3042 vss.n3041 9.3
R12925 vss.n3026 vss.n3025 9.3
R12926 vss.n3009 vss.n3008 9.3
R12927 vss.n2993 vss.n2992 9.3
R12928 vss.n2973 vss.n2972 9.3
R12929 vss.n2947 vss.n2946 9.3
R12930 vss.n2915 vss.n2914 9.3
R12931 vss.n2882 vss.n2881 9.3
R12932 vss.n2850 vss.n2849 9.3
R12933 vss.n2846 vss.n2845 9.3
R12934 vss.n2818 vss.n2817 9.3
R12935 vss.n2803 vss.n2802 9.3
R12936 vss.n2787 vss.n2786 9.3
R12937 vss.n2771 vss.n2770 9.3
R12938 vss.n2755 vss.n2754 9.3
R12939 vss.n2735 vss.n2734 9.3
R12940 vss.n2729 vss.n2728 9.3
R12941 vss.n2692 vss.n2691 9.3
R12942 vss.n2660 vss.n2659 9.3
R12943 vss.n2628 vss.n2627 9.3
R12944 vss.n2607 vss.n2606 9.3
R12945 vss.n2591 vss.n2590 9.3
R12946 vss.n2575 vss.n2574 9.3
R12947 vss.n2559 vss.n2558 9.3
R12948 vss.n2543 vss.n2542 9.3
R12949 vss.n2527 vss.n2526 9.3
R12950 vss.n2511 vss.n2510 9.3
R12951 vss.n2490 vss.n2489 9.3
R12952 vss.n2464 vss.n2463 9.3
R12953 vss.n2432 vss.n2431 9.3
R12954 vss.n2400 vss.n2399 9.3
R12955 vss.n2367 vss.n2366 9.3
R12956 vss.n2363 vss.n2362 9.3
R12957 vss.n2347 vss.n2346 9.3
R12958 vss.n2331 vss.n2330 9.3
R12959 vss.n2315 vss.n2314 9.3
R12960 vss.n2299 vss.n2298 9.3
R12961 vss.n2282 vss.n2281 9.3
R12962 vss.n2266 vss.n2265 9.3
R12963 vss.n2246 vss.n2245 9.3
R12964 vss.n2240 vss.n2239 9.3
R12965 vss.n2204 vss.n2203 9.3
R12966 vss.n2171 vss.n2170 9.3
R12967 vss.n2139 vss.n2138 9.3
R12968 vss.n2119 vss.n2118 9.3
R12969 vss.n2103 vss.n2102 9.3
R12970 vss.n2086 vss.n2085 9.3
R12971 vss.n2070 vss.n2069 9.3
R12972 vss.n2054 vss.n2053 9.3
R12973 vss.n2038 vss.n2037 9.3
R12974 vss.n2022 vss.n2021 9.3
R12975 vss.n2002 vss.n2001 9.3
R12976 vss.n1975 vss.n1974 9.3
R12977 vss.n1943 vss.n1942 9.3
R12978 vss.n1911 vss.n1910 9.3
R12979 vss.n1878 vss.n1877 9.3
R12980 vss.n1874 vss.n1873 9.3
R12981 vss.n1859 vss.n1858 9.3
R12982 vss.n1844 vss.n1843 9.3
R12983 vss.n1829 vss.n1828 9.3
R12984 vss.n1814 vss.n1813 9.3
R12985 vss.n1799 vss.n1798 9.3
R12986 vss.n1801 vss.n1800 9.3
R12987 vss.n1812 vss.n1811 9.3
R12988 vss.n1811 vss.n1810 9.3
R12989 vss.n1810 vss.n1809 9.3
R12990 vss.n1827 vss.n1826 9.3
R12991 vss.n1826 vss.n1825 9.3
R12992 vss.n1825 vss.n1824 9.3
R12993 vss.n1816 vss.n1815 9.3
R12994 vss.n1831 vss.n1830 9.3
R12995 vss.n1842 vss.n1841 9.3
R12996 vss.n1841 vss.n1840 9.3
R12997 vss.n1840 vss.n1839 9.3
R12998 vss.n1857 vss.n1856 9.3
R12999 vss.n1856 vss.n1855 9.3
R13000 vss.n1855 vss.n1854 9.3
R13001 vss.n1846 vss.n1845 9.3
R13002 vss.n1861 vss.n1860 9.3
R13003 vss.n1872 vss.n1871 9.3
R13004 vss.n1871 vss.n1870 9.3
R13005 vss.n1870 vss.n1869 9.3
R13006 vss.n1649 vss.n1648 9.3
R13007 vss.n1648 vss.n1647 9.3
R13008 vss.n1637 vss.n1636 9.3
R13009 vss.n1636 vss.n1635 9.3
R13010 vss.n1891 vss.n1890 9.3
R13011 vss.n1890 vss.n1889 9.3
R13012 vss.n1889 vss.n1888 9.3
R13013 vss.n1895 vss.n1894 9.3
R13014 vss.n1893 vss.n1892 9.3
R13015 vss.n1909 vss.n1908 9.3
R13016 vss.n1907 vss.n1906 9.3
R13017 vss.n1906 vss.n1905 9.3
R13018 vss.n1905 vss.n1904 9.3
R13019 vss.n1923 vss.n1922 9.3
R13020 vss.n1922 vss.n1921 9.3
R13021 vss.n1921 vss.n1920 9.3
R13022 vss.n1927 vss.n1926 9.3
R13023 vss.n1925 vss.n1924 9.3
R13024 vss.n1941 vss.n1940 9.3
R13025 vss.n1939 vss.n1938 9.3
R13026 vss.n1938 vss.n1937 9.3
R13027 vss.n1937 vss.n1936 9.3
R13028 vss.n1955 vss.n1954 9.3
R13029 vss.n1954 vss.n1953 9.3
R13030 vss.n1953 vss.n1952 9.3
R13031 vss.n1959 vss.n1958 9.3
R13032 vss.n1957 vss.n1956 9.3
R13033 vss.n1973 vss.n1972 9.3
R13034 vss.n1971 vss.n1970 9.3
R13035 vss.n1970 vss.n1969 9.3
R13036 vss.n1969 vss.n1968 9.3
R13037 vss.n1991 vss.n1990 9.3
R13038 vss.n1990 vss.n1989 9.3
R13039 vss.n1989 vss.n1988 9.3
R13040 vss.n1995 vss.n1994 9.3
R13041 vss.n1993 vss.n1992 9.3
R13042 vss.n2020 vss.n2019 9.3
R13043 vss.n2019 vss.n2018 9.3
R13044 vss.n2018 vss.n2017 9.3
R13045 vss.n2004 vss.n2003 9.3
R13046 vss.n2024 vss.n2023 9.3
R13047 vss.n2036 vss.n2035 9.3
R13048 vss.n2035 vss.n2034 9.3
R13049 vss.n2034 vss.n2033 9.3
R13050 vss.n2052 vss.n2051 9.3
R13051 vss.n2051 vss.n2050 9.3
R13052 vss.n2050 vss.n2049 9.3
R13053 vss.n2040 vss.n2039 9.3
R13054 vss.n2056 vss.n2055 9.3
R13055 vss.n2068 vss.n2067 9.3
R13056 vss.n2067 vss.n2066 9.3
R13057 vss.n2066 vss.n2065 9.3
R13058 vss.n2084 vss.n2083 9.3
R13059 vss.n2083 vss.n2082 9.3
R13060 vss.n2082 vss.n2081 9.3
R13061 vss.n2072 vss.n2071 9.3
R13062 vss.n2088 vss.n2087 9.3
R13063 vss.n2100 vss.n2099 9.3
R13064 vss.n2099 vss.n2098 9.3
R13065 vss.n2098 vss.n2097 9.3
R13066 vss.n2117 vss.n2116 9.3
R13067 vss.n2116 vss.n2115 9.3
R13068 vss.n2115 vss.n2114 9.3
R13069 vss.n2105 vss.n2104 9.3
R13070 vss.n1622 vss.n1621 9.3
R13071 vss.n1621 vss.n1620 9.3
R13072 vss.n1610 vss.n1609 9.3
R13073 vss.n1609 vss.n1608 9.3
R13074 vss.n2123 vss.n2122 9.3
R13075 vss.n2137 vss.n2136 9.3
R13076 vss.n2135 vss.n2134 9.3
R13077 vss.n2134 vss.n2133 9.3
R13078 vss.n2133 vss.n2132 9.3
R13079 vss.n2151 vss.n2150 9.3
R13080 vss.n2150 vss.n2149 9.3
R13081 vss.n2149 vss.n2148 9.3
R13082 vss.n2155 vss.n2154 9.3
R13083 vss.n2153 vss.n2152 9.3
R13084 vss.n2169 vss.n2168 9.3
R13085 vss.n2167 vss.n2166 9.3
R13086 vss.n2166 vss.n2165 9.3
R13087 vss.n2165 vss.n2164 9.3
R13088 vss.n2183 vss.n2182 9.3
R13089 vss.n2182 vss.n2181 9.3
R13090 vss.n2181 vss.n2180 9.3
R13091 vss.n2187 vss.n2186 9.3
R13092 vss.n2185 vss.n2184 9.3
R13093 vss.n2202 vss.n2201 9.3
R13094 vss.n2200 vss.n2199 9.3
R13095 vss.n2199 vss.n2198 9.3
R13096 vss.n2198 vss.n2197 9.3
R13097 vss.n2216 vss.n2215 9.3
R13098 vss.n2215 vss.n2214 9.3
R13099 vss.n2214 vss.n2213 9.3
R13100 vss.n2220 vss.n2219 9.3
R13101 vss.n2218 vss.n2217 9.3
R13102 vss.n2238 vss.n2237 9.3
R13103 vss.n2236 vss.n2235 9.3
R13104 vss.n2235 vss.n2234 9.3
R13105 vss.n2234 vss.n2233 9.3
R13106 vss.n2248 vss.n2247 9.3
R13107 vss.n2264 vss.n2263 9.3
R13108 vss.n2263 vss.n2262 9.3
R13109 vss.n2262 vss.n2261 9.3
R13110 vss.n2280 vss.n2279 9.3
R13111 vss.n2279 vss.n2278 9.3
R13112 vss.n2278 vss.n2277 9.3
R13113 vss.n2268 vss.n2267 9.3
R13114 vss.n2284 vss.n2283 9.3
R13115 vss.n2296 vss.n2295 9.3
R13116 vss.n2295 vss.n2294 9.3
R13117 vss.n2294 vss.n2293 9.3
R13118 vss.n2313 vss.n2312 9.3
R13119 vss.n2312 vss.n2311 9.3
R13120 vss.n2311 vss.n2310 9.3
R13121 vss.n2301 vss.n2300 9.3
R13122 vss.n2317 vss.n2316 9.3
R13123 vss.n2329 vss.n2328 9.3
R13124 vss.n2328 vss.n2327 9.3
R13125 vss.n2327 vss.n2326 9.3
R13126 vss.n2345 vss.n2344 9.3
R13127 vss.n2344 vss.n2343 9.3
R13128 vss.n2343 vss.n2342 9.3
R13129 vss.n2333 vss.n2332 9.3
R13130 vss.n2349 vss.n2348 9.3
R13131 vss.n2361 vss.n2360 9.3
R13132 vss.n2360 vss.n2359 9.3
R13133 vss.n2359 vss.n2358 9.3
R13134 vss.n1597 vss.n1596 9.3
R13135 vss.n1596 vss.n1595 9.3
R13136 vss.n1585 vss.n1584 9.3
R13137 vss.n1584 vss.n1583 9.3
R13138 vss.n2379 vss.n2378 9.3
R13139 vss.n2378 vss.n2377 9.3
R13140 vss.n2377 vss.n2376 9.3
R13141 vss.n2383 vss.n2382 9.3
R13142 vss.n2381 vss.n2380 9.3
R13143 vss.n2397 vss.n2396 9.3
R13144 vss.n2395 vss.n2394 9.3
R13145 vss.n2394 vss.n2393 9.3
R13146 vss.n2393 vss.n2392 9.3
R13147 vss.n2412 vss.n2411 9.3
R13148 vss.n2411 vss.n2410 9.3
R13149 vss.n2410 vss.n2409 9.3
R13150 vss.n2416 vss.n2415 9.3
R13151 vss.n2414 vss.n2413 9.3
R13152 vss.n2430 vss.n2429 9.3
R13153 vss.n2428 vss.n2427 9.3
R13154 vss.n2427 vss.n2426 9.3
R13155 vss.n2426 vss.n2425 9.3
R13156 vss.n2444 vss.n2443 9.3
R13157 vss.n2443 vss.n2442 9.3
R13158 vss.n2442 vss.n2441 9.3
R13159 vss.n2448 vss.n2447 9.3
R13160 vss.n2446 vss.n2445 9.3
R13161 vss.n2462 vss.n2461 9.3
R13162 vss.n2460 vss.n2459 9.3
R13163 vss.n2459 vss.n2458 9.3
R13164 vss.n2458 vss.n2457 9.3
R13165 vss.n2480 vss.n2479 9.3
R13166 vss.n2479 vss.n2478 9.3
R13167 vss.n2478 vss.n2477 9.3
R13168 vss.n2484 vss.n2483 9.3
R13169 vss.n2482 vss.n2481 9.3
R13170 vss.n2508 vss.n2507 9.3
R13171 vss.n2507 vss.n2506 9.3
R13172 vss.n2506 vss.n2505 9.3
R13173 vss.n2492 vss.n2491 9.3
R13174 vss.n2513 vss.n2512 9.3
R13175 vss.n2525 vss.n2524 9.3
R13176 vss.n2524 vss.n2523 9.3
R13177 vss.n2523 vss.n2522 9.3
R13178 vss.n2541 vss.n2540 9.3
R13179 vss.n2540 vss.n2539 9.3
R13180 vss.n2539 vss.n2538 9.3
R13181 vss.n2529 vss.n2528 9.3
R13182 vss.n2545 vss.n2544 9.3
R13183 vss.n2557 vss.n2556 9.3
R13184 vss.n2556 vss.n2555 9.3
R13185 vss.n2555 vss.n2554 9.3
R13186 vss.n2573 vss.n2572 9.3
R13187 vss.n2572 vss.n2571 9.3
R13188 vss.n2571 vss.n2570 9.3
R13189 vss.n2561 vss.n2560 9.3
R13190 vss.n2577 vss.n2576 9.3
R13191 vss.n2589 vss.n2588 9.3
R13192 vss.n2588 vss.n2587 9.3
R13193 vss.n2587 vss.n2586 9.3
R13194 vss.n2605 vss.n2604 9.3
R13195 vss.n2604 vss.n2603 9.3
R13196 vss.n2603 vss.n2602 9.3
R13197 vss.n2593 vss.n2592 9.3
R13198 vss.n1572 vss.n1571 9.3
R13199 vss.n1571 vss.n1570 9.3
R13200 vss.n1559 vss.n1558 9.3
R13201 vss.n1558 vss.n1557 9.3
R13202 vss.n2612 vss.n2611 9.3
R13203 vss.n2626 vss.n2625 9.3
R13204 vss.n2624 vss.n2623 9.3
R13205 vss.n2623 vss.n2622 9.3
R13206 vss.n2622 vss.n2621 9.3
R13207 vss.n2640 vss.n2639 9.3
R13208 vss.n2639 vss.n2638 9.3
R13209 vss.n2638 vss.n2637 9.3
R13210 vss.n2644 vss.n2643 9.3
R13211 vss.n2642 vss.n2641 9.3
R13212 vss.n2658 vss.n2657 9.3
R13213 vss.n2656 vss.n2655 9.3
R13214 vss.n2655 vss.n2654 9.3
R13215 vss.n2654 vss.n2653 9.3
R13216 vss.n2672 vss.n2671 9.3
R13217 vss.n2671 vss.n2670 9.3
R13218 vss.n2670 vss.n2669 9.3
R13219 vss.n2676 vss.n2675 9.3
R13220 vss.n2674 vss.n2673 9.3
R13221 vss.n2690 vss.n2689 9.3
R13222 vss.n2688 vss.n2687 9.3
R13223 vss.n2687 vss.n2686 9.3
R13224 vss.n2686 vss.n2685 9.3
R13225 vss.n2704 vss.n2703 9.3
R13226 vss.n2703 vss.n2702 9.3
R13227 vss.n2702 vss.n2701 9.3
R13228 vss.n2708 vss.n2707 9.3
R13229 vss.n2706 vss.n2705 9.3
R13230 vss.n2727 vss.n2726 9.3
R13231 vss.n2725 vss.n2724 9.3
R13232 vss.n2724 vss.n2723 9.3
R13233 vss.n2723 vss.n2722 9.3
R13234 vss.n2737 vss.n2736 9.3
R13235 vss.n2753 vss.n2752 9.3
R13236 vss.n2752 vss.n2751 9.3
R13237 vss.n2751 vss.n2750 9.3
R13238 vss.n2769 vss.n2768 9.3
R13239 vss.n2768 vss.n2767 9.3
R13240 vss.n2767 vss.n2766 9.3
R13241 vss.n2757 vss.n2756 9.3
R13242 vss.n2773 vss.n2772 9.3
R13243 vss.n2785 vss.n2784 9.3
R13244 vss.n2784 vss.n2783 9.3
R13245 vss.n2783 vss.n2782 9.3
R13246 vss.n2801 vss.n2800 9.3
R13247 vss.n2800 vss.n2799 9.3
R13248 vss.n2799 vss.n2798 9.3
R13249 vss.n2789 vss.n2788 9.3
R13250 vss.n2805 vss.n2804 9.3
R13251 vss.n2816 vss.n2815 9.3
R13252 vss.n2815 vss.n2814 9.3
R13253 vss.n2814 vss.n2813 9.3
R13254 vss.n2831 vss.n2830 9.3
R13255 vss.n2830 vss.n2829 9.3
R13256 vss.n2829 vss.n2828 9.3
R13257 vss.n2821 vss.n2820 9.3
R13258 vss.n2842 vss.n2834 9.3
R13259 vss.n2842 vss.n2841 9.3
R13260 vss.n2841 vss.n2840 9.3
R13261 vss.n1542 vss.n1541 9.3
R13262 vss.n1541 vss.n1540 9.3
R13263 vss.n1527 vss.n1526 9.3
R13264 vss.n1526 vss.n1525 9.3
R13265 vss.n2862 vss.n2861 9.3
R13266 vss.n2861 vss.n2860 9.3
R13267 vss.n2860 vss.n2859 9.3
R13268 vss.n2866 vss.n2865 9.3
R13269 vss.n2864 vss.n2863 9.3
R13270 vss.n2880 vss.n2879 9.3
R13271 vss.n2878 vss.n2877 9.3
R13272 vss.n2877 vss.n2876 9.3
R13273 vss.n2876 vss.n2875 9.3
R13274 vss.n2894 vss.n2893 9.3
R13275 vss.n2893 vss.n2892 9.3
R13276 vss.n2892 vss.n2891 9.3
R13277 vss.n2898 vss.n2897 9.3
R13278 vss.n2896 vss.n2895 9.3
R13279 vss.n2912 vss.n2911 9.3
R13280 vss.n2910 vss.n2909 9.3
R13281 vss.n2909 vss.n2908 9.3
R13282 vss.n2908 vss.n2907 9.3
R13283 vss.n2927 vss.n2926 9.3
R13284 vss.n2926 vss.n2925 9.3
R13285 vss.n2925 vss.n2924 9.3
R13286 vss.n2931 vss.n2930 9.3
R13287 vss.n2929 vss.n2928 9.3
R13288 vss.n2945 vss.n2944 9.3
R13289 vss.n2943 vss.n2942 9.3
R13290 vss.n2942 vss.n2941 9.3
R13291 vss.n2941 vss.n2940 9.3
R13292 vss.n2963 vss.n2962 9.3
R13293 vss.n2962 vss.n2961 9.3
R13294 vss.n2961 vss.n2960 9.3
R13295 vss.n2967 vss.n2966 9.3
R13296 vss.n2965 vss.n2964 9.3
R13297 vss.n2991 vss.n2990 9.3
R13298 vss.n2990 vss.n2989 9.3
R13299 vss.n2989 vss.n2988 9.3
R13300 vss.n2975 vss.n2974 9.3
R13301 vss.n2995 vss.n2994 9.3
R13302 vss.n3007 vss.n3006 9.3
R13303 vss.n3006 vss.n3005 9.3
R13304 vss.n3005 vss.n3004 9.3
R13305 vss.n3024 vss.n3023 9.3
R13306 vss.n3023 vss.n3022 9.3
R13307 vss.n3022 vss.n3021 9.3
R13308 vss.n3011 vss.n3010 9.3
R13309 vss.n3028 vss.n3027 9.3
R13310 vss.n3040 vss.n3039 9.3
R13311 vss.n3039 vss.n3038 9.3
R13312 vss.n3038 vss.n3037 9.3
R13313 vss.n3056 vss.n3055 9.3
R13314 vss.n3055 vss.n3054 9.3
R13315 vss.n3054 vss.n3053 9.3
R13316 vss.n3044 vss.n3043 9.3
R13317 vss.n3060 vss.n3059 9.3
R13318 vss.n3072 vss.n3071 9.3
R13319 vss.n3071 vss.n3070 9.3
R13320 vss.n3070 vss.n3069 9.3
R13321 vss.n3088 vss.n3087 9.3
R13322 vss.n3087 vss.n3086 9.3
R13323 vss.n3086 vss.n3085 9.3
R13324 vss.n3076 vss.n3075 9.3
R13325 vss.n1514 vss.n1513 9.3
R13326 vss.n1513 vss.n1512 9.3
R13327 vss.n1502 vss.n1501 9.3
R13328 vss.n1501 vss.n1500 9.3
R13329 vss.n3094 vss.n3093 9.3
R13330 vss.n3108 vss.n3107 9.3
R13331 vss.n3106 vss.n3105 9.3
R13332 vss.n3105 vss.n3104 9.3
R13333 vss.n3104 vss.n3103 9.3
R13334 vss.n3123 vss.n3122 9.3
R13335 vss.n3122 vss.n3121 9.3
R13336 vss.n3121 vss.n3120 9.3
R13337 vss.n3127 vss.n3126 9.3
R13338 vss.n3125 vss.n3124 9.3
R13339 vss.n3141 vss.n3140 9.3
R13340 vss.n3139 vss.n3138 9.3
R13341 vss.n3138 vss.n3137 9.3
R13342 vss.n3137 vss.n3136 9.3
R13343 vss.n3155 vss.n3154 9.3
R13344 vss.n3154 vss.n3153 9.3
R13345 vss.n3153 vss.n3152 9.3
R13346 vss.n3159 vss.n3158 9.3
R13347 vss.n3157 vss.n3156 9.3
R13348 vss.n3173 vss.n3172 9.3
R13349 vss.n3171 vss.n3170 9.3
R13350 vss.n3170 vss.n3169 9.3
R13351 vss.n3169 vss.n3168 9.3
R13352 vss.n3187 vss.n3186 9.3
R13353 vss.n3186 vss.n3185 9.3
R13354 vss.n3185 vss.n3184 9.3
R13355 vss.n3191 vss.n3190 9.3
R13356 vss.n3189 vss.n3188 9.3
R13357 vss.n3209 vss.n3208 9.3
R13358 vss.n3207 vss.n3206 9.3
R13359 vss.n3206 vss.n3205 9.3
R13360 vss.n3205 vss.n3204 9.3
R13361 vss.n3220 vss.n3219 9.3
R13362 vss.n3236 vss.n3235 9.3
R13363 vss.n3235 vss.n3234 9.3
R13364 vss.n3234 vss.n3233 9.3
R13365 vss.n3252 vss.n3251 9.3
R13366 vss.n3251 vss.n3250 9.3
R13367 vss.n3250 vss.n3249 9.3
R13368 vss.n3240 vss.n3239 9.3
R13369 vss.n3256 vss.n3255 9.3
R13370 vss.n3268 vss.n3267 9.3
R13371 vss.n3267 vss.n3266 9.3
R13372 vss.n3266 vss.n3265 9.3
R13373 vss.n3284 vss.n3283 9.3
R13374 vss.n3283 vss.n3282 9.3
R13375 vss.n3282 vss.n3281 9.3
R13376 vss.n3272 vss.n3271 9.3
R13377 vss.n3288 vss.n3287 9.3
R13378 vss.n3300 vss.n3299 9.3
R13379 vss.n3299 vss.n3298 9.3
R13380 vss.n3298 vss.n3297 9.3
R13381 vss.n3316 vss.n3315 9.3
R13382 vss.n3315 vss.n3314 9.3
R13383 vss.n3314 vss.n3313 9.3
R13384 vss.n3304 vss.n3303 9.3
R13385 vss.n3320 vss.n3319 9.3
R13386 vss.n3332 vss.n3331 9.3
R13387 vss.n3331 vss.n3330 9.3
R13388 vss.n3330 vss.n3329 9.3
R13389 vss.n1487 vss.n1486 9.3
R13390 vss.n1486 vss.n1485 9.3
R13391 vss.n1475 vss.n1474 9.3
R13392 vss.n1474 vss.n1473 9.3
R13393 vss.n3350 vss.n3349 9.3
R13394 vss.n3349 vss.n3348 9.3
R13395 vss.n3348 vss.n3347 9.3
R13396 vss.n3354 vss.n3353 9.3
R13397 vss.n3352 vss.n3351 9.3
R13398 vss.n3367 vss.n3366 9.3
R13399 vss.n3365 vss.n3364 9.3
R13400 vss.n3364 vss.n3363 9.3
R13401 vss.n3363 vss.n3362 9.3
R13402 vss.n3380 vss.n3379 9.3
R13403 vss.n3379 vss.n3378 9.3
R13404 vss.n3378 vss.n3377 9.3
R13405 vss.n3384 vss.n3383 9.3
R13406 vss.n3382 vss.n3381 9.3
R13407 vss.n3397 vss.n3396 9.3
R13408 vss.n3395 vss.n3394 9.3
R13409 vss.n3394 vss.n3393 9.3
R13410 vss.n3393 vss.n3392 9.3
R13411 vss.n3410 vss.n3409 9.3
R13412 vss.n3409 vss.n3408 9.3
R13413 vss.n3408 vss.n3407 9.3
R13414 vss.n3414 vss.n3413 9.3
R13415 vss.n3412 vss.n3411 9.3
R13416 vss.n3441 vss.n3440 9.3
R13417 vss.n3439 vss.n3438 9.3
R13418 vss.n3446 vss.n3445 9.3
R13419 vss.n3444 vss.n3443 9.3
R13420 vss.n3449 vss.n3448 9.3
R13421 vss.n3424 vss.n3423 9.3
R13422 vss.n3423 vss.n3422 9.3
R13423 vss.n3431 vss.n3430 9.3
R13424 vss.n3435 vss.n3434 9.3
R13425 vss.n3433 vss.n3432 9.3
R13426 vss.n3488 vss.n3487 9.3
R13427 vss.n3487 vss.n3486 9.3
R13428 vss.n15172 vss.n15171 9.3
R13429 vss.n15209 vss.n15208 9.3
R13430 vss.n15208 vss.n15207 9.3
R13431 vss.n15207 vss.n15206 9.3
R13432 vss.n15189 vss.n15188 9.3
R13433 vss.n15188 vss.n15187 9.3
R13434 vss.n15187 vss.n15186 9.3
R13435 vss.n3465 vss.n3464 9.3
R13436 vss.n3464 vss.n3463 9.3
R13437 vss.n3476 vss.n3475 9.3
R13438 vss.n3475 vss.n3474 9.3
R13439 vss.n15170 vss.n15169 9.3
R13440 vss.n15168 vss.n15167 9.3
R13441 vss.n15167 vss.n15166 9.3
R13442 vss.n15166 vss.n15165 9.3
R13443 vss.n16236 vss.n16235 9.3
R13444 vss.n16235 vss.n16234 9.3
R13445 vss.n16222 vss.n16221 9.3
R13446 vss.n16221 vss.n16220 9.3
R13447 vss.n16208 vss.n16207 9.3
R13448 vss.n16207 vss.n16206 9.3
R13449 vss.n16194 vss.n16193 9.3
R13450 vss.n16193 vss.n16192 9.3
R13451 vss.n16170 vss.n16169 9.3
R13452 vss.n16169 vss.n16168 9.3
R13453 vss.n16156 vss.n16155 9.3
R13454 vss.n16155 vss.n16154 9.3
R13455 vss.n16142 vss.n16141 9.3
R13456 vss.n16141 vss.n16140 9.3
R13457 vss.n16128 vss.n16127 9.3
R13458 vss.n16127 vss.n16126 9.3
R13459 vss.n16114 vss.n16113 9.3
R13460 vss.n16113 vss.n16112 9.3
R13461 vss.n16100 vss.n16099 9.3
R13462 vss.n16099 vss.n16098 9.3
R13463 vss.n16086 vss.n16085 9.3
R13464 vss.n16085 vss.n16084 9.3
R13465 vss.n16072 vss.n16071 9.3
R13466 vss.n16071 vss.n16070 9.3
R13467 vss.n16056 vss.n16055 9.3
R13468 vss.n16055 vss.n16054 9.3
R13469 vss.n16042 vss.n16041 9.3
R13470 vss.n16041 vss.n16040 9.3
R13471 vss.n16028 vss.n16027 9.3
R13472 vss.n16027 vss.n16026 9.3
R13473 vss.n16014 vss.n16013 9.3
R13474 vss.n16013 vss.n16012 9.3
R13475 vss.n16000 vss.n15999 9.3
R13476 vss.n15999 vss.n15998 9.3
R13477 vss.n15986 vss.n15985 9.3
R13478 vss.n15985 vss.n15984 9.3
R13479 vss.n15972 vss.n15971 9.3
R13480 vss.n15971 vss.n15970 9.3
R13481 vss.n15958 vss.n15957 9.3
R13482 vss.n15957 vss.n15956 9.3
R13483 vss.n15934 vss.n15933 9.3
R13484 vss.n15933 vss.n15932 9.3
R13485 vss.n15920 vss.n15919 9.3
R13486 vss.n15919 vss.n15918 9.3
R13487 vss.n15906 vss.n15905 9.3
R13488 vss.n15905 vss.n15904 9.3
R13489 vss.n15892 vss.n15891 9.3
R13490 vss.n15891 vss.n15890 9.3
R13491 vss.n15330 vss.n15329 9.3
R13492 vss.n15344 vss.n15343 9.3
R13493 vss.n15359 vss.n15358 9.3
R13494 vss.n15373 vss.n15372 9.3
R13495 vss.n15387 vss.n15386 9.3
R13496 vss.n15401 vss.n15400 9.3
R13497 vss.n15415 vss.n15414 9.3
R13498 vss.n15434 vss.n15433 9.3
R13499 vss.n15448 vss.n15447 9.3
R13500 vss.n15462 vss.n15461 9.3
R13501 vss.n15476 vss.n15475 9.3
R13502 vss.n15490 vss.n15489 9.3
R13503 vss.n15504 vss.n15503 9.3
R13504 vss.n15518 vss.n15517 9.3
R13505 vss.n15532 vss.n15531 9.3
R13506 vss.n15553 vss.n15552 9.3
R13507 vss.n15567 vss.n15566 9.3
R13508 vss.n15581 vss.n15580 9.3
R13509 vss.n15595 vss.n15594 9.3
R13510 vss.n15609 vss.n15608 9.3
R13511 vss.n15623 vss.n15622 9.3
R13512 vss.n15637 vss.n15636 9.3
R13513 vss.n15651 vss.n15650 9.3
R13514 vss.n15670 vss.n15669 9.3
R13515 vss.n15684 vss.n15683 9.3
R13516 vss.n15698 vss.n15697 9.3
R13517 vss.n15712 vss.n15711 9.3
R13518 vss.n15726 vss.n15725 9.3
R13519 vss.n15740 vss.n15739 9.3
R13520 vss.n15754 vss.n15753 9.3
R13521 vss.n15768 vss.n15767 9.3
R13522 vss.n15823 vss.n15822 9.3
R13523 vss.n15837 vss.n15836 9.3
R13524 vss.n15851 vss.n15850 9.3
R13525 vss.n15863 vss.n15862 9.3
R13526 vss.n15305 vss.n15304 9.3
R13527 vss.n15248 vss.n15247 9.3
R13528 vss.n15247 vss.n15246 9.3
R13529 vss.n15238 vss.n15237 9.3
R13530 vss.n15237 vss.n15236 9.3
R13531 vss.n15321 vss.n15320 9.3
R13532 vss.n15320 vss.n15319 9.3
R13533 vss.n15226 vss.n15225 9.3
R13534 vss.n15225 vss.n15224 9.3
R13535 vss.n15328 vss.n15327 9.3
R13536 vss.n15340 vss.n15339 9.3
R13537 vss.n15339 vss.n15338 9.3
R13538 vss.n15338 vss.n15337 9.3
R13539 vss.n15342 vss.n15341 9.3
R13540 vss.n15354 vss.n15353 9.3
R13541 vss.n15353 vss.n15352 9.3
R13542 vss.n15352 vss.n15351 9.3
R13543 vss.n15356 vss.n15355 9.3
R13544 vss.n15369 vss.n15368 9.3
R13545 vss.n15368 vss.n15367 9.3
R13546 vss.n15367 vss.n15366 9.3
R13547 vss.n15371 vss.n15370 9.3
R13548 vss.n15383 vss.n15382 9.3
R13549 vss.n15382 vss.n15381 9.3
R13550 vss.n15381 vss.n15380 9.3
R13551 vss.n15385 vss.n15384 9.3
R13552 vss.n15397 vss.n15396 9.3
R13553 vss.n15396 vss.n15395 9.3
R13554 vss.n15395 vss.n15394 9.3
R13555 vss.n15399 vss.n15398 9.3
R13556 vss.n15411 vss.n15410 9.3
R13557 vss.n15410 vss.n15409 9.3
R13558 vss.n15409 vss.n15408 9.3
R13559 vss.n15413 vss.n15412 9.3
R13560 vss.n15422 vss.n15421 9.3
R13561 vss.n15436 vss.n15435 9.3
R13562 vss.n15432 vss.n15431 9.3
R13563 vss.n15431 vss.n15430 9.3
R13564 vss.n15430 vss.n15429 9.3
R13565 vss.n15450 vss.n15449 9.3
R13566 vss.n15446 vss.n15445 9.3
R13567 vss.n15445 vss.n15444 9.3
R13568 vss.n15444 vss.n15443 9.3
R13569 vss.n15464 vss.n15463 9.3
R13570 vss.n15460 vss.n15459 9.3
R13571 vss.n15459 vss.n15458 9.3
R13572 vss.n15458 vss.n15457 9.3
R13573 vss.n15478 vss.n15477 9.3
R13574 vss.n15474 vss.n15473 9.3
R13575 vss.n15473 vss.n15472 9.3
R13576 vss.n15472 vss.n15471 9.3
R13577 vss.n15492 vss.n15491 9.3
R13578 vss.n15488 vss.n15487 9.3
R13579 vss.n15487 vss.n15486 9.3
R13580 vss.n15486 vss.n15485 9.3
R13581 vss.n15506 vss.n15505 9.3
R13582 vss.n15502 vss.n15501 9.3
R13583 vss.n15501 vss.n15500 9.3
R13584 vss.n15500 vss.n15499 9.3
R13585 vss.n15520 vss.n15519 9.3
R13586 vss.n15516 vss.n15515 9.3
R13587 vss.n15515 vss.n15514 9.3
R13588 vss.n15514 vss.n15513 9.3
R13589 vss.n15534 vss.n15533 9.3
R13590 vss.n15530 vss.n15529 9.3
R13591 vss.n15529 vss.n15528 9.3
R13592 vss.n15528 vss.n15527 9.3
R13593 vss.n15546 vss.n15545 9.3
R13594 vss.n15545 vss.n15544 9.3
R13595 vss.n15551 vss.n15550 9.3
R13596 vss.n15563 vss.n15562 9.3
R13597 vss.n15562 vss.n15561 9.3
R13598 vss.n15561 vss.n15560 9.3
R13599 vss.n15565 vss.n15564 9.3
R13600 vss.n15577 vss.n15576 9.3
R13601 vss.n15576 vss.n15575 9.3
R13602 vss.n15575 vss.n15574 9.3
R13603 vss.n15579 vss.n15578 9.3
R13604 vss.n15591 vss.n15590 9.3
R13605 vss.n15590 vss.n15589 9.3
R13606 vss.n15589 vss.n15588 9.3
R13607 vss.n15593 vss.n15592 9.3
R13608 vss.n15605 vss.n15604 9.3
R13609 vss.n15604 vss.n15603 9.3
R13610 vss.n15603 vss.n15602 9.3
R13611 vss.n15607 vss.n15606 9.3
R13612 vss.n15619 vss.n15618 9.3
R13613 vss.n15618 vss.n15617 9.3
R13614 vss.n15617 vss.n15616 9.3
R13615 vss.n15621 vss.n15620 9.3
R13616 vss.n15633 vss.n15632 9.3
R13617 vss.n15632 vss.n15631 9.3
R13618 vss.n15631 vss.n15630 9.3
R13619 vss.n15635 vss.n15634 9.3
R13620 vss.n15647 vss.n15646 9.3
R13621 vss.n15646 vss.n15645 9.3
R13622 vss.n15645 vss.n15644 9.3
R13623 vss.n15649 vss.n15648 9.3
R13624 vss.n15658 vss.n15657 9.3
R13625 vss.n15672 vss.n15671 9.3
R13626 vss.n15668 vss.n15667 9.3
R13627 vss.n15667 vss.n15666 9.3
R13628 vss.n15666 vss.n15665 9.3
R13629 vss.n15686 vss.n15685 9.3
R13630 vss.n15682 vss.n15681 9.3
R13631 vss.n15681 vss.n15680 9.3
R13632 vss.n15680 vss.n15679 9.3
R13633 vss.n15700 vss.n15699 9.3
R13634 vss.n15696 vss.n15695 9.3
R13635 vss.n15695 vss.n15694 9.3
R13636 vss.n15694 vss.n15693 9.3
R13637 vss.n15714 vss.n15713 9.3
R13638 vss.n15710 vss.n15709 9.3
R13639 vss.n15709 vss.n15708 9.3
R13640 vss.n15708 vss.n15707 9.3
R13641 vss.n15728 vss.n15727 9.3
R13642 vss.n15724 vss.n15723 9.3
R13643 vss.n15723 vss.n15722 9.3
R13644 vss.n15722 vss.n15721 9.3
R13645 vss.n15742 vss.n15741 9.3
R13646 vss.n15738 vss.n15737 9.3
R13647 vss.n15737 vss.n15736 9.3
R13648 vss.n15736 vss.n15735 9.3
R13649 vss.n15756 vss.n15755 9.3
R13650 vss.n15752 vss.n15751 9.3
R13651 vss.n15751 vss.n15750 9.3
R13652 vss.n15750 vss.n15749 9.3
R13653 vss.n15770 vss.n15769 9.3
R13654 vss.n15766 vss.n15765 9.3
R13655 vss.n15765 vss.n15764 9.3
R13656 vss.n15764 vss.n15763 9.3
R13657 vss.n15780 vss.n15779 9.3
R13658 vss.n15779 vss.n15778 9.3
R13659 vss.n15792 vss.n15791 9.3
R13660 vss.n15791 vss.n15790 9.3
R13661 vss.n15804 vss.n15803 9.3
R13662 vss.n15803 vss.n15802 9.3
R13663 vss.n15814 vss.n15813 9.3
R13664 vss.n15813 vss.n15812 9.3
R13665 vss.n15821 vss.n15820 9.3
R13666 vss.n15833 vss.n15832 9.3
R13667 vss.n15832 vss.n15831 9.3
R13668 vss.n15831 vss.n15830 9.3
R13669 vss.n15835 vss.n15834 9.3
R13670 vss.n15847 vss.n15846 9.3
R13671 vss.n15846 vss.n15845 9.3
R13672 vss.n15845 vss.n15844 9.3
R13673 vss.n15849 vss.n15848 9.3
R13674 vss.n15861 vss.n15860 9.3
R13675 vss.n15860 vss.n15859 9.3
R13676 vss.n15859 vss.n15858 9.3
R13677 vss.n15872 vss.n15871 9.3
R13678 vss.n15871 vss.n15870 9.3
R13679 vss.n16286 vss.n16285 9.3
R13680 vss.n16272 vss.n16271 9.3
R13681 vss.n15261 vss.n15260 9.3
R13682 vss.n15275 vss.n15274 9.3
R13683 vss.n15289 vss.n15288 9.3
R13684 vss.n15303 vss.n15302 9.3
R13685 vss.n16284 vss.n16283 9.3
R13686 vss.n16270 vss.n16269 9.3
R13687 vss.n16282 vss.n16281 9.3
R13688 vss.n16281 vss.n16280 9.3
R13689 vss.n16280 vss.n16279 9.3
R13690 vss.n15263 vss.n15262 9.3
R13691 vss.n15259 vss.n15258 9.3
R13692 vss.n15258 vss.n15257 9.3
R13693 vss.n15257 vss.n15256 9.3
R13694 vss.n15277 vss.n15276 9.3
R13695 vss.n15273 vss.n15272 9.3
R13696 vss.n15272 vss.n15271 9.3
R13697 vss.n15271 vss.n15270 9.3
R13698 vss.n15291 vss.n15290 9.3
R13699 vss.n15287 vss.n15286 9.3
R13700 vss.n15286 vss.n15285 9.3
R13701 vss.n15285 vss.n15284 9.3
R13702 vss.n15301 vss.n15300 9.3
R13703 vss.n15300 vss.n15299 9.3
R13704 vss.n15299 vss.n15298 9.3
R13705 vss.n16293 vss.n16292 9.3
R13706 vss.n16292 vss.n16291 9.3
R13707 vss.n16291 vss.n16290 9.3
R13708 vss.n16657 vss.n16656 9.3
R13709 vss.n16656 vss.n16655 9.3
R13710 vss.n16655 vss.n16654 9.3
R13711 vss.n16633 vss.n16632 9.3
R13712 vss.n16596 vss.n16595 9.3
R13713 vss.n16582 vss.n16581 9.3
R13714 vss.n16568 vss.n16567 9.3
R13715 vss.n16554 vss.n16553 9.3
R13716 vss.n16540 vss.n16539 9.3
R13717 vss.n16526 vss.n16525 9.3
R13718 vss.n16512 vss.n16511 9.3
R13719 vss.n16498 vss.n16497 9.3
R13720 vss.n16467 vss.n16466 9.3
R13721 vss.n16439 vss.n16438 9.3
R13722 vss.n16411 vss.n16410 9.3
R13723 vss.n16383 vss.n16382 9.3
R13724 vss.n16360 vss.n16359 9.3
R13725 vss.n16346 vss.n16345 9.3
R13726 vss.n16332 vss.n16331 9.3
R13727 vss.n16318 vss.n16317 9.3
R13728 vss.n16304 vss.n16303 9.3
R13729 vss.n16316 vss.n16315 9.3
R13730 vss.n16315 vss.n16314 9.3
R13731 vss.n16314 vss.n16313 9.3
R13732 vss.n16306 vss.n16305 9.3
R13733 vss.n16320 vss.n16319 9.3
R13734 vss.n16330 vss.n16329 9.3
R13735 vss.n16329 vss.n16328 9.3
R13736 vss.n16328 vss.n16327 9.3
R13737 vss.n16344 vss.n16343 9.3
R13738 vss.n16343 vss.n16342 9.3
R13739 vss.n16342 vss.n16341 9.3
R13740 vss.n16334 vss.n16333 9.3
R13741 vss.n16348 vss.n16347 9.3
R13742 vss.n16358 vss.n16357 9.3
R13743 vss.n16357 vss.n16356 9.3
R13744 vss.n16356 vss.n16355 9.3
R13745 vss.n16369 vss.n16368 9.3
R13746 vss.n16362 vss.n16361 9.3
R13747 vss.n16381 vss.n16380 9.3
R13748 vss.n16379 vss.n16378 9.3
R13749 vss.n16378 vss.n16377 9.3
R13750 vss.n16377 vss.n16376 9.3
R13751 vss.n16393 vss.n16392 9.3
R13752 vss.n16392 vss.n16391 9.3
R13753 vss.n16391 vss.n16390 9.3
R13754 vss.n16397 vss.n16396 9.3
R13755 vss.n16395 vss.n16394 9.3
R13756 vss.n16409 vss.n16408 9.3
R13757 vss.n16407 vss.n16406 9.3
R13758 vss.n16406 vss.n16405 9.3
R13759 vss.n16405 vss.n16404 9.3
R13760 vss.n16421 vss.n16420 9.3
R13761 vss.n16420 vss.n16419 9.3
R13762 vss.n16419 vss.n16418 9.3
R13763 vss.n16425 vss.n16424 9.3
R13764 vss.n16423 vss.n16422 9.3
R13765 vss.n16437 vss.n16436 9.3
R13766 vss.n16435 vss.n16434 9.3
R13767 vss.n16434 vss.n16433 9.3
R13768 vss.n16433 vss.n16432 9.3
R13769 vss.n16449 vss.n16448 9.3
R13770 vss.n16448 vss.n16447 9.3
R13771 vss.n16447 vss.n16446 9.3
R13772 vss.n16453 vss.n16452 9.3
R13773 vss.n16451 vss.n16450 9.3
R13774 vss.n16465 vss.n16464 9.3
R13775 vss.n16463 vss.n16462 9.3
R13776 vss.n16462 vss.n16461 9.3
R13777 vss.n16461 vss.n16460 9.3
R13778 vss.n16477 vss.n16476 9.3
R13779 vss.n16476 vss.n16475 9.3
R13780 vss.n16475 vss.n16474 9.3
R13781 vss.n16481 vss.n16480 9.3
R13782 vss.n16479 vss.n16478 9.3
R13783 vss.n16493 vss.n16492 9.3
R13784 vss.n16492 vss.n16491 9.3
R13785 vss.n16510 vss.n16509 9.3
R13786 vss.n16509 vss.n16508 9.3
R13787 vss.n16508 vss.n16507 9.3
R13788 vss.n16500 vss.n16499 9.3
R13789 vss.n16514 vss.n16513 9.3
R13790 vss.n16524 vss.n16523 9.3
R13791 vss.n16523 vss.n16522 9.3
R13792 vss.n16522 vss.n16521 9.3
R13793 vss.n16538 vss.n16537 9.3
R13794 vss.n16537 vss.n16536 9.3
R13795 vss.n16536 vss.n16535 9.3
R13796 vss.n16528 vss.n16527 9.3
R13797 vss.n16542 vss.n16541 9.3
R13798 vss.n16552 vss.n16551 9.3
R13799 vss.n16551 vss.n16550 9.3
R13800 vss.n16550 vss.n16549 9.3
R13801 vss.n16566 vss.n16565 9.3
R13802 vss.n16565 vss.n16564 9.3
R13803 vss.n16564 vss.n16563 9.3
R13804 vss.n16556 vss.n16555 9.3
R13805 vss.n16570 vss.n16569 9.3
R13806 vss.n16580 vss.n16579 9.3
R13807 vss.n16579 vss.n16578 9.3
R13808 vss.n16578 vss.n16577 9.3
R13809 vss.n16594 vss.n16593 9.3
R13810 vss.n16593 vss.n16592 9.3
R13811 vss.n16592 vss.n16591 9.3
R13812 vss.n16584 vss.n16583 9.3
R13813 vss.n16598 vss.n16597 9.3
R13814 vss.n16605 vss.n16604 9.3
R13815 vss.n16615 vss.n16614 9.3
R13816 vss.n16614 vss.n16613 9.3
R13817 vss.n16613 vss.n16612 9.3
R13818 vss.n16619 vss.n16618 9.3
R13819 vss.n16617 vss.n16616 9.3
R13820 vss.n16631 vss.n16630 9.3
R13821 vss.n16629 vss.n16628 9.3
R13822 vss.n16628 vss.n16627 9.3
R13823 vss.n16627 vss.n16626 9.3
R13824 vss.n16643 vss.n16642 9.3
R13825 vss.n16642 vss.n16641 9.3
R13826 vss.n16641 vss.n16640 9.3
R13827 vss.n16647 vss.n16646 9.3
R13828 vss.n16645 vss.n16644 9.3
R13829 vss.n16659 vss.n16658 9.3
R13830 vss.n16661 vss.n16660 9.3
R13831 vss.n22081 vss.n22080 9.3
R13832 vss.n22080 vss.n22079 9.3
R13833 vss.n22097 vss.n22096 9.3
R13834 vss.n22096 vss.n22095 9.3
R13835 vss.n22111 vss.n22110 9.3
R13836 vss.n22110 vss.n22109 9.3
R13837 vss.n22125 vss.n22124 9.3
R13838 vss.n22124 vss.n22123 9.3
R13839 vss.n22139 vss.n22138 9.3
R13840 vss.n22138 vss.n22137 9.3
R13841 vss.n22153 vss.n22152 9.3
R13842 vss.n22152 vss.n22151 9.3
R13843 vss.n22167 vss.n22166 9.3
R13844 vss.n22166 vss.n22165 9.3
R13845 vss.n17395 vss.n17394 9.3
R13846 vss.n17394 vss.n17393 9.3
R13847 vss.n17384 vss.n17383 9.3
R13848 vss.n17383 vss.n17382 9.3
R13849 vss.n22186 vss.n22185 9.3
R13850 vss.n22185 vss.n22184 9.3
R13851 vss.n22200 vss.n22199 9.3
R13852 vss.n22199 vss.n22198 9.3
R13853 vss.n22214 vss.n22213 9.3
R13854 vss.n22213 vss.n22212 9.3
R13855 vss.n22228 vss.n22227 9.3
R13856 vss.n22227 vss.n22226 9.3
R13857 vss.n22242 vss.n22241 9.3
R13858 vss.n22241 vss.n22240 9.3
R13859 vss.n22256 vss.n22255 9.3
R13860 vss.n22255 vss.n22254 9.3
R13861 vss.n22272 vss.n22271 9.3
R13862 vss.n22271 vss.n22270 9.3
R13863 vss.n22291 vss.n22290 9.3
R13864 vss.n22290 vss.n22289 9.3
R13865 vss.n22305 vss.n22304 9.3
R13866 vss.n22304 vss.n22303 9.3
R13867 vss.n22319 vss.n22318 9.3
R13868 vss.n22318 vss.n22317 9.3
R13869 vss.n22333 vss.n22332 9.3
R13870 vss.n22332 vss.n22331 9.3
R13871 vss.n22347 vss.n22346 9.3
R13872 vss.n22346 vss.n22345 9.3
R13873 vss.n22361 vss.n22360 9.3
R13874 vss.n22360 vss.n22359 9.3
R13875 vss.n22375 vss.n22374 9.3
R13876 vss.n22374 vss.n22373 9.3
R13877 vss.n17373 vss.n17372 9.3
R13878 vss.n17372 vss.n17371 9.3
R13879 vss.n17362 vss.n17361 9.3
R13880 vss.n17361 vss.n17360 9.3
R13881 vss.n22394 vss.n22393 9.3
R13882 vss.n22393 vss.n22392 9.3
R13883 vss.n22408 vss.n22407 9.3
R13884 vss.n22407 vss.n22406 9.3
R13885 vss.n22422 vss.n22421 9.3
R13886 vss.n22421 vss.n22420 9.3
R13887 vss.n22436 vss.n22435 9.3
R13888 vss.n22435 vss.n22434 9.3
R13889 vss.n22450 vss.n22449 9.3
R13890 vss.n22449 vss.n22448 9.3
R13891 vss.n22464 vss.n22463 9.3
R13892 vss.n22463 vss.n22462 9.3
R13893 vss.n22480 vss.n22479 9.3
R13894 vss.n22479 vss.n22478 9.3
R13895 vss.n22499 vss.n22498 9.3
R13896 vss.n22498 vss.n22497 9.3
R13897 vss.n22513 vss.n22512 9.3
R13898 vss.n22512 vss.n22511 9.3
R13899 vss.n22527 vss.n22526 9.3
R13900 vss.n22526 vss.n22525 9.3
R13901 vss.n22541 vss.n22540 9.3
R13902 vss.n22540 vss.n22539 9.3
R13903 vss.n22555 vss.n22554 9.3
R13904 vss.n22554 vss.n22553 9.3
R13905 vss.n22569 vss.n22568 9.3
R13906 vss.n22568 vss.n22567 9.3
R13907 vss.n22583 vss.n22582 9.3
R13908 vss.n22582 vss.n22581 9.3
R13909 vss.n17351 vss.n17350 9.3
R13910 vss.n17350 vss.n17349 9.3
R13911 vss.n17340 vss.n17339 9.3
R13912 vss.n17339 vss.n17338 9.3
R13913 vss.n22602 vss.n22601 9.3
R13914 vss.n22601 vss.n22600 9.3
R13915 vss.n22616 vss.n22615 9.3
R13916 vss.n22615 vss.n22614 9.3
R13917 vss.n22630 vss.n22629 9.3
R13918 vss.n22629 vss.n22628 9.3
R13919 vss.n22644 vss.n22643 9.3
R13920 vss.n22643 vss.n22642 9.3
R13921 vss.n22658 vss.n22657 9.3
R13922 vss.n22657 vss.n22656 9.3
R13923 vss.n22672 vss.n22671 9.3
R13924 vss.n22671 vss.n22670 9.3
R13925 vss.n22688 vss.n22687 9.3
R13926 vss.n22687 vss.n22686 9.3
R13927 vss.n22707 vss.n22706 9.3
R13928 vss.n22706 vss.n22705 9.3
R13929 vss.n22721 vss.n22720 9.3
R13930 vss.n22720 vss.n22719 9.3
R13931 vss.n22735 vss.n22734 9.3
R13932 vss.n22734 vss.n22733 9.3
R13933 vss.n22749 vss.n22748 9.3
R13934 vss.n22748 vss.n22747 9.3
R13935 vss.n243 vss.n242 9.3
R13936 vss.n188 vss.n187 9.3
R13937 vss.n158 vss.n157 9.3
R13938 vss.n156 vss.n155 9.3
R13939 vss.n154 vss.n153 9.3
R13940 vss.n153 vss.n152 9.3
R13941 vss.n152 vss.n151 9.3
R13942 vss.n169 vss.n168 9.3
R13943 vss.n168 vss.n167 9.3
R13944 vss.n167 vss.n166 9.3
R13945 vss.n173 vss.n172 9.3
R13946 vss.n171 vss.n170 9.3
R13947 vss.n186 vss.n185 9.3
R13948 vss.n184 vss.n183 9.3
R13949 vss.n183 vss.n182 9.3
R13950 vss.n182 vss.n181 9.3
R13951 vss.n199 vss.n198 9.3
R13952 vss.n198 vss.n197 9.3
R13953 vss.n197 vss.n196 9.3
R13954 vss.n203 vss.n202 9.3
R13955 vss.n201 vss.n200 9.3
R13956 vss.n221 vss.n220 9.3
R13957 vss.n220 vss.n219 9.3
R13958 vss.n219 vss.n218 9.3
R13959 vss.n241 vss.n240 9.3
R13960 vss.n240 vss.n239 9.3
R13961 vss.n239 vss.n238 9.3
R13962 vss.n258 vss.n257 9.3
R13963 vss.n257 vss.n256 9.3
R13964 vss.n256 vss.n255 9.3
R13965 vss.n245 vss.n244 9.3
R13966 vss.n22859 vss.n22858 9.3
R13967 vss.n22889 vss.n22888 9.3
R13968 vss.n22919 vss.n22918 9.3
R13969 vss.n22923 vss.n22922 9.3
R13970 vss.n22940 vss.n22939 9.3
R13971 vss.n22956 vss.n22955 9.3
R13972 vss.n22972 vss.n22971 9.3
R13973 vss.n22988 vss.n22987 9.3
R13974 vss.n23004 vss.n23003 9.3
R13975 vss.n23020 vss.n23019 9.3
R13976 vss.n23040 vss.n23039 9.3
R13977 vss.n23047 vss.n23046 9.3
R13978 vss.n23083 vss.n23082 9.3
R13979 vss.n23115 vss.n23114 9.3
R13980 vss.n23148 vss.n23147 9.3
R13981 vss.n23168 vss.n23167 9.3
R13982 vss.n23184 vss.n23183 9.3
R13983 vss.n23200 vss.n23199 9.3
R13984 vss.n23216 vss.n23215 9.3
R13985 vss.n23232 vss.n23231 9.3
R13986 vss.n23249 vss.n23248 9.3
R13987 vss.n23265 vss.n23264 9.3
R13988 vss.n23285 vss.n23284 9.3
R13989 vss.n23311 vss.n23310 9.3
R13990 vss.n23343 vss.n23342 9.3
R13991 vss.n23375 vss.n23374 9.3
R13992 vss.n23407 vss.n23406 9.3
R13993 vss.n23411 vss.n23410 9.3
R13994 vss.n1297 vss.n1296 9.3
R13995 vss.n1280 vss.n1279 9.3
R13996 vss.n1264 vss.n1263 9.3
R13997 vss.n1248 vss.n1247 9.3
R13998 vss.n1232 vss.n1231 9.3
R13999 vss.n1216 vss.n1215 9.3
R14000 vss.n1196 vss.n1195 9.3
R14001 vss.n1190 vss.n1189 9.3
R14002 vss.n1153 vss.n1152 9.3
R14003 vss.n1121 vss.n1120 9.3
R14004 vss.n1089 vss.n1088 9.3
R14005 vss.n1068 vss.n1067 9.3
R14006 vss.n1052 vss.n1051 9.3
R14007 vss.n1036 vss.n1035 9.3
R14008 vss.n1020 vss.n1019 9.3
R14009 vss.n1004 vss.n1003 9.3
R14010 vss.n988 vss.n987 9.3
R14011 vss.n972 vss.n971 9.3
R14012 vss.n951 vss.n950 9.3
R14013 vss.n925 vss.n924 9.3
R14014 vss.n893 vss.n892 9.3
R14015 vss.n861 vss.n860 9.3
R14016 vss.n828 vss.n827 9.3
R14017 vss.n824 vss.n823 9.3
R14018 vss.n808 vss.n807 9.3
R14019 vss.n792 vss.n791 9.3
R14020 vss.n776 vss.n775 9.3
R14021 vss.n760 vss.n759 9.3
R14022 vss.n743 vss.n742 9.3
R14023 vss.n727 vss.n726 9.3
R14024 vss.n707 vss.n706 9.3
R14025 vss.n701 vss.n700 9.3
R14026 vss.n665 vss.n664 9.3
R14027 vss.n632 vss.n631 9.3
R14028 vss.n600 vss.n599 9.3
R14029 vss.n580 vss.n579 9.3
R14030 vss.n564 vss.n563 9.3
R14031 vss.n547 vss.n546 9.3
R14032 vss.n531 vss.n530 9.3
R14033 vss.n515 vss.n514 9.3
R14034 vss.n499 vss.n498 9.3
R14035 vss.n483 vss.n482 9.3
R14036 vss.n463 vss.n462 9.3
R14037 vss.n436 vss.n435 9.3
R14038 vss.n404 vss.n403 9.3
R14039 vss.n372 vss.n371 9.3
R14040 vss.n339 vss.n338 9.3
R14041 vss.n335 vss.n334 9.3
R14042 vss.n320 vss.n319 9.3
R14043 vss.n305 vss.n304 9.3
R14044 vss.n290 vss.n289 9.3
R14045 vss.n275 vss.n274 9.3
R14046 vss.n260 vss.n259 9.3
R14047 vss.n262 vss.n261 9.3
R14048 vss.n273 vss.n272 9.3
R14049 vss.n272 vss.n271 9.3
R14050 vss.n271 vss.n270 9.3
R14051 vss.n288 vss.n287 9.3
R14052 vss.n287 vss.n286 9.3
R14053 vss.n286 vss.n285 9.3
R14054 vss.n277 vss.n276 9.3
R14055 vss.n292 vss.n291 9.3
R14056 vss.n303 vss.n302 9.3
R14057 vss.n302 vss.n301 9.3
R14058 vss.n301 vss.n300 9.3
R14059 vss.n318 vss.n317 9.3
R14060 vss.n317 vss.n316 9.3
R14061 vss.n316 vss.n315 9.3
R14062 vss.n307 vss.n306 9.3
R14063 vss.n322 vss.n321 9.3
R14064 vss.n333 vss.n332 9.3
R14065 vss.n332 vss.n331 9.3
R14066 vss.n331 vss.n330 9.3
R14067 vss.n110 vss.n109 9.3
R14068 vss.n109 vss.n108 9.3
R14069 vss.n98 vss.n97 9.3
R14070 vss.n97 vss.n96 9.3
R14071 vss.n352 vss.n351 9.3
R14072 vss.n351 vss.n350 9.3
R14073 vss.n350 vss.n349 9.3
R14074 vss.n356 vss.n355 9.3
R14075 vss.n354 vss.n353 9.3
R14076 vss.n370 vss.n369 9.3
R14077 vss.n368 vss.n367 9.3
R14078 vss.n367 vss.n366 9.3
R14079 vss.n366 vss.n365 9.3
R14080 vss.n384 vss.n383 9.3
R14081 vss.n383 vss.n382 9.3
R14082 vss.n382 vss.n381 9.3
R14083 vss.n388 vss.n387 9.3
R14084 vss.n386 vss.n385 9.3
R14085 vss.n402 vss.n401 9.3
R14086 vss.n400 vss.n399 9.3
R14087 vss.n399 vss.n398 9.3
R14088 vss.n398 vss.n397 9.3
R14089 vss.n416 vss.n415 9.3
R14090 vss.n415 vss.n414 9.3
R14091 vss.n414 vss.n413 9.3
R14092 vss.n420 vss.n419 9.3
R14093 vss.n418 vss.n417 9.3
R14094 vss.n434 vss.n433 9.3
R14095 vss.n432 vss.n431 9.3
R14096 vss.n431 vss.n430 9.3
R14097 vss.n430 vss.n429 9.3
R14098 vss.n452 vss.n451 9.3
R14099 vss.n451 vss.n450 9.3
R14100 vss.n450 vss.n449 9.3
R14101 vss.n456 vss.n455 9.3
R14102 vss.n454 vss.n453 9.3
R14103 vss.n481 vss.n480 9.3
R14104 vss.n480 vss.n479 9.3
R14105 vss.n479 vss.n478 9.3
R14106 vss.n465 vss.n464 9.3
R14107 vss.n485 vss.n484 9.3
R14108 vss.n497 vss.n496 9.3
R14109 vss.n496 vss.n495 9.3
R14110 vss.n495 vss.n494 9.3
R14111 vss.n513 vss.n512 9.3
R14112 vss.n512 vss.n511 9.3
R14113 vss.n511 vss.n510 9.3
R14114 vss.n501 vss.n500 9.3
R14115 vss.n517 vss.n516 9.3
R14116 vss.n529 vss.n528 9.3
R14117 vss.n528 vss.n527 9.3
R14118 vss.n527 vss.n526 9.3
R14119 vss.n545 vss.n544 9.3
R14120 vss.n544 vss.n543 9.3
R14121 vss.n543 vss.n542 9.3
R14122 vss.n533 vss.n532 9.3
R14123 vss.n549 vss.n548 9.3
R14124 vss.n561 vss.n560 9.3
R14125 vss.n560 vss.n559 9.3
R14126 vss.n559 vss.n558 9.3
R14127 vss.n578 vss.n577 9.3
R14128 vss.n577 vss.n576 9.3
R14129 vss.n576 vss.n575 9.3
R14130 vss.n566 vss.n565 9.3
R14131 vss.n83 vss.n82 9.3
R14132 vss.n82 vss.n81 9.3
R14133 vss.n71 vss.n70 9.3
R14134 vss.n70 vss.n69 9.3
R14135 vss.n584 vss.n583 9.3
R14136 vss.n598 vss.n597 9.3
R14137 vss.n596 vss.n595 9.3
R14138 vss.n595 vss.n594 9.3
R14139 vss.n594 vss.n593 9.3
R14140 vss.n612 vss.n611 9.3
R14141 vss.n611 vss.n610 9.3
R14142 vss.n610 vss.n609 9.3
R14143 vss.n616 vss.n615 9.3
R14144 vss.n614 vss.n613 9.3
R14145 vss.n630 vss.n629 9.3
R14146 vss.n628 vss.n627 9.3
R14147 vss.n627 vss.n626 9.3
R14148 vss.n626 vss.n625 9.3
R14149 vss.n644 vss.n643 9.3
R14150 vss.n643 vss.n642 9.3
R14151 vss.n642 vss.n641 9.3
R14152 vss.n648 vss.n647 9.3
R14153 vss.n646 vss.n645 9.3
R14154 vss.n663 vss.n662 9.3
R14155 vss.n661 vss.n660 9.3
R14156 vss.n660 vss.n659 9.3
R14157 vss.n659 vss.n658 9.3
R14158 vss.n677 vss.n676 9.3
R14159 vss.n676 vss.n675 9.3
R14160 vss.n675 vss.n674 9.3
R14161 vss.n681 vss.n680 9.3
R14162 vss.n679 vss.n678 9.3
R14163 vss.n699 vss.n698 9.3
R14164 vss.n697 vss.n696 9.3
R14165 vss.n696 vss.n695 9.3
R14166 vss.n695 vss.n694 9.3
R14167 vss.n709 vss.n708 9.3
R14168 vss.n725 vss.n724 9.3
R14169 vss.n724 vss.n723 9.3
R14170 vss.n723 vss.n722 9.3
R14171 vss.n741 vss.n740 9.3
R14172 vss.n740 vss.n739 9.3
R14173 vss.n739 vss.n738 9.3
R14174 vss.n729 vss.n728 9.3
R14175 vss.n745 vss.n744 9.3
R14176 vss.n757 vss.n756 9.3
R14177 vss.n756 vss.n755 9.3
R14178 vss.n755 vss.n754 9.3
R14179 vss.n774 vss.n773 9.3
R14180 vss.n773 vss.n772 9.3
R14181 vss.n772 vss.n771 9.3
R14182 vss.n762 vss.n761 9.3
R14183 vss.n778 vss.n777 9.3
R14184 vss.n790 vss.n789 9.3
R14185 vss.n789 vss.n788 9.3
R14186 vss.n788 vss.n787 9.3
R14187 vss.n806 vss.n805 9.3
R14188 vss.n805 vss.n804 9.3
R14189 vss.n804 vss.n803 9.3
R14190 vss.n794 vss.n793 9.3
R14191 vss.n810 vss.n809 9.3
R14192 vss.n822 vss.n821 9.3
R14193 vss.n821 vss.n820 9.3
R14194 vss.n820 vss.n819 9.3
R14195 vss.n58 vss.n57 9.3
R14196 vss.n57 vss.n56 9.3
R14197 vss.n46 vss.n45 9.3
R14198 vss.n45 vss.n44 9.3
R14199 vss.n840 vss.n839 9.3
R14200 vss.n839 vss.n838 9.3
R14201 vss.n838 vss.n837 9.3
R14202 vss.n844 vss.n843 9.3
R14203 vss.n842 vss.n841 9.3
R14204 vss.n858 vss.n857 9.3
R14205 vss.n856 vss.n855 9.3
R14206 vss.n855 vss.n854 9.3
R14207 vss.n854 vss.n853 9.3
R14208 vss.n873 vss.n872 9.3
R14209 vss.n872 vss.n871 9.3
R14210 vss.n871 vss.n870 9.3
R14211 vss.n877 vss.n876 9.3
R14212 vss.n875 vss.n874 9.3
R14213 vss.n891 vss.n890 9.3
R14214 vss.n889 vss.n888 9.3
R14215 vss.n888 vss.n887 9.3
R14216 vss.n887 vss.n886 9.3
R14217 vss.n905 vss.n904 9.3
R14218 vss.n904 vss.n903 9.3
R14219 vss.n903 vss.n902 9.3
R14220 vss.n909 vss.n908 9.3
R14221 vss.n907 vss.n906 9.3
R14222 vss.n923 vss.n922 9.3
R14223 vss.n921 vss.n920 9.3
R14224 vss.n920 vss.n919 9.3
R14225 vss.n919 vss.n918 9.3
R14226 vss.n941 vss.n940 9.3
R14227 vss.n940 vss.n939 9.3
R14228 vss.n939 vss.n938 9.3
R14229 vss.n945 vss.n944 9.3
R14230 vss.n943 vss.n942 9.3
R14231 vss.n969 vss.n968 9.3
R14232 vss.n968 vss.n967 9.3
R14233 vss.n967 vss.n966 9.3
R14234 vss.n953 vss.n952 9.3
R14235 vss.n974 vss.n973 9.3
R14236 vss.n986 vss.n985 9.3
R14237 vss.n985 vss.n984 9.3
R14238 vss.n984 vss.n983 9.3
R14239 vss.n1002 vss.n1001 9.3
R14240 vss.n1001 vss.n1000 9.3
R14241 vss.n1000 vss.n999 9.3
R14242 vss.n990 vss.n989 9.3
R14243 vss.n1006 vss.n1005 9.3
R14244 vss.n1018 vss.n1017 9.3
R14245 vss.n1017 vss.n1016 9.3
R14246 vss.n1016 vss.n1015 9.3
R14247 vss.n1034 vss.n1033 9.3
R14248 vss.n1033 vss.n1032 9.3
R14249 vss.n1032 vss.n1031 9.3
R14250 vss.n1022 vss.n1021 9.3
R14251 vss.n1038 vss.n1037 9.3
R14252 vss.n1050 vss.n1049 9.3
R14253 vss.n1049 vss.n1048 9.3
R14254 vss.n1048 vss.n1047 9.3
R14255 vss.n1066 vss.n1065 9.3
R14256 vss.n1065 vss.n1064 9.3
R14257 vss.n1064 vss.n1063 9.3
R14258 vss.n1054 vss.n1053 9.3
R14259 vss.n33 vss.n32 9.3
R14260 vss.n32 vss.n31 9.3
R14261 vss.n20 vss.n19 9.3
R14262 vss.n19 vss.n18 9.3
R14263 vss.n1073 vss.n1072 9.3
R14264 vss.n1087 vss.n1086 9.3
R14265 vss.n1085 vss.n1084 9.3
R14266 vss.n1084 vss.n1083 9.3
R14267 vss.n1083 vss.n1082 9.3
R14268 vss.n1101 vss.n1100 9.3
R14269 vss.n1100 vss.n1099 9.3
R14270 vss.n1099 vss.n1098 9.3
R14271 vss.n1105 vss.n1104 9.3
R14272 vss.n1103 vss.n1102 9.3
R14273 vss.n1119 vss.n1118 9.3
R14274 vss.n1117 vss.n1116 9.3
R14275 vss.n1116 vss.n1115 9.3
R14276 vss.n1115 vss.n1114 9.3
R14277 vss.n1133 vss.n1132 9.3
R14278 vss.n1132 vss.n1131 9.3
R14279 vss.n1131 vss.n1130 9.3
R14280 vss.n1137 vss.n1136 9.3
R14281 vss.n1135 vss.n1134 9.3
R14282 vss.n1151 vss.n1150 9.3
R14283 vss.n1149 vss.n1148 9.3
R14284 vss.n1148 vss.n1147 9.3
R14285 vss.n1147 vss.n1146 9.3
R14286 vss.n1165 vss.n1164 9.3
R14287 vss.n1164 vss.n1163 9.3
R14288 vss.n1163 vss.n1162 9.3
R14289 vss.n1169 vss.n1168 9.3
R14290 vss.n1167 vss.n1166 9.3
R14291 vss.n1188 vss.n1187 9.3
R14292 vss.n1186 vss.n1185 9.3
R14293 vss.n1185 vss.n1184 9.3
R14294 vss.n1184 vss.n1183 9.3
R14295 vss.n1198 vss.n1197 9.3
R14296 vss.n1214 vss.n1213 9.3
R14297 vss.n1213 vss.n1212 9.3
R14298 vss.n1212 vss.n1211 9.3
R14299 vss.n1230 vss.n1229 9.3
R14300 vss.n1229 vss.n1228 9.3
R14301 vss.n1228 vss.n1227 9.3
R14302 vss.n1218 vss.n1217 9.3
R14303 vss.n1234 vss.n1233 9.3
R14304 vss.n1246 vss.n1245 9.3
R14305 vss.n1245 vss.n1244 9.3
R14306 vss.n1244 vss.n1243 9.3
R14307 vss.n1262 vss.n1261 9.3
R14308 vss.n1261 vss.n1260 9.3
R14309 vss.n1260 vss.n1259 9.3
R14310 vss.n1250 vss.n1249 9.3
R14311 vss.n1266 vss.n1265 9.3
R14312 vss.n1278 vss.n1277 9.3
R14313 vss.n1277 vss.n1276 9.3
R14314 vss.n1276 vss.n1275 9.3
R14315 vss.n1295 vss.n1294 9.3
R14316 vss.n1294 vss.n1293 9.3
R14317 vss.n1293 vss.n1292 9.3
R14318 vss.n1283 vss.n1282 9.3
R14319 vss.n1299 vss.n1298 9.3
R14320 vss.n1311 vss.n1310 9.3
R14321 vss.n1310 vss.n1309 9.3
R14322 vss.n1309 vss.n1308 9.3
R14323 vss.n1322 vss.n1321 9.3
R14324 vss.n1321 vss.n1320 9.3
R14325 vss.n1334 vss.n1333 9.3
R14326 vss.n1333 vss.n1332 9.3
R14327 vss.n23405 vss.n23404 9.3
R14328 vss.n23404 vss.n23403 9.3
R14329 vss.n23403 vss.n23402 9.3
R14330 vss.n23391 vss.n23390 9.3
R14331 vss.n23393 vss.n23392 9.3
R14332 vss.n23377 vss.n23376 9.3
R14333 vss.n23389 vss.n23388 9.3
R14334 vss.n23388 vss.n23387 9.3
R14335 vss.n23387 vss.n23386 9.3
R14336 vss.n23373 vss.n23372 9.3
R14337 vss.n23372 vss.n23371 9.3
R14338 vss.n23371 vss.n23370 9.3
R14339 vss.n23359 vss.n23358 9.3
R14340 vss.n23361 vss.n23360 9.3
R14341 vss.n23345 vss.n23344 9.3
R14342 vss.n23357 vss.n23356 9.3
R14343 vss.n23356 vss.n23355 9.3
R14344 vss.n23355 vss.n23354 9.3
R14345 vss.n23341 vss.n23340 9.3
R14346 vss.n23340 vss.n23339 9.3
R14347 vss.n23339 vss.n23338 9.3
R14348 vss.n23327 vss.n23326 9.3
R14349 vss.n23329 vss.n23328 9.3
R14350 vss.n23313 vss.n23312 9.3
R14351 vss.n23325 vss.n23324 9.3
R14352 vss.n23324 vss.n23323 9.3
R14353 vss.n23323 vss.n23322 9.3
R14354 vss.n23309 vss.n23308 9.3
R14355 vss.n23308 vss.n23307 9.3
R14356 vss.n23307 vss.n23306 9.3
R14357 vss.n23291 vss.n23290 9.3
R14358 vss.n23293 vss.n23292 9.3
R14359 vss.n23281 vss.n23280 9.3
R14360 vss.n23280 vss.n23279 9.3
R14361 vss.n23279 vss.n23278 9.3
R14362 vss.n23283 vss.n23282 9.3
R14363 vss.n23263 vss.n23262 9.3
R14364 vss.n23261 vss.n23260 9.3
R14365 vss.n23260 vss.n23259 9.3
R14366 vss.n23259 vss.n23258 9.3
R14367 vss.n23244 vss.n23243 9.3
R14368 vss.n23243 vss.n23242 9.3
R14369 vss.n23242 vss.n23241 9.3
R14370 vss.n23247 vss.n23246 9.3
R14371 vss.n23230 vss.n23229 9.3
R14372 vss.n23228 vss.n23227 9.3
R14373 vss.n23227 vss.n23226 9.3
R14374 vss.n23226 vss.n23225 9.3
R14375 vss.n23212 vss.n23211 9.3
R14376 vss.n23211 vss.n23210 9.3
R14377 vss.n23210 vss.n23209 9.3
R14378 vss.n23214 vss.n23213 9.3
R14379 vss.n23198 vss.n23197 9.3
R14380 vss.n23196 vss.n23195 9.3
R14381 vss.n23195 vss.n23194 9.3
R14382 vss.n23194 vss.n23193 9.3
R14383 vss.n23180 vss.n23179 9.3
R14384 vss.n23179 vss.n23178 9.3
R14385 vss.n23178 vss.n23177 9.3
R14386 vss.n23182 vss.n23181 9.3
R14387 vss.n1348 vss.n1347 9.3
R14388 vss.n1347 vss.n1346 9.3
R14389 vss.n1360 vss.n1359 9.3
R14390 vss.n1359 vss.n1358 9.3
R14391 vss.n23164 vss.n23163 9.3
R14392 vss.n23150 vss.n23149 9.3
R14393 vss.n23162 vss.n23161 9.3
R14394 vss.n23161 vss.n23160 9.3
R14395 vss.n23160 vss.n23159 9.3
R14396 vss.n23145 vss.n23144 9.3
R14397 vss.n23144 vss.n23143 9.3
R14398 vss.n23143 vss.n23142 9.3
R14399 vss.n23131 vss.n23130 9.3
R14400 vss.n23133 vss.n23132 9.3
R14401 vss.n23117 vss.n23116 9.3
R14402 vss.n23129 vss.n23128 9.3
R14403 vss.n23128 vss.n23127 9.3
R14404 vss.n23127 vss.n23126 9.3
R14405 vss.n23113 vss.n23112 9.3
R14406 vss.n23112 vss.n23111 9.3
R14407 vss.n23111 vss.n23110 9.3
R14408 vss.n23099 vss.n23098 9.3
R14409 vss.n23101 vss.n23100 9.3
R14410 vss.n23085 vss.n23084 9.3
R14411 vss.n23097 vss.n23096 9.3
R14412 vss.n23096 vss.n23095 9.3
R14413 vss.n23095 vss.n23094 9.3
R14414 vss.n23081 vss.n23080 9.3
R14415 vss.n23080 vss.n23079 9.3
R14416 vss.n23079 vss.n23078 9.3
R14417 vss.n23067 vss.n23066 9.3
R14418 vss.n23069 vss.n23068 9.3
R14419 vss.n23049 vss.n23048 9.3
R14420 vss.n23065 vss.n23064 9.3
R14421 vss.n23064 vss.n23063 9.3
R14422 vss.n23063 vss.n23062 9.3
R14423 vss.n23038 vss.n23037 9.3
R14424 vss.n23036 vss.n23035 9.3
R14425 vss.n23035 vss.n23034 9.3
R14426 vss.n23034 vss.n23033 9.3
R14427 vss.n23016 vss.n23015 9.3
R14428 vss.n23015 vss.n23014 9.3
R14429 vss.n23014 vss.n23013 9.3
R14430 vss.n23018 vss.n23017 9.3
R14431 vss.n23002 vss.n23001 9.3
R14432 vss.n23000 vss.n22999 9.3
R14433 vss.n22999 vss.n22998 9.3
R14434 vss.n22998 vss.n22997 9.3
R14435 vss.n22984 vss.n22983 9.3
R14436 vss.n22983 vss.n22982 9.3
R14437 vss.n22982 vss.n22981 9.3
R14438 vss.n22986 vss.n22985 9.3
R14439 vss.n22970 vss.n22969 9.3
R14440 vss.n22968 vss.n22967 9.3
R14441 vss.n22967 vss.n22966 9.3
R14442 vss.n22966 vss.n22965 9.3
R14443 vss.n22952 vss.n22951 9.3
R14444 vss.n22951 vss.n22950 9.3
R14445 vss.n22950 vss.n22949 9.3
R14446 vss.n22954 vss.n22953 9.3
R14447 vss.n22938 vss.n22937 9.3
R14448 vss.n22936 vss.n22935 9.3
R14449 vss.n22935 vss.n22934 9.3
R14450 vss.n22934 vss.n22933 9.3
R14451 vss.n1375 vss.n1374 9.3
R14452 vss.n1374 vss.n1373 9.3
R14453 vss.n1387 vss.n1386 9.3
R14454 vss.n1386 vss.n1385 9.3
R14455 vss.n22917 vss.n22916 9.3
R14456 vss.n22916 vss.n22915 9.3
R14457 vss.n22915 vss.n22914 9.3
R14458 vss.n22904 vss.n22903 9.3
R14459 vss.n22906 vss.n22905 9.3
R14460 vss.n22891 vss.n22890 9.3
R14461 vss.n22902 vss.n22901 9.3
R14462 vss.n22901 vss.n22900 9.3
R14463 vss.n22900 vss.n22899 9.3
R14464 vss.n22887 vss.n22886 9.3
R14465 vss.n22886 vss.n22885 9.3
R14466 vss.n22885 vss.n22884 9.3
R14467 vss.n22874 vss.n22873 9.3
R14468 vss.n22876 vss.n22875 9.3
R14469 vss.n22861 vss.n22860 9.3
R14470 vss.n22872 vss.n22871 9.3
R14471 vss.n22871 vss.n22870 9.3
R14472 vss.n22870 vss.n22869 9.3
R14473 vss.n22857 vss.n22856 9.3
R14474 vss.n22856 vss.n22855 9.3
R14475 vss.n22855 vss.n22854 9.3
R14476 vss.n22844 vss.n22843 9.3
R14477 vss.n22846 vss.n22845 9.3
R14478 vss.n1416 vss.n1415 9.3
R14479 vss.n1414 vss.n1413 9.3
R14480 vss.n1421 vss.n1420 9.3
R14481 vss.n1419 vss.n1418 9.3
R14482 vss.n1424 vss.n1423 9.3
R14483 vss.n22839 vss.n22838 9.3
R14484 vss.n22838 vss.n22837 9.3
R14485 vss.n1406 vss.n1405 9.3
R14486 vss.n1410 vss.n1409 9.3
R14487 vss.n1408 vss.n1407 9.3
R14488 vss.n1463 vss.n1462 9.3
R14489 vss.n1462 vss.n1461 9.3
R14490 vss.n22806 vss.n22805 9.3
R14491 vss.n22842 vss.n1401 9.3
R14492 vss.n1401 vss.n1400 9.3
R14493 vss.n1400 vss.n1399 9.3
R14494 vss.n22823 vss.n22822 9.3
R14495 vss.n22822 vss.n22821 9.3
R14496 vss.n22821 vss.n22820 9.3
R14497 vss.n1440 vss.n1439 9.3
R14498 vss.n1439 vss.n1438 9.3
R14499 vss.n1451 vss.n1450 9.3
R14500 vss.n1450 vss.n1449 9.3
R14501 vss.n22804 vss.n22803 9.3
R14502 vss.n22802 vss.n22801 9.3
R14503 vss.n22801 vss.n22800 9.3
R14504 vss.n22800 vss.n22799 9.3
R14505 vss.n19014 vss.n17635 9.154
R14506 vss.n17635 vss.n17634 9.154
R14507 vss.n18889 vss.n18888 9.154
R14508 vss.n18888 vss.n18887 9.154
R14509 vss.n18767 vss.n17841 9.154
R14510 vss.n17841 vss.n17840 9.154
R14511 vss.n18648 vss.n18647 9.154
R14512 vss.n18647 vss.n18646 9.154
R14513 vss.n18526 vss.n18054 9.154
R14514 vss.n18054 vss.n18053 9.154
R14515 vss.n18407 vss.n18406 9.154
R14516 vss.n18406 vss.n18405 9.154
R14517 vss.n18285 vss.n18267 9.154
R14518 vss.n18267 vss.n18266 9.154
R14519 vss.n20311 vss.n17612 9.154
R14520 vss.n20281 vss.n20280 9.154
R14521 vss.n20282 vss.n20281 9.154
R14522 vss.n20160 vss.n19141 9.154
R14523 vss.n19141 vss.n19140 9.154
R14524 vss.n20035 vss.n20034 9.154
R14525 vss.n20034 vss.n20033 9.154
R14526 vss.n19913 vss.n19348 9.154
R14527 vss.n19348 vss.n19347 9.154
R14528 vss.n19788 vss.n19787 9.154
R14529 vss.n19787 vss.n19786 9.154
R14530 vss.n19666 vss.n19555 9.154
R14531 vss.n19555 vss.n19554 9.154
R14532 vss.n9651 vss.n9650 9.154
R14533 vss.n10216 vss.n10215 9.154
R14534 vss.n9639 vss.n9638 9.154
R14535 vss.n9638 vss.n9637 9.154
R14536 vss.n9645 vss.n9644 9.154
R14537 vss.n9644 vss.n9643 9.154
R14538 vss.n9159 vss.n9158 9.154
R14539 vss.n9158 vss.n9157 9.154
R14540 vss.n9654 vss.n9653 9.154
R14541 vss.n9653 vss.n9652 9.154
R14542 vss.n10219 vss.n10218 9.154
R14543 vss.n10218 vss.n10217 9.154
R14544 vss.n10213 vss.n10212 9.154
R14545 vss.n10212 vss.n10211 9.154
R14546 vss.n10207 vss.n10206 9.154
R14547 vss.n10206 vss.n10205 9.154
R14548 vss.n10201 vss.n10200 9.154
R14549 vss.n10200 vss.n10199 9.154
R14550 vss.n10195 vss.n10194 9.154
R14551 vss.n10194 vss.n10193 9.154
R14552 vss.n10190 vss.n10189 9.154
R14553 vss.n10189 vss.n10188 9.154
R14554 vss.n9702 vss.n9701 9.154
R14555 vss.n9701 vss.n9700 9.154
R14556 vss.n9708 vss.n9707 9.154
R14557 vss.n9707 vss.n9706 9.154
R14558 vss.n9712 vss.n9711 9.154
R14559 vss.n9711 vss.n9710 9.154
R14560 vss.n9699 vss.n9698 9.154
R14561 vss.n9698 vss.n9697 9.154
R14562 vss.n9719 vss.n9718 9.154
R14563 vss.n9718 vss.n9717 9.154
R14564 vss.n9725 vss.n9724 9.154
R14565 vss.n9724 vss.n9723 9.154
R14566 vss.n9731 vss.n9730 9.154
R14567 vss.n9730 vss.n9729 9.154
R14568 vss.n9737 vss.n9736 9.154
R14569 vss.n9736 vss.n9735 9.154
R14570 vss.n9743 vss.n9742 9.154
R14571 vss.n9742 vss.n9741 9.154
R14572 vss.n10182 vss.n10181 9.154
R14573 vss.n10181 vss.n10180 9.154
R14574 vss.n13307 vss.n13306 9.154
R14575 vss.n12574 vss.n12572 9.154
R14576 vss.n11168 vss.n11167 9.154
R14577 vss.n14409 vss.n14408 9.154
R14578 vss.n5624 vss.n4245 9.154
R14579 vss.n4245 vss.n4244 9.154
R14580 vss.n5499 vss.n5498 9.154
R14581 vss.n5498 vss.n5497 9.154
R14582 vss.n5377 vss.n4451 9.154
R14583 vss.n4451 vss.n4450 9.154
R14584 vss.n5258 vss.n5257 9.154
R14585 vss.n5257 vss.n5256 9.154
R14586 vss.n5136 vss.n4664 9.154
R14587 vss.n4664 vss.n4663 9.154
R14588 vss.n5017 vss.n5016 9.154
R14589 vss.n5016 vss.n5015 9.154
R14590 vss.n4895 vss.n4877 9.154
R14591 vss.n4877 vss.n4876 9.154
R14592 vss.n6921 vss.n4222 9.154
R14593 vss.n6891 vss.n6890 9.154
R14594 vss.n6892 vss.n6891 9.154
R14595 vss.n6770 vss.n5751 9.154
R14596 vss.n5751 vss.n5750 9.154
R14597 vss.n6645 vss.n6644 9.154
R14598 vss.n6644 vss.n6643 9.154
R14599 vss.n6523 vss.n5958 9.154
R14600 vss.n5958 vss.n5957 9.154
R14601 vss.n6398 vss.n6397 9.154
R14602 vss.n6397 vss.n6396 9.154
R14603 vss.n6276 vss.n6165 9.154
R14604 vss.n6165 vss.n6164 9.154
R14605 vss.n15421 vss.n15420 9.154
R14606 vss.n15420 vss.n15419 9.154
R14607 vss.n15657 vss.n15656 9.154
R14608 vss.n15656 vss.n15655 9.154
R14609 vss.n16301 vss.n16300 9.154
R14610 vss.n16300 vss.n16299 9.154
R14611 vss.n16368 vss.n16367 9.154
R14612 vss.n16367 vss.n16366 9.154
R14613 vss.n16604 vss.n16603 9.154
R14614 vss.n16603 vss.n16602 9.154
R14615 vss.n16697 vss.n16694 9.154
R14616 vss.n16694 vss.n16693 9.154
R14617 vss.n16711 vss.n16708 9.154
R14618 vss.n16708 vss.n16707 9.154
R14619 vss.n16725 vss.n16722 9.154
R14620 vss.n16722 vss.n16721 9.154
R14621 vss.n16739 vss.n16736 9.154
R14622 vss.n16736 vss.n16735 9.154
R14623 vss.n16753 vss.n16750 9.154
R14624 vss.n16750 vss.n16749 9.154
R14625 vss.n16683 vss.n16682 9.154
R14626 vss.n16682 vss.n16681 9.154
R14627 vss.n16765 vss.n16764 9.154
R14628 vss.n16764 vss.n16763 9.154
R14629 vss.n16777 vss.n16776 9.154
R14630 vss.n16776 vss.n16775 9.154
R14631 vss.n16795 vss.n16794 9.154
R14632 vss.n16794 vss.n16793 9.154
R14633 vss.n16806 vss.n16805 9.154
R14634 vss.n16805 vss.n16804 9.154
R14635 vss.n16820 vss.n16819 9.154
R14636 vss.n16819 vss.n16818 9.154
R14637 vss.n16834 vss.n16833 9.154
R14638 vss.n16833 vss.n16832 9.154
R14639 vss.n16848 vss.n16847 9.154
R14640 vss.n16847 vss.n16846 9.154
R14641 vss.n16876 vss.n16873 9.154
R14642 vss.n16873 vss.n16872 9.154
R14643 vss.n16890 vss.n16887 9.154
R14644 vss.n16887 vss.n16886 9.154
R14645 vss.n16913 vss.n16910 9.154
R14646 vss.n16910 vss.n16909 9.154
R14647 vss.n16927 vss.n16924 9.154
R14648 vss.n16924 vss.n16923 9.154
R14649 vss.n16941 vss.n16938 9.154
R14650 vss.n16938 vss.n16937 9.154
R14651 vss.n16955 vss.n16952 9.154
R14652 vss.n16952 vss.n16951 9.154
R14653 vss.n16969 vss.n16966 9.154
R14654 vss.n16966 vss.n16965 9.154
R14655 vss.n16983 vss.n16980 9.154
R14656 vss.n16980 vss.n16979 9.154
R14657 vss.n16997 vss.n16994 9.154
R14658 vss.n16994 vss.n16993 9.154
R14659 vss.n17011 vss.n17008 9.154
R14660 vss.n17008 vss.n17007 9.154
R14661 vss.n16862 vss.n16859 9.154
R14662 vss.n16859 vss.n16858 9.154
R14663 vss.n17264 vss.n17263 9.154
R14664 vss.n17263 vss.n17262 9.154
R14665 vss.n17028 vss.n17025 9.154
R14666 vss.n17025 vss.n17024 9.154
R14667 vss.n17042 vss.n17039 9.154
R14668 vss.n17039 vss.n17038 9.154
R14669 vss.n17056 vss.n17053 9.154
R14670 vss.n17053 vss.n17052 9.154
R14671 vss.n17070 vss.n17067 9.154
R14672 vss.n17067 vss.n17066 9.154
R14673 vss.n17084 vss.n17081 9.154
R14674 vss.n17081 vss.n17080 9.154
R14675 vss.n17098 vss.n17095 9.154
R14676 vss.n17095 vss.n17094 9.154
R14677 vss.n17112 vss.n17109 9.154
R14678 vss.n17109 vss.n17108 9.154
R14679 vss.n17126 vss.n17123 9.154
R14680 vss.n17123 vss.n17122 9.154
R14681 vss.n17149 vss.n17146 9.154
R14682 vss.n17146 vss.n17145 9.154
R14683 vss.n17163 vss.n17160 9.154
R14684 vss.n17160 vss.n17159 9.154
R14685 vss.n17177 vss.n17174 9.154
R14686 vss.n17174 vss.n17173 9.154
R14687 vss.n17191 vss.n17188 9.154
R14688 vss.n17188 vss.n17187 9.154
R14689 vss.n17205 vss.n17202 9.154
R14690 vss.n17202 vss.n17201 9.154
R14691 vss.n17219 vss.n17216 9.154
R14692 vss.n17216 vss.n17215 9.154
R14693 vss.n17233 vss.n17230 9.154
R14694 vss.n17230 vss.n17229 9.154
R14695 vss.n17247 vss.n17244 9.154
R14696 vss.n17244 vss.n17243 9.154
R14697 vss.n16264 vss.n16263 9.154
R14698 vss.n16263 vss.n16262 9.154
R14699 vss.n17274 vss.n17271 9.154
R14700 vss.n17271 vss.n17270 9.154
R14701 vss.n17284 vss.n17283 9.154
R14702 vss.n17283 vss.n17282 9.154
R14703 vss.n17295 vss.n17294 9.154
R14704 vss.n17294 vss.n17293 9.154
R14705 vss.n17305 vss.n17304 9.154
R14706 vss.n17304 vss.n17303 9.154
R14707 vss.n17326 vss.n17323 9.154
R14708 vss.n17323 vss.n17322 9.154
R14709 vss.n17315 vss.n17312 9.154
R14710 vss.n17312 vss.n17311 9.154
R14711 vss.n12566 vss.n12564 9.095
R14712 vss.n14389 vss.n14388 9.095
R14713 vss.n13287 vss.n13286 9.095
R14714 vss.n9028 vss.n9027 9.086
R14715 vss.n15880 vss.n15879 9.013
R14716 vss.n15879 vss.n15878 9.013
R14717 vss.n15945 vss.n15944 9.013
R14718 vss.n15944 vss.n15943 9.013
R14719 vss.n16181 vss.n16180 9.013
R14720 vss.n16180 vss.n16179 9.013
R14721 vss.n16901 vss.n16899 9.013
R14722 vss.n16899 vss.n16898 9.013
R14723 vss.n17137 vss.n17135 9.013
R14724 vss.n17135 vss.n17134 9.013
R14725 vss.n20331 vss.n17575 8.918
R14726 vss.n6941 vss.n4185 8.918
R14727 vss.n11166 vss.n11165 8.897
R14728 vss.n3454 vss.n3453 8.87
R14729 vss.n1429 vss.n1428 8.87
R14730 vss.n11538 vss.n11537 8.855
R14731 vss.n12378 vss.n12377 8.855
R14732 vss.n13180 vss.n13179 8.855
R14733 vss.n12939 vss.n12938 8.855
R14734 vss.n11965 vss.n11964 8.855
R14735 vss.n12094 vss.n12092 8.855
R14736 vss.n10994 vss.n10993 8.855
R14737 vss.n10719 vss.n10718 8.855
R14738 vss.n13009 vss.n13008 8.855
R14739 vss.n10557 vss.n10556 8.855
R14740 vss.n12970 vss.n12969 8.855
R14741 vss.n12342 vss.n12341 8.855
R14742 vss.n13766 vss.n13765 8.855
R14743 vss.n13806 vss.n13805 8.855
R14744 vss.n11502 vss.n11501 8.855
R14745 vss.n14763 vss.n14762 8.855
R14746 vss.n13553 vss.n13552 8.855
R14747 vss.n14438 vss.n14437 8.855
R14748 vss.n21796 vss.n21661 8.804
R14749 vss.n3745 vss.n3610 8.804
R14750 vss.n21796 vss.n21649 8.737
R14751 vss.n3745 vss.n3598 8.737
R14752 vss.n20303 vss.n17610 8.57
R14753 vss.n6913 vss.n4220 8.57
R14754 vss.n11529 vss.n11528 8.57
R14755 vss.n12368 vss.n12367 8.57
R14756 vss.n13169 vss.n13168 8.57
R14757 vss.n12927 vss.n12926 8.57
R14758 vss.n10710 vss.n10709 8.57
R14759 vss.n12999 vss.n12998 8.57
R14760 vss.n10563 vss.n10562 8.57
R14761 vss.n12348 vss.n12347 8.57
R14762 vss.n11508 vss.n11507 8.57
R14763 vss.n9059 vss.n9058 8.568
R14764 vss.n1746 vss.n1745 8.541
R14765 vss.n207 vss.n206 8.541
R14766 vss.n20317 vss.n17608 8.533
R14767 vss.n6927 vss.n4218 8.533
R14768 vss.n17544 vss.n17543 8.5
R14769 vss.n17499 vss.n17498 8.5
R14770 vss.n4154 vss.n4153 8.5
R14771 vss.n4109 vss.n4108 8.5
R14772 vss.n3448 vss.n3447 8.5
R14773 vss.n1423 vss.n1422 8.5
R14774 vss.n14178 vss.n14177 8.45
R14775 vss.n10869 vss.n10868 8.45
R14776 vss.n13811 vss.n13810 8.45
R14777 vss.n12286 vss.n12285 8.45
R14778 vss.n10766 vss.n10765 8.45
R14779 vss.n13485 vss.n13484 8.45
R14780 vss.n13394 vss.n13393 8.45
R14781 vss.n13170 vss.n13169 8.45
R14782 vss.n12929 vss.n12927 8.45
R14783 vss.n12101 vss.n12099 8.45
R14784 vss.n11236 vss.n11234 8.45
R14785 vss.n10711 vss.n10710 8.45
R14786 vss.n10565 vss.n10563 8.45
R14787 vss.n11342 vss.n11341 8.45
R14788 vss.n13723 vss.n13722 8.45
R14789 vss.n14148 vss.n14147 8.45
R14790 vss.n13604 vss.n13603 8.45
R14791 vss.n11335 vss.n11334 8.45
R14792 vss.n13001 vss.n12999 8.45
R14793 vss.n12960 vss.n12958 8.45
R14794 vss.n13062 vss.n13061 8.45
R14795 vss.n13051 vss.n13050 8.45
R14796 vss.n12370 vss.n12368 8.45
R14797 vss.n12350 vss.n12348 8.45
R14798 vss.n12445 vss.n12444 8.45
R14799 vss.n13774 vss.n13772 8.45
R14800 vss.n13716 vss.n13715 8.45
R14801 vss.n11510 vss.n11508 8.45
R14802 vss.n11530 vss.n11529 8.45
R14803 vss.n14023 vss.n14022 8.45
R14804 vss.n14287 vss.n14286 8.45
R14805 vss.n11710 vss.n11709 8.45
R14806 vss.n13282 vss.n13281 8.45
R14807 vss.n13523 vss.n13522 8.45
R14808 vss.n12786 vss.n12785 8.45
R14809 vss.n13209 vss.n13208 8.45
R14810 vss.n20317 vss.n17609 8.228
R14811 vss.n20306 vss.n17610 8.228
R14812 vss.n6927 vss.n4219 8.228
R14813 vss.n6916 vss.n4220 8.228
R14814 vss.n21789 vss.n21692 8.139
R14815 vss.n3738 vss.n3641 8.139
R14816 vss.n10257 vss.n10256 8.116
R14817 vss.n21789 vss.n21788 8.111
R14818 vss.n3738 vss.n3737 8.111
R14819 vss.n14135 vss.n14134 8.11
R14820 vss.n12275 vss.n12274 8.11
R14821 vss.n10465 vss.n10464 8.11
R14822 vss.n10606 vss.n10605 8.11
R14823 vss.n21790 vss.n21789 8.083
R14824 vss.n3739 vss.n3738 8.083
R14825 vss.n21789 vss.n21695 8.056
R14826 vss.n3738 vss.n3644 8.056
R14827 vss.n21789 vss.n21693 8.029
R14828 vss.n3738 vss.n3642 8.029
R14829 vss.n21789 vss.n21787 8.003
R14830 vss.n3738 vss.n3736 8.003
R14831 vss.n19028 vss.n17626 7.88
R14832 vss.n19000 vss.n17643 7.88
R14833 vss.n18897 vss.n17722 7.88
R14834 vss.n18876 vss.n17745 7.88
R14835 vss.n18780 vss.n17828 7.88
R14836 vss.n18759 vss.n17852 7.88
R14837 vss.n18656 vss.n17935 7.88
R14838 vss.n18635 vss.n17958 7.88
R14839 vss.n18539 vss.n18041 7.88
R14840 vss.n18518 vss.n18065 7.88
R14841 vss.n18415 vss.n18148 7.88
R14842 vss.n18394 vss.n18171 7.88
R14843 vss.n18298 vss.n18254 7.88
R14844 vss.n20269 vss.n19041 7.88
R14845 vss.n20173 vss.n19128 7.88
R14846 vss.n20146 vss.n19150 7.88
R14847 vss.n20043 vss.n19229 7.88
R14848 vss.n20022 vss.n19252 7.88
R14849 vss.n19926 vss.n19335 7.88
R14850 vss.n19899 vss.n19357 7.88
R14851 vss.n19796 vss.n19436 7.88
R14852 vss.n19775 vss.n19459 7.88
R14853 vss.n19679 vss.n19542 7.88
R14854 vss.n19652 vss.n19564 7.88
R14855 vss.n20320 vss.n17605 7.88
R14856 vss.n20297 vss.n20295 7.88
R14857 vss.n5638 vss.n4236 7.88
R14858 vss.n5610 vss.n4253 7.88
R14859 vss.n5507 vss.n4332 7.88
R14860 vss.n5486 vss.n4355 7.88
R14861 vss.n5390 vss.n4438 7.88
R14862 vss.n5369 vss.n4462 7.88
R14863 vss.n5266 vss.n4545 7.88
R14864 vss.n5245 vss.n4568 7.88
R14865 vss.n5149 vss.n4651 7.88
R14866 vss.n5128 vss.n4675 7.88
R14867 vss.n5025 vss.n4758 7.88
R14868 vss.n5004 vss.n4781 7.88
R14869 vss.n4908 vss.n4864 7.88
R14870 vss.n6879 vss.n5651 7.88
R14871 vss.n6783 vss.n5738 7.88
R14872 vss.n6756 vss.n5760 7.88
R14873 vss.n6653 vss.n5839 7.88
R14874 vss.n6632 vss.n5862 7.88
R14875 vss.n6536 vss.n5945 7.88
R14876 vss.n6509 vss.n5967 7.88
R14877 vss.n6406 vss.n6046 7.88
R14878 vss.n6385 vss.n6069 7.88
R14879 vss.n6289 vss.n6152 7.88
R14880 vss.n6262 vss.n6174 7.88
R14881 vss.n6930 vss.n4215 7.88
R14882 vss.n6907 vss.n6905 7.88
R14883 vss.n16694 vss.n16690 7.88
R14884 vss.n16873 vss.n16869 7.88
R14885 vss.n16924 vss.n16920 7.88
R14886 vss.n17109 vss.n17105 7.88
R14887 vss.n17160 vss.n17156 7.88
R14888 vss.n17271 vss.n17267 7.88
R14889 vss.n15879 vss.n15876 7.88
R14890 vss.n15919 vss.n15915 7.88
R14891 vss.n15971 vss.n15967 7.88
R14892 vss.n16155 vss.n16151 7.88
R14893 vss.n16207 vss.n16203 7.88
R14894 vss.n16280 vss.n16276 7.88
R14895 vss.n15395 vss.n15391 7.88
R14896 vss.n15444 vss.n15440 7.88
R14897 vss.n15631 vss.n15627 7.88
R14898 vss.n15680 vss.n15676 7.88
R14899 vss.n15859 vss.n15855 7.88
R14900 vss.n16300 vss.n16297 7.88
R14901 vss.n16342 vss.n16338 7.88
R14902 vss.n16391 vss.n16387 7.88
R14903 vss.n16578 vss.n16574 7.88
R14904 vss.n16627 vss.n16623 7.88
R14905 vss.n10259 vss.n10258 7.863
R14906 vss.n12427 vss.n12423 7.801
R14907 vss.n12600 vss.n12596 7.801
R14908 vss.n14493 vss.n14489 7.801
R14909 vss.n14400 vss.n14396 7.801
R14910 vss.n14663 vss.n14659 7.801
R14911 vss.n13582 vss.n13578 7.801
R14912 vss.n15017 vss.n15013 7.801
R14913 vss.n10508 vss.n10504 7.801
R14914 vss.n13300 vss.n13296 7.801
R14915 vss.n13341 vss.n13337 7.801
R14916 vss.n13242 vss.n13238 7.801
R14917 vss.n14963 vss.n14959 7.801
R14918 vss.n14359 vss.n14355 7.801
R14919 vss.n13865 vss.n13861 7.801
R14920 vss.n13980 vss.n13976 7.801
R14921 vss.n11575 vss.n11571 7.801
R14922 vss.n11762 vss.n11758 7.801
R14923 vss.n11052 vss.n11048 7.801
R14924 vss.n10826 vss.n10822 7.801
R14925 vss.n10900 vss.n10896 7.801
R14926 vss.n10953 vss.n10949 7.801
R14927 vss.n11013 vss.n11009 7.801
R14928 vss.n12585 vss.n12581 7.801
R14929 vss.n12081 vss.n12077 7.801
R14930 vss.n17604 vss.n17575 7.787
R14931 vss.n4214 vss.n4185 7.787
R14932 vss.n20307 vss.n20306 7.771
R14933 vss.n6917 vss.n6916 7.771
R14934 vss.n22718 vss.n22715 7.725
R14935 vss.n22669 vss.n22666 7.725
R14936 vss.n22510 vss.n22507 7.725
R14937 vss.n22461 vss.n22458 7.725
R14938 vss.n22302 vss.n22299 7.725
R14939 vss.n22253 vss.n22250 7.725
R14940 vss.n22094 vss.n22091 7.725
R14941 vss.n21585 vss.n21582 7.725
R14942 vss.n21438 vss.n21435 7.725
R14943 vss.n21389 vss.n21386 7.725
R14944 vss.n21230 vss.n21227 7.725
R14945 vss.n21181 vss.n21178 7.725
R14946 vss.n21022 vss.n21019 7.725
R14947 vss.n20973 vss.n20970 7.725
R14948 vss.n8881 vss.n8878 7.725
R14949 vss.n8832 vss.n8829 7.725
R14950 vss.n8673 vss.n8670 7.725
R14951 vss.n8624 vss.n8621 7.725
R14952 vss.n8465 vss.n8462 7.725
R14953 vss.n8416 vss.n8413 7.725
R14954 vss.n8257 vss.n8254 7.725
R14955 vss.n8208 vss.n8205 7.725
R14956 vss.n8049 vss.n8046 7.725
R14957 vss.n8000 vss.n7997 7.725
R14958 vss.n7840 vss.n7837 7.725
R14959 vss.n7791 vss.n7788 7.725
R14960 vss.n7632 vss.n7629 7.725
R14961 vss.n7583 vss.n7580 7.725
R14962 vss.n13709 vss.n13708 7.645
R14963 vss.n13032 vss.n13031 7.645
R14964 vss.n14348 vss.n14347 7.645
R14965 vss.n14481 vss.n14480 7.645
R14966 vss.n10757 vss.n10756 7.645
R14967 vss.n12794 vss.n12793 7.645
R14968 vss.n13043 vss.n13042 7.645
R14969 vss.n13696 vss.n13695 7.645
R14970 vss.n17610 vss.n17608 7.585
R14971 vss.n4220 vss.n4218 7.585
R14972 vss.n12571 vss.n12570 7.583
R14973 vss.n11166 vss.n11164 7.582
R14974 vss.n21925 vss.n21924 7.512
R14975 vss.n21952 vss.n21951 7.512
R14976 vss.n3874 vss.n3873 7.512
R14977 vss.n3901 vss.n3900 7.512
R14978 vss.n9005 vss.n9004 7.356
R14979 vss.n17610 vss.n17609 7.314
R14980 vss.n4220 vss.n4219 7.314
R14981 vss.n11350 vss.n11347 7.272
R14982 vss.n10759 vss.n10758 7.272
R14983 vss.n13045 vss.n13044 7.272
R14984 vss.n12796 vss.n12795 7.272
R14985 vss.n13710 vss.n13706 7.271
R14986 vss.n10747 vss.n10744 7.271
R14987 vss.n9090 vss.n9089 7.267
R14988 vss.n10460 vss.n10459 7.248
R14989 vss.n10868 vss.n10866 7.231
R14990 vss.n12927 vss.n12924 7.231
R14991 vss.n10589 vss.n10588 7.231
R14992 vss.n10496 vss.n10495 7.231
R14993 vss.n11394 vss.n11393 7.231
R14994 vss.n13622 vss.n13621 7.229
R14995 vss.n13134 vss.n13133 7.224
R14996 vss.n13674 vss.n13673 7.224
R14997 vss.n13124 vss.n13123 7.224
R14998 vss.n13125 vss.n13124 7.224
R14999 vss.n13643 vss.n13642 7.224
R15000 vss.n11467 vss.n11466 7.224
R15001 vss.n11466 vss.n11465 7.224
R15002 vss.n10661 vss.n10660 7.224
R15003 vss.n10654 vss.n10653 7.224
R15004 vss.n11458 vss.n11457 7.224
R15005 vss.n13675 vss.n13674 7.224
R15006 vss.n13133 vss.n13132 7.224
R15007 vss.n10662 vss.n10661 7.224
R15008 vss.n11459 vss.n11458 7.224
R15009 vss.n10653 vss.n10652 7.224
R15010 vss.n13642 vss.n13641 7.224
R15011 vss.n11964 vss.n11963 7.189
R15012 vss.n13923 vss.n13922 7.175
R15013 vss.n11269 vss.n11268 7.175
R15014 vss.n13425 vss.n13424 7.175
R15015 vss.n13610 vss.n13609 7.175
R15016 vss.n11022 vss.n11021 7.175
R15017 vss.n12235 vss.n12234 7.175
R15018 vss.n12516 vss.n12515 7.175
R15019 vss.n13196 vss.n13195 7.175
R15020 vss.n13434 vss.n13433 7.175
R15021 vss.n13620 vss.n13619 7.175
R15022 vss.n11392 vss.n11391 7.175
R15023 vss.n11649 vss.n11648 7.175
R15024 vss.n20314 vss.n17610 7.152
R15025 vss.n20304 vss.n17610 7.152
R15026 vss.n6924 vss.n4220 7.152
R15027 vss.n6914 vss.n4220 7.152
R15028 vss.n13060 vss.t176 7.049
R15029 vss.n12784 vss.t147 7.049
R15030 vss.n13207 vss.t168 7.049
R15031 vss.n9035 vss.n9034 6.977
R15032 vss.n20530 vss.t153 6.94
R15033 vss.n17525 vss.n17524 6.94
R15034 vss.n17512 vss.n17511 6.94
R15035 vss.n20775 vss.t131 6.94
R15036 vss.n7140 vss.t92 6.94
R15037 vss.n4135 vss.n4134 6.94
R15038 vss.n4122 vss.n4121 6.94
R15039 vss.n7385 vss.t126 6.94
R15040 vss.n1647 vss.n1646 6.94
R15041 vss.n1635 vss.n1634 6.94
R15042 vss.n1620 vss.n1619 6.94
R15043 vss.n1608 vss.n1607 6.94
R15044 vss.n1595 vss.n1594 6.94
R15045 vss.n1583 vss.n1582 6.94
R15046 vss.n2476 vss.t51 6.94
R15047 vss.n1570 vss.n1569 6.94
R15048 vss.n1557 vss.n1556 6.94
R15049 vss.n2743 vss.t71 6.94
R15050 vss.n1540 vss.n1539 6.94
R15051 vss.n1525 vss.n1524 6.94
R15052 vss.n1512 vss.n1511 6.94
R15053 vss.n1500 vss.n1499 6.94
R15054 vss.n1485 vss.n1484 6.94
R15055 vss.n1473 vss.n1472 6.94
R15056 vss.n108 vss.n107 6.94
R15057 vss.n96 vss.n95 6.94
R15058 vss.n81 vss.n80 6.94
R15059 vss.n69 vss.n68 6.94
R15060 vss.n56 vss.n55 6.94
R15061 vss.n44 vss.n43 6.94
R15062 vss.n937 vss.t295 6.94
R15063 vss.n31 vss.n30 6.94
R15064 vss.n18 vss.n17 6.94
R15065 vss.n1204 vss.t251 6.94
R15066 vss.n1320 vss.n1319 6.94
R15067 vss.n1332 vss.n1331 6.94
R15068 vss.n1346 vss.n1345 6.94
R15069 vss.n1358 vss.n1357 6.94
R15070 vss.n1373 vss.n1372 6.94
R15071 vss.n1385 vss.n1384 6.94
R15072 vss.n13552 vss.n13551 6.922
R15073 vss.n12341 vss.n12340 6.883
R15074 vss.n13765 vss.n13764 6.883
R15075 vss.n10993 vss.n10992 6.883
R15076 vss.n12092 vss.n12091 6.883
R15077 vss.n20336 vss.n17600 6.815
R15078 vss.n20333 vss.n17600 6.815
R15079 vss.n6946 vss.n4210 6.815
R15080 vss.n6943 vss.n4210 6.815
R15081 vss.n14177 vss.n14175 6.674
R15082 vss.n2915 vss.n2913 6.64
R15083 vss.n23343 vss.n1336 6.64
R15084 vss.n1879 vss.n1626 6.639
R15085 vss.n3111 vss.n1491 6.639
R15086 vss.n3333 vss.n1489 6.639
R15087 vss.n340 vss.n87 6.639
R15088 vss.n23146 vss.n1362 6.639
R15089 vss.n22924 vss.n1364 6.639
R15090 vss.n2400 vss.n2398 6.638
R15091 vss.n3216 vss.n1490 6.638
R15092 vss.n861 vss.n859 6.638
R15093 vss.n23041 vss.n1363 6.638
R15094 vss.n12958 vss.n12956 6.638
R15095 vss.n11234 vss.n11232 6.638
R15096 vss.n1996 vss.n1625 6.638
R15097 vss.n2101 vss.n1624 6.638
R15098 vss.n2188 vss.n1599 6.638
R15099 vss.n2299 vss.n2297 6.638
R15100 vss.n2509 vss.n1574 6.638
R15101 vss.n2609 vss.n1561 6.638
R15102 vss.n2709 vss.n1548 6.638
R15103 vss.n3012 vss.n1516 6.638
R15104 vss.n457 vss.n86 6.638
R15105 vss.n562 vss.n85 6.638
R15106 vss.n649 vss.n60 6.638
R15107 vss.n760 vss.n758 6.638
R15108 vss.n970 vss.n35 6.638
R15109 vss.n1070 vss.n22 6.638
R15110 vss.n1170 vss.n9 6.638
R15111 vss.n23245 vss.n1337 6.638
R15112 vss.n2819 vss.n1547 6.636
R15113 vss.n1281 vss.n8 6.636
R15114 vss.n20547 vss.n17530 6.606
R15115 vss.n7157 vss.n4140 6.606
R15116 vss.n21619 vss.n21617 6.605
R15117 vss.n3568 vss.n3566 6.605
R15118 vss.n21863 vss.n21862 6.604
R15119 vss.n3812 vss.n3811 6.604
R15120 vss.n20749 vss.n17504 6.601
R15121 vss.n7359 vss.n4114 6.601
R15122 vss.n20655 vss.n17516 6.601
R15123 vss.n7265 vss.n4126 6.601
R15124 vss.n20524 vss.n20523 6.586
R15125 vss.n20552 vss.n20551 6.586
R15126 vss.n20753 vss.n20752 6.586
R15127 vss.n20774 vss.n20773 6.586
R15128 vss.n7134 vss.n7133 6.586
R15129 vss.n7162 vss.n7161 6.586
R15130 vss.n7363 vss.n7362 6.586
R15131 vss.n7384 vss.n7383 6.586
R15132 vss.n1750 vss.n1749 6.586
R15133 vss.n1771 vss.n1770 6.586
R15134 vss.n1979 vss.n1978 6.586
R15135 vss.n2009 vss.n2008 6.586
R15136 vss.n2224 vss.n2223 6.586
R15137 vss.n2253 vss.n2252 6.586
R15138 vss.n2468 vss.n2467 6.586
R15139 vss.n2497 vss.n2496 6.586
R15140 vss.n2713 vss.n2712 6.586
R15141 vss.n2742 vss.n2741 6.586
R15142 vss.n2951 vss.n2950 6.586
R15143 vss.n2980 vss.n2979 6.586
R15144 vss.n3195 vss.n3194 6.586
R15145 vss.n3225 vss.n3224 6.586
R15146 vss.n15199 vss.n15198 6.586
R15147 vss.n15180 vss.n15179 6.586
R15148 vss.n211 vss.n210 6.586
R15149 vss.n232 vss.n231 6.586
R15150 vss.n440 vss.n439 6.586
R15151 vss.n470 vss.n469 6.586
R15152 vss.n685 vss.n684 6.586
R15153 vss.n714 vss.n713 6.586
R15154 vss.n929 vss.n928 6.586
R15155 vss.n958 vss.n957 6.586
R15156 vss.n1174 vss.n1173 6.586
R15157 vss.n1203 vss.n1202 6.586
R15158 vss.n23297 vss.n23296 6.586
R15159 vss.n23270 vss.n23269 6.586
R15160 vss.n23053 vss.n23052 6.586
R15161 vss.n23025 vss.n23024 6.586
R15162 vss.n1392 vss.n1391 6.586
R15163 vss.n22814 vss.n22813 6.586
R15164 vss.n1797 vss.n1786 6.477
R15165 vss.n258 vss.n247 6.477
R15166 vss.n20317 vss.n20316 6.344
R15167 vss.n6927 vss.n6926 6.344
R15168 vss.n20658 vss.n17515 6.208
R15169 vss.n7268 vss.n4125 6.208
R15170 vss.n12485 vss.n12469 6.143
R15171 vss.n9114 vss.n9113 6.119
R15172 vss.n17518 vss.n17517 6.023
R15173 vss.n17506 vss.n17505 6.023
R15174 vss.n21830 vss.n21829 6.023
R15175 vss.n21837 vss.n21836 6.023
R15176 vss.n21721 vss.n21720 6.023
R15177 vss.n21729 vss.n21718 6.023
R15178 vss.n21730 vss.n21716 6.023
R15179 vss.n21737 vss.n21736 6.023
R15180 vss.n21764 vss.n21763 6.023
R15181 vss.n21771 vss.n21761 6.023
R15182 vss.n21682 vss.n21664 6.023
R15183 vss.n21677 vss.n21676 6.023
R15184 vss.n12048 vss.n12047 6.023
R15185 vss.n12038 vss.n12037 6.023
R15186 vss.n10967 vss.n10966 6.023
R15187 vss.n10977 vss.n10976 6.023
R15188 vss.n13830 vss.n13829 6.023
R15189 vss.n13820 vss.n13819 6.023
R15190 vss.n11122 vss.n11121 6.023
R15191 vss.n11112 vss.n11111 6.023
R15192 vss.n13361 vss.n13360 6.023
R15193 vss.n13381 vss.n13380 6.023
R15194 vss.n14193 vss.n14192 6.023
R15195 vss.n14203 vss.n14202 6.023
R15196 vss.n12880 vss.n12879 6.023
R15197 vss.n12471 vss.n12470 6.023
R15198 vss.n3779 vss.n3778 6.023
R15199 vss.n3786 vss.n3785 6.023
R15200 vss.n3670 vss.n3669 6.023
R15201 vss.n3678 vss.n3667 6.023
R15202 vss.n3679 vss.n3665 6.023
R15203 vss.n3686 vss.n3685 6.023
R15204 vss.n3713 vss.n3712 6.023
R15205 vss.n3720 vss.n3710 6.023
R15206 vss.n3631 vss.n3613 6.023
R15207 vss.n3626 vss.n3625 6.023
R15208 vss.n4128 vss.n4127 6.023
R15209 vss.n4116 vss.n4115 6.023
R15210 vss.n1640 vss.n1639 6.023
R15211 vss.n1628 vss.n1627 6.023
R15212 vss.n1613 vss.n1612 6.023
R15213 vss.n1601 vss.n1600 6.023
R15214 vss.n1588 vss.n1587 6.023
R15215 vss.n1576 vss.n1575 6.023
R15216 vss.n1563 vss.n1562 6.023
R15217 vss.n1550 vss.n1549 6.023
R15218 vss.n1530 vss.n1529 6.023
R15219 vss.n1518 vss.n1517 6.023
R15220 vss.n1505 vss.n1504 6.023
R15221 vss.n1493 vss.n1492 6.023
R15222 vss.n1478 vss.n1477 6.023
R15223 vss.n1466 vss.n1465 6.023
R15224 vss.n101 vss.n100 6.023
R15225 vss.n89 vss.n88 6.023
R15226 vss.n74 vss.n73 6.023
R15227 vss.n62 vss.n61 6.023
R15228 vss.n49 vss.n48 6.023
R15229 vss.n37 vss.n36 6.023
R15230 vss.n24 vss.n23 6.023
R15231 vss.n11 vss.n10 6.023
R15232 vss.n1313 vss.n1312 6.023
R15233 vss.n1325 vss.n1324 6.023
R15234 vss.n1339 vss.n1338 6.023
R15235 vss.n1351 vss.n1350 6.023
R15236 vss.n1366 vss.n1365 6.023
R15237 vss.n1378 vss.n1377 6.023
R15238 vss.n18965 vss.n17671 5.91
R15239 vss.n17699 vss.n17696 5.91
R15240 vss.n18841 vss.n17778 5.91
R15241 vss.n18815 vss.n17800 5.91
R15242 vss.n17886 vss.n17880 5.91
R15243 vss.n17912 vss.n17909 5.91
R15244 vss.n18600 vss.n17991 5.91
R15245 vss.n18574 vss.n18013 5.91
R15246 vss.n18099 vss.n18093 5.91
R15247 vss.n18125 vss.n18122 5.91
R15248 vss.n18359 vss.n18204 5.91
R15249 vss.n18333 vss.n18226 5.91
R15250 vss.n20234 vss.n19078 5.91
R15251 vss.n20208 vss.n19100 5.91
R15252 vss.n20111 vss.n19178 5.91
R15253 vss.n19206 vss.n19203 5.91
R15254 vss.n19987 vss.n19285 5.91
R15255 vss.n19961 vss.n19307 5.91
R15256 vss.n19864 vss.n19385 5.91
R15257 vss.n19413 vss.n19410 5.91
R15258 vss.n19740 vss.n19492 5.91
R15259 vss.n19714 vss.n19514 5.91
R15260 vss.n19606 vss.n19603 5.91
R15261 vss.n5575 vss.n4281 5.91
R15262 vss.n4309 vss.n4306 5.91
R15263 vss.n5451 vss.n4388 5.91
R15264 vss.n5425 vss.n4410 5.91
R15265 vss.n4496 vss.n4490 5.91
R15266 vss.n4522 vss.n4519 5.91
R15267 vss.n5210 vss.n4601 5.91
R15268 vss.n5184 vss.n4623 5.91
R15269 vss.n4709 vss.n4703 5.91
R15270 vss.n4735 vss.n4732 5.91
R15271 vss.n4969 vss.n4814 5.91
R15272 vss.n4943 vss.n4836 5.91
R15273 vss.n6844 vss.n5688 5.91
R15274 vss.n6818 vss.n5710 5.91
R15275 vss.n6721 vss.n5788 5.91
R15276 vss.n5816 vss.n5813 5.91
R15277 vss.n6597 vss.n5895 5.91
R15278 vss.n6571 vss.n5917 5.91
R15279 vss.n6474 vss.n5995 5.91
R15280 vss.n6023 vss.n6020 5.91
R15281 vss.n6350 vss.n6102 5.91
R15282 vss.n6324 vss.n6124 5.91
R15283 vss.n6216 vss.n6213 5.91
R15284 vss.n16760 vss.n16759 5.91
R15285 vss.n16801 vss.n16800 5.91
R15286 vss.n16990 vss.n16989 5.91
R15287 vss.n17035 vss.n17034 5.91
R15288 vss.n17226 vss.n17225 5.91
R15289 vss.n17290 vss.n17289 5.91
R15290 vss.n16039 vss.n16036 5.91
R15291 vss.n16083 vss.n16080 5.91
R15292 vss.n15243 vss.n15242 5.91
R15293 vss.n15221 vss.n15220 5.91
R15294 vss.n15510 vss.n15509 5.91
R15295 vss.n15557 vss.n15556 5.91
R15296 vss.n15746 vss.n15745 5.91
R15297 vss.n15787 vss.n15786 5.91
R15298 vss.n16457 vss.n16456 5.91
R15299 vss.n16504 vss.n16503 5.91
R15300 vss.n21852 vss.n21850 5.896
R15301 vss.n21743 vss.n21713 5.896
R15302 vss.n3801 vss.n3799 5.896
R15303 vss.n3692 vss.n3662 5.896
R15304 vss.n10490 vss.n10489 5.88
R15305 vss.n10520 vss.n10519 5.88
R15306 vss.n10537 vss.n10533 5.851
R15307 vss.n12990 vss.n12986 5.851
R15308 vss.n12980 vss.n12976 5.851
R15309 vss.n14585 vss.n14581 5.851
R15310 vss.n14721 vss.n14717 5.851
R15311 vss.n14585 vss.n14583 5.851
R15312 vss.n14993 vss.n14989 5.851
R15313 vss.n14721 vss.n14719 5.851
R15314 vss.n12949 vss.n12945 5.851
R15315 vss.n13160 vss.n13156 5.851
R15316 vss.n13947 vss.n13945 5.851
R15317 vss.n13784 vss.n13780 5.851
R15318 vss.n13795 vss.n13791 5.851
R15319 vss.n13947 vss.n13946 5.851
R15320 vss.n11685 vss.n11682 5.851
R15321 vss.n11551 vss.n11547 5.851
R15322 vss.n11520 vss.n11516 5.851
R15323 vss.n11685 vss.n11684 5.851
R15324 vss.n12259 vss.n12257 5.851
R15325 vss.n11935 vss.n11932 5.851
R15326 vss.n11935 vss.n11934 5.851
R15327 vss.n14161 vss.n14157 5.851
R15328 vss.n14118 vss.n14114 5.851
R15329 vss.n13737 vss.n13733 5.851
R15330 vss.n11434 vss.n11430 5.851
R15331 vss.n11874 vss.n11870 5.851
R15332 vss.n11910 vss.n11906 5.851
R15333 vss.n12390 vss.n12386 5.851
R15334 vss.n12363 vss.n12359 5.851
R15335 vss.n10694 vss.n10690 5.851
R15336 vss.n10704 vss.n10700 5.851
R15337 vss.n13417 vss.n13413 5.851
R15338 vss.n13496 vss.n13492 5.851
R15339 vss.n13076 vss.n13072 5.851
R15340 vss.n10629 vss.n10625 5.851
R15341 vss.n10789 vss.n10785 5.851
R15342 vss.n12297 vss.n12293 5.851
R15343 vss.n12259 vss.n12258 5.851
R15344 vss.n22601 vss.n22597 5.794
R15345 vss.n22582 vss.n22578 5.794
R15346 vss.n22393 vss.n22389 5.794
R15347 vss.n22374 vss.n22370 5.794
R15348 vss.n22185 vss.n22181 5.794
R15349 vss.n22166 vss.n22162 5.794
R15350 vss.n21529 vss.n21525 5.794
R15351 vss.n21510 vss.n21506 5.794
R15352 vss.n21321 vss.n21317 5.794
R15353 vss.n21302 vss.n21298 5.794
R15354 vss.n21113 vss.n21109 5.794
R15355 vss.n21094 vss.n21090 5.794
R15356 vss.n20905 vss.n20901 5.794
R15357 vss.n12054 vss.n12051 5.794
R15358 vss.n12044 vss.n12041 5.794
R15359 vss.n10973 vss.n10970 5.794
R15360 vss.n10983 vss.n10980 5.794
R15361 vss.n13836 vss.n13833 5.794
R15362 vss.n13826 vss.n13823 5.794
R15363 vss.n11128 vss.n11125 5.794
R15364 vss.n11118 vss.n11115 5.794
R15365 vss.n13367 vss.n13364 5.794
R15366 vss.n13387 vss.n13384 5.794
R15367 vss.n14199 vss.n14196 5.794
R15368 vss.n14209 vss.n14206 5.794
R15369 vss.n12892 vss.n12889 5.794
R15370 vss.n12884 vss.n12883 5.794
R15371 vss.n12483 vss.n12480 5.794
R15372 vss.n12475 vss.n12474 5.794
R15373 vss.n8764 vss.n8760 5.794
R15374 vss.n8745 vss.n8741 5.794
R15375 vss.n8556 vss.n8552 5.794
R15376 vss.n8537 vss.n8533 5.794
R15377 vss.n8348 vss.n8344 5.794
R15378 vss.n8329 vss.n8325 5.794
R15379 vss.n8140 vss.n8136 5.794
R15380 vss.n8121 vss.n8117 5.794
R15381 vss.n7932 vss.n7928 5.794
R15382 vss.n7913 vss.n7909 5.794
R15383 vss.n7723 vss.n7719 5.794
R15384 vss.n7704 vss.n7700 5.794
R15385 vss.n7515 vss.n7511 5.794
R15386 vss.n14992 vss.n14990 5.75
R15387 vss.n10536 vss.n10534 5.75
R15388 vss.n14407 vss.n14406 5.705
R15389 vss.n13305 vss.n13304 5.705
R15390 vss.n14404 vss.n14403 5.683
R15391 vss.n11056 vss.n11055 5.683
R15392 vss.n13302 vss.n13292 5.683
R15393 vss.n12587 vss.n12577 5.683
R15394 vss.n20533 vss.n20522 5.647
R15395 vss.n20560 vss.n20549 5.647
R15396 vss.n20762 vss.n20751 5.647
R15397 vss.n20782 vss.n20771 5.647
R15398 vss.n12121 vss.n12114 5.647
R15399 vss.n12131 vss.n12124 5.647
R15400 vss.n10881 vss.n10874 5.647
R15401 vss.n11949 vss.n11942 5.647
R15402 vss.n14420 vss.n14413 5.647
R15403 vss.n14374 vss.n14367 5.647
R15404 vss.n11638 vss.n11631 5.647
R15405 vss.n11665 vss.n11658 5.647
R15406 vss.n13275 vss.n13268 5.647
R15407 vss.n13259 vss.n13252 5.647
R15408 vss.n13544 vss.n13537 5.647
R15409 vss.n14596 vss.n14589 5.647
R15410 vss.n14836 vss.n14829 5.647
R15411 vss.n14864 vss.n14857 5.647
R15412 vss.n10489 vss.n10482 5.647
R15413 vss.n10519 vss.n10512 5.647
R15414 vss.n7143 vss.n7132 5.647
R15415 vss.n7170 vss.n7159 5.647
R15416 vss.n7372 vss.n7361 5.647
R15417 vss.n7392 vss.n7381 5.647
R15418 vss.n1759 vss.n1748 5.647
R15419 vss.n1779 vss.n1768 5.647
R15420 vss.n1990 vss.n1977 5.647
R15421 vss.n2019 vss.n2006 5.647
R15422 vss.n2235 vss.n2222 5.647
R15423 vss.n2263 vss.n2250 5.647
R15424 vss.n2479 vss.n2466 5.647
R15425 vss.n2507 vss.n2494 5.647
R15426 vss.n2724 vss.n2711 5.647
R15427 vss.n2752 vss.n2739 5.647
R15428 vss.n2962 vss.n2949 5.647
R15429 vss.n2990 vss.n2977 5.647
R15430 vss.n3206 vss.n3193 5.647
R15431 vss.n3235 vss.n3222 5.647
R15432 vss.n15208 vss.n15197 5.647
R15433 vss.n15188 vss.n15177 5.647
R15434 vss.n220 vss.n209 5.647
R15435 vss.n240 vss.n229 5.647
R15436 vss.n451 vss.n438 5.647
R15437 vss.n480 vss.n467 5.647
R15438 vss.n696 vss.n683 5.647
R15439 vss.n724 vss.n711 5.647
R15440 vss.n940 vss.n927 5.647
R15441 vss.n968 vss.n955 5.647
R15442 vss.n1185 vss.n1172 5.647
R15443 vss.n1213 vss.n1200 5.647
R15444 vss.n23308 vss.n23295 5.647
R15445 vss.n23280 vss.n23267 5.647
R15446 vss.n23064 vss.n23051 5.647
R15447 vss.n23035 vss.n23022 5.647
R15448 vss.n1401 vss.n1390 5.647
R15449 vss.n22822 vss.n22811 5.647
R15450 vss.n12468 vss.n12458 5.611
R15451 bandgapmd_0.pnp_groupm_0.vss vss.n14820 5.584
R15452 vss.n12442 vss.t172 5.548
R15453 vss.n14020 vss.t166 5.548
R15454 vss.n21752 vss.n21708 5.495
R15455 vss.n3701 vss.n3657 5.495
R15456 vss.n9066 vss.n9065 5.449
R15457 vss.n9143 vss.n9142 5.449
R15458 vss.n10550 vss.n10549 5.337
R15459 vss.n15795 vss.n15794 5.325
R15460 vss.n10191 vss.n10190 5.307
R15461 vss.n22082 vss.n22070 5.307
R15462 vss.n22068 vss.n21607 5.282
R15463 vss.n4018 vss.n3556 5.282
R15464 vss.n21787 vss.n21774 5.282
R15465 vss.n3736 vss.n3723 5.282
R15466 vss.n22000 vss.n21999 5.28
R15467 vss.n3949 vss.n3948 5.28
R15468 vss.n20642 vss.n20641 5.27
R15469 vss.n20660 vss.n20659 5.27
R15470 vss.n21848 vss.n21847 5.27
R15471 vss.n21673 vss.n21662 5.27
R15472 vss.n12065 vss.n12064 5.27
R15473 vss.n10794 vss.n10793 5.27
R15474 vss.n10957 vss.n10956 5.27
R15475 vss.n10997 vss.n10996 5.27
R15476 vss.n13847 vss.n13846 5.27
R15477 vss.n14068 vss.n14067 5.27
R15478 vss.n11714 vss.n11713 5.27
R15479 vss.n11058 vss.n11057 5.27
R15480 vss.n13345 vss.n13344 5.27
R15481 vss.n14690 vss.n14689 5.27
R15482 vss.n14183 vss.n14182 5.27
R15483 vss.n14225 vss.n14224 5.27
R15484 vss.n12865 vss.n12864 5.27
R15485 vss.n12908 vss.n12907 5.27
R15486 vss.n12460 vss.n12459 5.27
R15487 vss.n12495 vss.n12494 5.27
R15488 vss.n3797 vss.n3796 5.27
R15489 vss.n3622 vss.n3611 5.27
R15490 vss.n7252 vss.n7251 5.27
R15491 vss.n7270 vss.n7269 5.27
R15492 vss.n1863 vss.n1862 5.27
R15493 vss.n1881 vss.n1880 5.27
R15494 vss.n2107 vss.n2106 5.27
R15495 vss.n2125 vss.n2124 5.27
R15496 vss.n2351 vss.n2350 5.27
R15497 vss.n2369 vss.n2368 5.27
R15498 vss.n2595 vss.n2594 5.27
R15499 vss.n2614 vss.n2613 5.27
R15500 vss.n1546 vss.n1545 5.27
R15501 vss.n2844 vss.n2843 5.27
R15502 vss.n2852 vss.n2851 5.27
R15503 vss.n3078 vss.n3077 5.27
R15504 vss.n3096 vss.n3095 5.27
R15505 vss.n3322 vss.n3321 5.27
R15506 vss.n3341 vss.n3340 5.27
R15507 vss.n324 vss.n323 5.27
R15508 vss.n342 vss.n341 5.27
R15509 vss.n568 vss.n567 5.27
R15510 vss.n586 vss.n585 5.27
R15511 vss.n812 vss.n811 5.27
R15512 vss.n830 vss.n829 5.27
R15513 vss.n1056 vss.n1055 5.27
R15514 vss.n1075 vss.n1074 5.27
R15515 vss.n1301 vss.n1300 5.27
R15516 vss.n23395 vss.n23394 5.27
R15517 vss.n23170 vss.n23169 5.27
R15518 vss.n23152 vss.n23151 5.27
R15519 vss.n22926 vss.n22925 5.27
R15520 vss.n22908 vss.n22907 5.27
R15521 vss.n21767 vss.n21696 5.268
R15522 vss.n21681 vss.n21663 5.268
R15523 vss.n3716 vss.n3645 5.268
R15524 vss.n3630 vss.n3612 5.268
R15525 vss.n21995 vss.n21994 5.268
R15526 vss.n3944 vss.n3943 5.268
R15527 vss.n21765 vss.n21696 5.267
R15528 vss.n21678 vss.n21663 5.267
R15529 vss.n3714 vss.n3645 5.267
R15530 vss.n3627 vss.n3612 5.267
R15531 vss.n3477 vss.n3476 5.148
R15532 vss.n1452 vss.n1451 5.148
R15533 vss.n13924 vss.n13923 5
R15534 vss.n13612 vss.n13610 5
R15535 vss.n11023 vss.n11022 5
R15536 vss.n11270 vss.n11269 5
R15537 vss.n10915 vss.n10914 5
R15538 vss.n10835 vss.n10834 5
R15539 vss.n12236 vss.n12235 5
R15540 vss.n12518 vss.n12516 5
R15541 vss.n10597 vss.n10596 5
R15542 vss.n10496 vss.n10494 5
R15543 vss.n13197 vss.n13196 5
R15544 vss.n13435 vss.n13434 5
R15545 vss.n13622 vss.n13620 5
R15546 vss.n13426 vss.n13425 5
R15547 vss.n10589 vss.n10587 5
R15548 vss.n11402 vss.n11401 5
R15549 vss.n11394 vss.n11392 5
R15550 vss.n11650 vss.n11649 5
R15551 vss.n3489 vss.n3478 4.919
R15552 vss.n1464 vss.n1453 4.919
R15553 vss.n20515 vss.n20507 4.894
R15554 vss.n20575 vss.n20567 4.894
R15555 vss.n20743 vss.n20735 4.894
R15556 vss.n20797 vss.n20789 4.894
R15557 vss.n12145 vss.n12138 4.894
R15558 vss.n11977 vss.n11970 4.894
R15559 vss.n11923 vss.n11916 4.894
R15560 vss.n14339 vss.n14332 4.894
R15561 vss.n11627 vss.n11620 4.894
R15562 vss.n11676 vss.n11669 4.894
R15563 vss.n14817 vss.n14810 4.894
R15564 vss.n14616 vss.n14609 4.894
R15565 vss.n14556 vss.n14549 4.894
R15566 vss.n14907 vss.n14900 4.894
R15567 vss.n10549 vss.n10542 4.894
R15568 vss.n7125 vss.n7117 4.894
R15569 vss.n7185 vss.n7177 4.894
R15570 vss.n7353 vss.n7345 4.894
R15571 vss.n7407 vss.n7399 4.894
R15572 vss.n1737 vss.n1729 4.894
R15573 vss.n1796 vss.n1788 4.894
R15574 vss.n1970 vss.n1961 4.894
R15575 vss.n2035 vss.n2026 4.894
R15576 vss.n2215 vss.n2206 4.894
R15577 vss.n2279 vss.n2270 4.894
R15578 vss.n2459 vss.n2450 4.894
R15579 vss.n2524 vss.n2515 4.894
R15580 vss.n2703 vss.n2694 4.894
R15581 vss.n2768 vss.n2759 4.894
R15582 vss.n2942 vss.n2933 4.894
R15583 vss.n3006 vss.n2997 4.894
R15584 vss.n3186 vss.n3177 4.894
R15585 vss.n3251 vss.n3242 4.894
R15586 vss.n3424 vss.n3416 4.894
R15587 vss.n3465 vss.n3457 4.894
R15588 vss.n198 vss.n190 4.894
R15589 vss.n257 vss.n249 4.894
R15590 vss.n431 vss.n422 4.894
R15591 vss.n496 vss.n487 4.894
R15592 vss.n676 vss.n667 4.894
R15593 vss.n740 vss.n731 4.894
R15594 vss.n920 vss.n911 4.894
R15595 vss.n985 vss.n976 4.894
R15596 vss.n1164 vss.n1155 4.894
R15597 vss.n1229 vss.n1220 4.894
R15598 vss.n23324 vss.n23315 4.894
R15599 vss.n23260 vss.n23251 4.894
R15600 vss.n23080 vss.n23071 4.894
R15601 vss.n23015 vss.n23006 4.894
R15602 vss.n22839 vss.n22831 4.894
R15603 vss.n1440 vss.n1432 4.894
R15604 vss.n20338 vss.n17598 4.884
R15605 vss.n20339 vss.n20338 4.884
R15606 vss.n6948 vss.n4208 4.884
R15607 vss.n6949 vss.n6948 4.884
R15608 vss.n22694 vss.n22692 4.835
R15609 vss.n22694 vss.n22693 4.835
R15610 vss.n22486 vss.n22484 4.835
R15611 vss.n22486 vss.n22485 4.835
R15612 vss.n22278 vss.n22276 4.835
R15613 vss.n22278 vss.n22277 4.835
R15614 vss.n22084 vss.n22083 4.835
R15615 vss.n21414 vss.n21412 4.835
R15616 vss.n21414 vss.n21413 4.835
R15617 vss.n21206 vss.n21204 4.835
R15618 vss.n21206 vss.n21205 4.835
R15619 vss.n20998 vss.n20996 4.835
R15620 vss.n20998 vss.n20997 4.835
R15621 vss.n8857 vss.n8855 4.835
R15622 vss.n8857 vss.n8856 4.835
R15623 vss.n8649 vss.n8647 4.835
R15624 vss.n8649 vss.n8648 4.835
R15625 vss.n8441 vss.n8439 4.835
R15626 vss.n8441 vss.n8440 4.835
R15627 vss.n8247 vss.n8245 4.835
R15628 vss.n8247 vss.n8246 4.835
R15629 vss.n8025 vss.n8023 4.835
R15630 vss.n8025 vss.n8024 4.835
R15631 vss.n7816 vss.n7814 4.835
R15632 vss.n7816 vss.n7815 4.835
R15633 vss.n7608 vss.n7606 4.835
R15634 vss.n7608 vss.n7607 4.835
R15635 vss.n21719 vss.n21688 4.734
R15636 vss.n3668 vss.n3637 4.734
R15637 vss.n21824 vss.n21823 4.734
R15638 vss.n3773 vss.n3772 4.734
R15639 vss.n19015 vss.n19014 4.711
R15640 vss.n19014 vss.n19013 4.711
R15641 vss.n18889 vss.n17734 4.711
R15642 vss.n18889 vss.n17735 4.711
R15643 vss.n18768 vss.n18767 4.711
R15644 vss.n18767 vss.n17842 4.711
R15645 vss.n18648 vss.n17947 4.711
R15646 vss.n18648 vss.n17948 4.711
R15647 vss.n18527 vss.n18526 4.711
R15648 vss.n18526 vss.n18055 4.711
R15649 vss.n18407 vss.n18160 4.711
R15650 vss.n18407 vss.n18161 4.711
R15651 vss.n18286 vss.n18285 4.711
R15652 vss.n18285 vss.n18268 4.711
R15653 vss.n20280 vss.n19034 4.711
R15654 vss.n20280 vss.n20279 4.711
R15655 vss.n20161 vss.n20160 4.711
R15656 vss.n20160 vss.n20159 4.711
R15657 vss.n20035 vss.n19241 4.711
R15658 vss.n20035 vss.n19242 4.711
R15659 vss.n19914 vss.n19913 4.711
R15660 vss.n19913 vss.n19912 4.711
R15661 vss.n19788 vss.n19448 4.711
R15662 vss.n19788 vss.n19449 4.711
R15663 vss.n19667 vss.n19666 4.711
R15664 vss.n19666 vss.n19665 4.711
R15665 vss.n5625 vss.n5624 4.711
R15666 vss.n5624 vss.n5623 4.711
R15667 vss.n5499 vss.n4344 4.711
R15668 vss.n5499 vss.n4345 4.711
R15669 vss.n5378 vss.n5377 4.711
R15670 vss.n5377 vss.n4452 4.711
R15671 vss.n5258 vss.n4557 4.711
R15672 vss.n5258 vss.n4558 4.711
R15673 vss.n5137 vss.n5136 4.711
R15674 vss.n5136 vss.n4665 4.711
R15675 vss.n5017 vss.n4770 4.711
R15676 vss.n5017 vss.n4771 4.711
R15677 vss.n4896 vss.n4895 4.711
R15678 vss.n4895 vss.n4878 4.711
R15679 vss.n6890 vss.n5644 4.711
R15680 vss.n6890 vss.n6889 4.711
R15681 vss.n6771 vss.n6770 4.711
R15682 vss.n6770 vss.n6769 4.711
R15683 vss.n6645 vss.n5851 4.711
R15684 vss.n6645 vss.n5852 4.711
R15685 vss.n6524 vss.n6523 4.711
R15686 vss.n6523 vss.n6522 4.711
R15687 vss.n6398 vss.n6058 4.711
R15688 vss.n6398 vss.n6059 4.711
R15689 vss.n6277 vss.n6276 4.711
R15690 vss.n6276 vss.n6275 4.711
R15691 vss.n10858 vss.n10857 4.684
R15692 vss.n14013 vss.n14012 4.684
R15693 vss.n13534 vss.n13533 4.684
R15694 vss.n1693 vss.n1682 4.681
R15695 vss.n154 vss.n143 4.681
R15696 vss.n16302 vss.n16301 4.655
R15697 vss.n12280 vss.n12279 4.65
R15698 vss.n13479 vss.n13478 4.65
R15699 vss.n10720 vss.n10719 4.65
R15700 vss.n13010 vss.n13009 4.65
R15701 vss.n12379 vss.n12378 4.65
R15702 vss.n11539 vss.n11538 4.65
R15703 vss.n19014 vss.n17631 4.65
R15704 vss.n18890 vss.n18889 4.65
R15705 vss.n18767 vss.n18766 4.65
R15706 vss.n18649 vss.n18648 4.65
R15707 vss.n18526 vss.n18525 4.65
R15708 vss.n18408 vss.n18407 4.65
R15709 vss.n18285 vss.n18284 4.65
R15710 vss.n19619 vss.n19589 4.65
R15711 vss.n20280 vss.n19033 4.65
R15712 vss.n20160 vss.n19142 4.65
R15713 vss.n20036 vss.n20035 4.65
R15714 vss.n19913 vss.n19349 4.65
R15715 vss.n19789 vss.n19788 4.65
R15716 vss.n19666 vss.n19556 4.65
R15717 vss.n20443 vss.n20442 4.65
R15718 vss.n20542 vss.n20541 4.65
R15719 vss.n20768 vss.n20767 4.65
R15720 vss.n20892 vss.n20891 4.65
R15721 vss.n21577 vss.n17408 4.65
R15722 vss.n21574 vss.n21573 4.65
R15723 vss.n21560 vss.n21559 4.65
R15724 vss.n21546 vss.n21545 4.65
R15725 vss.n21532 vss.n21531 4.65
R15726 vss.n21514 vss.n21513 4.65
R15727 vss.n21500 vss.n21499 4.65
R15728 vss.n21486 vss.n21485 4.65
R15729 vss.n21472 vss.n21471 4.65
R15730 vss.n21458 vss.n21457 4.65
R15731 vss.n21444 vss.n21443 4.65
R15732 vss.n21430 vss.n21429 4.65
R15733 vss.n21415 vss.n21414 4.65
R15734 vss.n21410 vss.n21409 4.65
R15735 vss.n21394 vss.n21393 4.65
R15736 vss.n21380 vss.n21379 4.65
R15737 vss.n21366 vss.n21365 4.65
R15738 vss.n21352 vss.n21351 4.65
R15739 vss.n21338 vss.n21337 4.65
R15740 vss.n21324 vss.n21323 4.65
R15741 vss.n21306 vss.n21305 4.65
R15742 vss.n21292 vss.n21291 4.65
R15743 vss.n21278 vss.n21277 4.65
R15744 vss.n21264 vss.n21263 4.65
R15745 vss.n21250 vss.n21249 4.65
R15746 vss.n21236 vss.n21235 4.65
R15747 vss.n21222 vss.n21221 4.65
R15748 vss.n21207 vss.n21206 4.65
R15749 vss.n21202 vss.n21201 4.65
R15750 vss.n21186 vss.n21185 4.65
R15751 vss.n21172 vss.n21171 4.65
R15752 vss.n21158 vss.n21157 4.65
R15753 vss.n21144 vss.n21143 4.65
R15754 vss.n21130 vss.n21129 4.65
R15755 vss.n21116 vss.n21115 4.65
R15756 vss.n21098 vss.n21097 4.65
R15757 vss.n21084 vss.n21083 4.65
R15758 vss.n21070 vss.n21069 4.65
R15759 vss.n21056 vss.n21055 4.65
R15760 vss.n21042 vss.n21041 4.65
R15761 vss.n21028 vss.n21027 4.65
R15762 vss.n21014 vss.n21013 4.65
R15763 vss.n20999 vss.n20998 4.65
R15764 vss.n20994 vss.n20993 4.65
R15765 vss.n20978 vss.n20977 4.65
R15766 vss.n20964 vss.n20963 4.65
R15767 vss.n20950 vss.n20949 4.65
R15768 vss.n20936 vss.n20935 4.65
R15769 vss.n20922 vss.n20921 4.65
R15770 vss.n20908 vss.n20907 4.65
R15771 vss.n22085 vss.n22084 4.65
R15772 vss.n10208 vss.n10207 4.65
R15773 vss.n10202 vss.n10201 4.65
R15774 vss.n10196 vss.n10195 4.65
R15775 vss.n10190 vss.n10187 4.65
R15776 vss.n9703 vss.n9702 4.65
R15777 vss.n9720 vss.n9719 4.65
R15778 vss.n9726 vss.n9725 4.65
R15779 vss.n9732 vss.n9731 4.65
R15780 vss.n9738 vss.n9737 4.65
R15781 vss.n9744 vss.n9743 4.65
R15782 vss.n10183 vss.n10182 4.65
R15783 vss.n12950 vss.n12949 4.65
R15784 vss.n12949 vss.n12948 4.65
R15785 vss.n13161 vss.n13160 4.65
R15786 vss.n13160 vss.n13159 4.65
R15787 vss.n12588 vss.n12574 4.65
R15788 vss.n12147 vss.n12109 4.65
R15789 vss.n11954 vss.n10910 4.65
R15790 vss.n11169 vss.n11168 4.65
R15791 vss.n11099 vss.n11098 4.65
R15792 vss.n11101 vss.n11100 4.65
R15793 vss.n11470 vss.n11469 4.65
R15794 vss.n11480 vss.n11479 4.65
R15795 vss.n11479 vss.n11478 4.65
R15796 vss.n13678 vss.n13677 4.65
R15797 vss.n13669 vss.n13668 4.65
R15798 vss.n13668 vss.n13667 4.65
R15799 vss.n12991 vss.n12990 4.65
R15800 vss.n12990 vss.n12989 4.65
R15801 vss.n12981 vss.n12980 4.65
R15802 vss.n12980 vss.n12979 4.65
R15803 vss.n13137 vss.n13136 4.65
R15804 vss.n13120 vss.n13119 4.65
R15805 vss.n13119 vss.n13118 4.65
R15806 vss.n13128 vss.n13127 4.65
R15807 vss.n13147 vss.n13146 4.65
R15808 vss.n13146 vss.n13145 4.65
R15809 vss.n12713 vss.n10538 4.65
R15810 vss.n10665 vss.n10664 4.65
R15811 vss.n12412 vss.n12411 4.65
R15812 vss.n12411 vss.n12410 4.65
R15813 vss.n12402 vss.n12401 4.65
R15814 vss.n12401 vss.n12400 4.65
R15815 vss.n12364 vss.n12363 4.65
R15816 vss.n12363 vss.n12362 4.65
R15817 vss.n12391 vss.n12390 4.65
R15818 vss.n12390 vss.n12389 4.65
R15819 vss.n10675 vss.n10674 4.65
R15820 vss.n10674 vss.n10673 4.65
R15821 vss.n11462 vss.n11461 4.65
R15822 vss.n10657 vss.n10656 4.65
R15823 vss.n10695 vss.n10694 4.65
R15824 vss.n10694 vss.n10693 4.65
R15825 vss.n10705 vss.n10704 4.65
R15826 vss.n10704 vss.n10703 4.65
R15827 vss.n12329 vss.n12328 4.65
R15828 vss.n12328 vss.n12327 4.65
R15829 vss.n11490 vss.n11489 4.65
R15830 vss.n11489 vss.n11488 4.65
R15831 vss.n13464 vss.n13463 4.65
R15832 vss.n13084 vss.n13083 4.65
R15833 vss.n13068 vss.n13067 4.65
R15834 vss.n10621 vss.n10620 4.65
R15835 vss.n10637 vss.n10636 4.65
R15836 vss.n12306 vss.n12305 4.65
R15837 vss.n13418 vss.n13417 4.65
R15838 vss.n13417 vss.n13416 4.65
R15839 vss.n13497 vss.n13496 4.65
R15840 vss.n13496 vss.n13495 4.65
R15841 vss.n13467 vss.n13466 4.65
R15842 vss.n13462 vss.n13461 4.65
R15843 vss.n13461 vss.n13460 4.65
R15844 vss.n13460 vss.n13459 4.65
R15845 vss.n13449 vss.n13448 4.65
R15846 vss.n13448 vss.n13447 4.65
R15847 vss.n13024 vss.n13023 4.65
R15848 vss.n13023 vss.n13022 4.65
R15849 vss.n13093 vss.n13092 4.65
R15850 vss.n13092 vss.n13091 4.65
R15851 vss.n13091 vss.n13090 4.65
R15852 vss.n13081 vss.n13080 4.65
R15853 vss.n13078 vss.n13077 4.65
R15854 vss.n13077 vss.n13076 4.65
R15855 vss.n13076 vss.n13075 4.65
R15856 vss.n13065 vss.n13064 4.65
R15857 vss.n10601 vss.n10600 4.65
R15858 vss.n10631 vss.n10630 4.65
R15859 vss.n10630 vss.n10629 4.65
R15860 vss.n10629 vss.n10628 4.65
R15861 vss.n10634 vss.n10633 4.65
R15862 vss.n10646 vss.n10645 4.65
R15863 vss.n10645 vss.n10644 4.65
R15864 vss.n10644 vss.n10643 4.65
R15865 vss.n10581 vss.n10580 4.65
R15866 vss.n10580 vss.n10579 4.65
R15867 vss.n10738 vss.n10737 4.65
R15868 vss.n10737 vss.n10736 4.65
R15869 vss.n12315 vss.n12314 4.65
R15870 vss.n12314 vss.n12313 4.65
R15871 vss.n12313 vss.n12312 4.65
R15872 vss.n12303 vss.n12302 4.65
R15873 vss.n10790 vss.n10789 4.65
R15874 vss.n10789 vss.n10788 4.65
R15875 vss.n12298 vss.n12297 4.65
R15876 vss.n12297 vss.n12296 4.65
R15877 vss.n10811 vss.n10810 4.65
R15878 vss.n10810 vss.n10809 4.65
R15879 vss.n12034 vss.n12033 4.65
R15880 vss.n12033 vss.n12032 4.65
R15881 vss.n12264 vss.n12263 4.65
R15882 vss.n14153 vss.n14152 4.65
R15883 vss.n14122 vss.n14121 4.65
R15884 vss.n14106 vss.n14105 4.65
R15885 vss.n13745 vss.n13744 4.65
R15886 vss.n13729 vss.n13728 4.65
R15887 vss.n11426 vss.n11425 4.65
R15888 vss.n11442 vss.n11441 4.65
R15889 vss.n11862 vss.n11861 4.65
R15890 vss.n11878 vss.n11877 4.65
R15891 vss.n11902 vss.n11901 4.65
R15892 vss.n14163 vss.n14162 4.65
R15893 vss.n14162 vss.n14161 4.65
R15894 vss.n14161 vss.n14160 4.65
R15895 vss.n14143 vss.n14142 4.65
R15896 vss.n14141 vss.n14140 4.65
R15897 vss.n14120 vss.n14119 4.65
R15898 vss.n14119 vss.n14118 4.65
R15899 vss.n14118 vss.n14117 4.65
R15900 vss.n14109 vss.n14108 4.65
R15901 vss.n14104 vss.n14103 4.65
R15902 vss.n14103 vss.n14102 4.65
R15903 vss.n14102 vss.n14101 4.65
R15904 vss.n13636 vss.n13635 4.65
R15905 vss.n13635 vss.n13634 4.65
R15906 vss.n13688 vss.n13687 4.65
R15907 vss.n13687 vss.n13686 4.65
R15908 vss.n13754 vss.n13753 4.65
R15909 vss.n13753 vss.n13752 4.65
R15910 vss.n13752 vss.n13751 4.65
R15911 vss.n13742 vss.n13741 4.65
R15912 vss.n13739 vss.n13738 4.65
R15913 vss.n13738 vss.n13737 4.65
R15914 vss.n13737 vss.n13736 4.65
R15915 vss.n13726 vss.n13725 4.65
R15916 vss.n11407 vss.n11406 4.65
R15917 vss.n11436 vss.n11435 4.65
R15918 vss.n11435 vss.n11434 4.65
R15919 vss.n11434 vss.n11433 4.65
R15920 vss.n11439 vss.n11438 4.65
R15921 vss.n11451 vss.n11450 4.65
R15922 vss.n11450 vss.n11449 4.65
R15923 vss.n11449 vss.n11448 4.65
R15924 vss.n11385 vss.n11384 4.65
R15925 vss.n11384 vss.n11383 4.65
R15926 vss.n11371 vss.n11370 4.65
R15927 vss.n11370 vss.n11369 4.65
R15928 vss.n11860 vss.n11859 4.65
R15929 vss.n11859 vss.n11858 4.65
R15930 vss.n11858 vss.n11857 4.65
R15931 vss.n11865 vss.n11864 4.65
R15932 vss.n11876 vss.n11875 4.65
R15933 vss.n11875 vss.n11874 4.65
R15934 vss.n11874 vss.n11873 4.65
R15935 vss.n11881 vss.n11880 4.65
R15936 vss.n11883 vss.n11882 4.65
R15937 vss.n11912 vss.n11911 4.65
R15938 vss.n11911 vss.n11910 4.65
R15939 vss.n11910 vss.n11909 4.65
R15940 vss.n10936 vss.n10935 4.65
R15941 vss.n10935 vss.n10934 4.65
R15942 vss.n11314 vss.n11313 4.65
R15943 vss.n11313 vss.n11312 4.65
R15944 vss.n11940 vss.n11939 4.65
R15945 vss.n13656 vss.n13655 4.65
R15946 vss.n13655 vss.n13654 4.65
R15947 vss.n13646 vss.n13645 4.65
R15948 vss.n13785 vss.n13784 4.65
R15949 vss.n13784 vss.n13783 4.65
R15950 vss.n13796 vss.n13795 4.65
R15951 vss.n13795 vss.n13794 4.65
R15952 vss.n11552 vss.n11551 4.65
R15953 vss.n11551 vss.n11550 4.65
R15954 vss.n11521 vss.n11520 4.65
R15955 vss.n11520 vss.n11519 4.65
R15956 vss.n11817 vss.n11689 4.65
R15957 vss.n14385 vss.n14384 4.65
R15958 vss.n11653 vss.n11584 4.65
R15959 vss.n14065 vss.n14064 4.65
R15960 vss.n14064 vss.n14063 4.65
R15961 vss.n11698 vss.n11697 4.65
R15962 vss.n11697 vss.n11696 4.65
R15963 vss.n13962 vss.n13961 4.65
R15964 vss.n13961 vss.n13960 4.65
R15965 vss.n11815 vss.n11814 4.65
R15966 vss.n11814 vss.n11813 4.65
R15967 vss.n13950 vss.n13949 4.65
R15968 vss.n14410 vss.n14409 4.65
R15969 vss.n14268 vss.n14267 4.65
R15970 vss.n14266 vss.n14265 4.65
R15971 vss.n14602 vss.n13591 4.65
R15972 vss.n14712 vss.n14711 4.65
R15973 vss.n14711 vss.n14710 4.65
R15974 vss.n13378 vss.n13377 4.65
R15975 vss.n13377 vss.n13376 4.65
R15976 vss.n14723 vss.n14722 4.65
R15977 vss.n14576 vss.n14575 4.65
R15978 vss.n14575 vss.n14574 4.65
R15979 vss.n14566 vss.n14565 4.65
R15980 vss.n14565 vss.n14564 4.65
R15981 vss.n14587 vss.n14586 4.65
R15982 vss.n15006 vss.n14995 4.65
R15983 vss.n13308 vss.n13307 4.65
R15984 vss.n15004 vss.n15003 4.65
R15985 vss.n15003 vss.n15002 4.65
R15986 vss.n14985 vss.n14984 4.65
R15987 vss.n14984 vss.n14983 4.65
R15988 vss.n14820 vss.n14819 4.65
R15989 vss.n5624 vss.n4241 4.65
R15990 vss.n5500 vss.n5499 4.65
R15991 vss.n5377 vss.n5376 4.65
R15992 vss.n5259 vss.n5258 4.65
R15993 vss.n5136 vss.n5135 4.65
R15994 vss.n5018 vss.n5017 4.65
R15995 vss.n4895 vss.n4894 4.65
R15996 vss.n6229 vss.n6199 4.65
R15997 vss.n6890 vss.n5643 4.65
R15998 vss.n6770 vss.n5752 4.65
R15999 vss.n6646 vss.n6645 4.65
R16000 vss.n6523 vss.n5959 4.65
R16001 vss.n6399 vss.n6398 4.65
R16002 vss.n6276 vss.n6166 4.65
R16003 vss.n7053 vss.n7052 4.65
R16004 vss.n7152 vss.n7151 4.65
R16005 vss.n7378 vss.n7377 4.65
R16006 vss.n7502 vss.n7501 4.65
R16007 vss.n8920 vss.n8919 4.65
R16008 vss.n8918 vss.n8917 4.65
R16009 vss.n8915 vss.n8914 4.65
R16010 vss.n8901 vss.n8900 4.65
R16011 vss.n8887 vss.n8886 4.65
R16012 vss.n8873 vss.n8872 4.65
R16013 vss.n8858 vss.n8857 4.65
R16014 vss.n8853 vss.n8852 4.65
R16015 vss.n8837 vss.n8836 4.65
R16016 vss.n8823 vss.n8822 4.65
R16017 vss.n8809 vss.n8808 4.65
R16018 vss.n8795 vss.n8794 4.65
R16019 vss.n8781 vss.n8780 4.65
R16020 vss.n8767 vss.n8766 4.65
R16021 vss.n8749 vss.n8748 4.65
R16022 vss.n8735 vss.n8734 4.65
R16023 vss.n8721 vss.n8720 4.65
R16024 vss.n8707 vss.n8706 4.65
R16025 vss.n8693 vss.n8692 4.65
R16026 vss.n8679 vss.n8678 4.65
R16027 vss.n8665 vss.n8664 4.65
R16028 vss.n8650 vss.n8649 4.65
R16029 vss.n8645 vss.n8644 4.65
R16030 vss.n8629 vss.n8628 4.65
R16031 vss.n8615 vss.n8614 4.65
R16032 vss.n8601 vss.n8600 4.65
R16033 vss.n8587 vss.n8586 4.65
R16034 vss.n8573 vss.n8572 4.65
R16035 vss.n8559 vss.n8558 4.65
R16036 vss.n8541 vss.n8540 4.65
R16037 vss.n8527 vss.n8526 4.65
R16038 vss.n8513 vss.n8512 4.65
R16039 vss.n8499 vss.n8498 4.65
R16040 vss.n8485 vss.n8484 4.65
R16041 vss.n8471 vss.n8470 4.65
R16042 vss.n8457 vss.n8456 4.65
R16043 vss.n8442 vss.n8441 4.65
R16044 vss.n8437 vss.n8436 4.65
R16045 vss.n8421 vss.n8420 4.65
R16046 vss.n8407 vss.n8406 4.65
R16047 vss.n8393 vss.n8392 4.65
R16048 vss.n8379 vss.n8378 4.65
R16049 vss.n8365 vss.n8364 4.65
R16050 vss.n8351 vss.n8350 4.65
R16051 vss.n8333 vss.n8332 4.65
R16052 vss.n8319 vss.n8318 4.65
R16053 vss.n8305 vss.n8304 4.65
R16054 vss.n8291 vss.n8290 4.65
R16055 vss.n8277 vss.n8276 4.65
R16056 vss.n8263 vss.n8262 4.65
R16057 vss.n8248 vss.n8247 4.65
R16058 vss.n8230 vss.n8229 4.65
R16059 vss.n8213 vss.n8212 4.65
R16060 vss.n8199 vss.n8198 4.65
R16061 vss.n8185 vss.n8184 4.65
R16062 vss.n8171 vss.n8170 4.65
R16063 vss.n8157 vss.n8156 4.65
R16064 vss.n8143 vss.n8142 4.65
R16065 vss.n8125 vss.n8124 4.65
R16066 vss.n8111 vss.n8110 4.65
R16067 vss.n8097 vss.n8096 4.65
R16068 vss.n8083 vss.n8082 4.65
R16069 vss.n8069 vss.n8068 4.65
R16070 vss.n8055 vss.n8054 4.65
R16071 vss.n8041 vss.n8040 4.65
R16072 vss.n8026 vss.n8025 4.65
R16073 vss.n8021 vss.n8020 4.65
R16074 vss.n8005 vss.n8004 4.65
R16075 vss.n7991 vss.n7990 4.65
R16076 vss.n7977 vss.n7976 4.65
R16077 vss.n7963 vss.n7962 4.65
R16078 vss.n7949 vss.n7948 4.65
R16079 vss.n7935 vss.n7934 4.65
R16080 vss.n7917 vss.n7916 4.65
R16081 vss.n7903 vss.n7902 4.65
R16082 vss.n7889 vss.n7888 4.65
R16083 vss.n7875 vss.n7874 4.65
R16084 vss.n7861 vss.n7860 4.65
R16085 vss.n7846 vss.n7845 4.65
R16086 vss.n7832 vss.n7831 4.65
R16087 vss.n7817 vss.n7816 4.65
R16088 vss.n7812 vss.n7811 4.65
R16089 vss.n7796 vss.n7795 4.65
R16090 vss.n7782 vss.n7781 4.65
R16091 vss.n7768 vss.n7767 4.65
R16092 vss.n7754 vss.n7753 4.65
R16093 vss.n7740 vss.n7739 4.65
R16094 vss.n7726 vss.n7725 4.65
R16095 vss.n7708 vss.n7707 4.65
R16096 vss.n7694 vss.n7693 4.65
R16097 vss.n7680 vss.n7679 4.65
R16098 vss.n7666 vss.n7665 4.65
R16099 vss.n7652 vss.n7651 4.65
R16100 vss.n7638 vss.n7637 4.65
R16101 vss.n7624 vss.n7623 4.65
R16102 vss.n7609 vss.n7608 4.65
R16103 vss.n7604 vss.n7603 4.65
R16104 vss.n7588 vss.n7587 4.65
R16105 vss.n7574 vss.n7573 4.65
R16106 vss.n7560 vss.n7559 4.65
R16107 vss.n7546 vss.n7545 4.65
R16108 vss.n7532 vss.n7531 4.65
R16109 vss.n7518 vss.n7517 4.65
R16110 vss.n1765 vss.n1764 4.65
R16111 vss.n2000 vss.n1999 4.65
R16112 vss.n2244 vss.n2243 4.65
R16113 vss.n2488 vss.n2487 4.65
R16114 vss.n2733 vss.n2732 4.65
R16115 vss.n2971 vss.n2970 4.65
R16116 vss.n3215 vss.n3214 4.65
R16117 vss.n15194 vss.n15193 4.65
R16118 vss.n15155 vss.n15154 4.65
R16119 vss.n16239 vss.n16238 4.65
R16120 vss.n16225 vss.n16224 4.65
R16121 vss.n16211 vss.n16210 4.65
R16122 vss.n16197 vss.n16196 4.65
R16123 vss.n16183 vss.n16182 4.65
R16124 vss.n16172 vss.n16171 4.65
R16125 vss.n16158 vss.n16157 4.65
R16126 vss.n16144 vss.n16143 4.65
R16127 vss.n16130 vss.n16129 4.65
R16128 vss.n16116 vss.n16115 4.65
R16129 vss.n16102 vss.n16101 4.65
R16130 vss.n16088 vss.n16087 4.65
R16131 vss.n16059 vss.n16058 4.65
R16132 vss.n16045 vss.n16044 4.65
R16133 vss.n16031 vss.n16030 4.65
R16134 vss.n16017 vss.n16016 4.65
R16135 vss.n16003 vss.n16002 4.65
R16136 vss.n15989 vss.n15988 4.65
R16137 vss.n15975 vss.n15974 4.65
R16138 vss.n15961 vss.n15960 4.65
R16139 vss.n15947 vss.n15946 4.65
R16140 vss.n15936 vss.n15935 4.65
R16141 vss.n15922 vss.n15921 4.65
R16142 vss.n15908 vss.n15907 4.65
R16143 vss.n15894 vss.n15893 4.65
R16144 vss.n15323 vss.n15322 4.65
R16145 vss.n15548 vss.n15547 4.65
R16146 vss.n15782 vss.n15781 4.65
R16147 vss.n16495 vss.n16494 4.65
R16148 vss.n16698 vss.n16697 4.65
R16149 vss.n16712 vss.n16711 4.65
R16150 vss.n16726 vss.n16725 4.65
R16151 vss.n16740 vss.n16739 4.65
R16152 vss.n16754 vss.n16753 4.65
R16153 vss.n16684 vss.n16683 4.65
R16154 vss.n16766 vss.n16765 4.65
R16155 vss.n16778 vss.n16777 4.65
R16156 vss.n16796 vss.n16795 4.65
R16157 vss.n16784 vss.n16783 4.65
R16158 vss.n16807 vss.n16806 4.65
R16159 vss.n16821 vss.n16820 4.65
R16160 vss.n16835 vss.n16834 4.65
R16161 vss.n16849 vss.n16848 4.65
R16162 vss.n16877 vss.n16876 4.65
R16163 vss.n16891 vss.n16890 4.65
R16164 vss.n16902 vss.n16901 4.65
R16165 vss.n16914 vss.n16913 4.65
R16166 vss.n16928 vss.n16927 4.65
R16167 vss.n16942 vss.n16941 4.65
R16168 vss.n16956 vss.n16955 4.65
R16169 vss.n16970 vss.n16969 4.65
R16170 vss.n16984 vss.n16983 4.65
R16171 vss.n16998 vss.n16997 4.65
R16172 vss.n17012 vss.n17011 4.65
R16173 vss.n16863 vss.n16862 4.65
R16174 vss.n17265 vss.n17264 4.65
R16175 vss.n17017 vss.n17016 4.65
R16176 vss.n17029 vss.n17028 4.65
R16177 vss.n17043 vss.n17042 4.65
R16178 vss.n17057 vss.n17056 4.65
R16179 vss.n17071 vss.n17070 4.65
R16180 vss.n17085 vss.n17084 4.65
R16181 vss.n17099 vss.n17098 4.65
R16182 vss.n17113 vss.n17112 4.65
R16183 vss.n17127 vss.n17126 4.65
R16184 vss.n17138 vss.n17137 4.65
R16185 vss.n17150 vss.n17149 4.65
R16186 vss.n17164 vss.n17163 4.65
R16187 vss.n17178 vss.n17177 4.65
R16188 vss.n17192 vss.n17191 4.65
R16189 vss.n17206 vss.n17205 4.65
R16190 vss.n17220 vss.n17219 4.65
R16191 vss.n17234 vss.n17233 4.65
R16192 vss.n17248 vss.n17247 4.65
R16193 vss.n17253 vss.n17252 4.65
R16194 vss.n16265 vss.n16264 4.65
R16195 vss.n16252 vss.n16251 4.65
R16196 vss.n22757 vss.n22756 4.65
R16197 vss.n22755 vss.n22754 4.65
R16198 vss.n22752 vss.n22751 4.65
R16199 vss.n22738 vss.n22737 4.65
R16200 vss.n22724 vss.n22723 4.65
R16201 vss.n22710 vss.n22709 4.65
R16202 vss.n22695 vss.n22694 4.65
R16203 vss.n22690 vss.n22689 4.65
R16204 vss.n22674 vss.n22673 4.65
R16205 vss.n22660 vss.n22659 4.65
R16206 vss.n22646 vss.n22645 4.65
R16207 vss.n22632 vss.n22631 4.65
R16208 vss.n22618 vss.n22617 4.65
R16209 vss.n22604 vss.n22603 4.65
R16210 vss.n22586 vss.n22585 4.65
R16211 vss.n22572 vss.n22571 4.65
R16212 vss.n22558 vss.n22557 4.65
R16213 vss.n22544 vss.n22543 4.65
R16214 vss.n22530 vss.n22529 4.65
R16215 vss.n22516 vss.n22515 4.65
R16216 vss.n22502 vss.n22501 4.65
R16217 vss.n22487 vss.n22486 4.65
R16218 vss.n22482 vss.n22481 4.65
R16219 vss.n22466 vss.n22465 4.65
R16220 vss.n22452 vss.n22451 4.65
R16221 vss.n22438 vss.n22437 4.65
R16222 vss.n22424 vss.n22423 4.65
R16223 vss.n22410 vss.n22409 4.65
R16224 vss.n22396 vss.n22395 4.65
R16225 vss.n22378 vss.n22377 4.65
R16226 vss.n22364 vss.n22363 4.65
R16227 vss.n22350 vss.n22349 4.65
R16228 vss.n22336 vss.n22335 4.65
R16229 vss.n22322 vss.n22321 4.65
R16230 vss.n22308 vss.n22307 4.65
R16231 vss.n22294 vss.n22293 4.65
R16232 vss.n22279 vss.n22278 4.65
R16233 vss.n22274 vss.n22273 4.65
R16234 vss.n22258 vss.n22257 4.65
R16235 vss.n22244 vss.n22243 4.65
R16236 vss.n22230 vss.n22229 4.65
R16237 vss.n22216 vss.n22215 4.65
R16238 vss.n22202 vss.n22201 4.65
R16239 vss.n22188 vss.n22187 4.65
R16240 vss.n22170 vss.n22169 4.65
R16241 vss.n22156 vss.n22155 4.65
R16242 vss.n22142 vss.n22141 4.65
R16243 vss.n22128 vss.n22127 4.65
R16244 vss.n22114 vss.n22113 4.65
R16245 vss.n22100 vss.n22099 4.65
R16246 vss.n226 vss.n225 4.65
R16247 vss.n461 vss.n460 4.65
R16248 vss.n705 vss.n704 4.65
R16249 vss.n949 vss.n948 4.65
R16250 vss.n1194 vss.n1193 4.65
R16251 vss.n23289 vss.n23288 4.65
R16252 vss.n23045 vss.n23044 4.65
R16253 vss.n22828 vss.n22827 4.65
R16254 vss.n22789 vss.n22788 4.65
R16255 vss.n17327 vss.n17326 4.65
R16256 vss.n12288 vss.n12287 4.649
R16257 vss.n10778 vss.n10777 4.649
R16258 vss.n13487 vss.n13486 4.649
R16259 vss.n13181 vss.n13180 4.649
R16260 vss.n12940 vss.n12939 4.649
R16261 vss.n12351 vss.n12350 4.649
R16262 vss.n13775 vss.n13774 4.649
R16263 vss.n13815 vss.n13806 4.649
R16264 vss.n11511 vss.n11510 4.649
R16265 vss.n10566 vss.n10565 4.649
R16266 vss.n12971 vss.n12970 4.649
R16267 vss.n21604 vss.n21603 4.644
R16268 vss.n15311 vss.n15310 4.644
R16269 vss.n16781 vss.n16780 4.643
R16270 vss.n18951 vss.n18950 4.629
R16271 vss.n18949 vss.n17685 4.629
R16272 vss.n17785 vss.n17782 4.629
R16273 vss.n17794 vss.n17792 4.629
R16274 vss.n18709 vss.n17892 4.629
R16275 vss.n18708 vss.n17895 4.629
R16276 vss.n17998 vss.n17995 4.629
R16277 vss.n18007 vss.n18005 4.629
R16278 vss.n18468 vss.n18105 4.629
R16279 vss.n18467 vss.n18108 4.629
R16280 vss.n18211 vss.n18208 4.629
R16281 vss.n18220 vss.n18218 4.629
R16282 vss.n19085 vss.n19082 4.629
R16283 vss.n19094 vss.n19092 4.629
R16284 vss.n20097 vss.n20096 4.629
R16285 vss.n20095 vss.n19192 4.629
R16286 vss.n19292 vss.n19289 4.629
R16287 vss.n19301 vss.n19299 4.629
R16288 vss.n19850 vss.n19849 4.629
R16289 vss.n19848 vss.n19398 4.629
R16290 vss.n19499 vss.n19496 4.629
R16291 vss.n19508 vss.n19506 4.629
R16292 vss.n5561 vss.n5560 4.629
R16293 vss.n5559 vss.n4295 4.629
R16294 vss.n4395 vss.n4392 4.629
R16295 vss.n4404 vss.n4402 4.629
R16296 vss.n5319 vss.n4502 4.629
R16297 vss.n5318 vss.n4505 4.629
R16298 vss.n4608 vss.n4605 4.629
R16299 vss.n4617 vss.n4615 4.629
R16300 vss.n5078 vss.n4715 4.629
R16301 vss.n5077 vss.n4718 4.629
R16302 vss.n4821 vss.n4818 4.629
R16303 vss.n4830 vss.n4828 4.629
R16304 vss.n5695 vss.n5692 4.629
R16305 vss.n5704 vss.n5702 4.629
R16306 vss.n6707 vss.n6706 4.629
R16307 vss.n6705 vss.n5802 4.629
R16308 vss.n5902 vss.n5899 4.629
R16309 vss.n5911 vss.n5909 4.629
R16310 vss.n6460 vss.n6459 4.629
R16311 vss.n6458 vss.n6008 4.629
R16312 vss.n6109 vss.n6106 4.629
R16313 vss.n6118 vss.n6116 4.629
R16314 vss.n11495 vss.n11471 4.619
R16315 vss.n13758 vss.n13679 4.619
R16316 vss.n13152 vss.n13129 4.619
R16317 vss.n13152 vss.n13138 4.619
R16318 vss.n10686 vss.n10666 4.619
R16319 vss.n12695 vss.n12403 4.619
R16320 vss.n10686 vss.n10658 4.619
R16321 vss.n11495 vss.n11463 4.619
R16322 vss.n12036 vss.n12035 4.619
R16323 vss.n11316 vss.n11315 4.619
R16324 vss.n13758 vss.n13647 4.619
R16325 vss.n14077 vss.n13963 4.619
R16326 vss.n11817 vss.n11816 4.619
R16327 vss.n14723 vss.n14713 4.619
R16328 vss.n14587 vss.n14577 4.619
R16329 vss.n15006 vss.n15005 4.619
R16330 vss.n21746 vss.n21708 4.612
R16331 vss.n3695 vss.n3657 4.612
R16332 vss.n12590 vss.n12532 4.588
R16333 vss.n12245 vss.n12063 4.588
R16334 vss.n11495 vss.n11481 4.588
R16335 vss.n13758 vss.n13670 4.588
R16336 vss.n13152 vss.n13121 4.588
R16337 vss.n13152 vss.n13148 4.588
R16338 vss.n12679 vss.n12419 4.588
R16339 vss.n12716 vss.n10527 4.588
R16340 vss.n10686 vss.n10676 4.588
R16341 vss.n12695 vss.n12413 4.588
R16342 vss.n11495 vss.n11491 4.588
R16343 vss.n12334 vss.n12330 4.588
R16344 vss.n12036 vss.n10812 4.588
R16345 vss.n12013 vss.n10818 4.588
R16346 vss.n11951 vss.n10925 4.588
R16347 vss.n11291 vss.n10943 4.588
R16348 vss.n11184 vss.n11034 4.588
R16349 vss.n11316 vss.n10937 4.588
R16350 vss.n13758 vss.n13657 4.588
R16351 vss.n14077 vss.n14066 4.588
R16352 vss.n11817 vss.n11699 4.588
R16353 vss.n14377 vss.n14280 4.588
R16354 vss.n13932 vss.n13845 4.588
R16355 vss.n14044 vss.n13971 4.588
R16356 vss.n11792 vss.n11705 4.588
R16357 vss.n11656 vss.n11565 4.588
R16358 vss.n14727 vss.n13359 4.588
R16359 vss.n14723 vss.n13379 4.588
R16360 vss.n14674 vss.n13507 4.588
R16361 vss.n14587 vss.n14567 4.588
R16362 vss.n14515 vss.n14172 4.588
R16363 vss.n14599 vss.n13597 4.588
R16364 vss.n15008 vss.n12831 4.588
R16365 vss.n14968 vss.n13191 4.588
R16366 vss.n13233 vss.n13232 4.588
R16367 vss.n15006 vss.n14986 4.588
R16368 vss.n15309 vss.n15239 4.587
R16369 vss.n15325 vss.n15227 4.587
R16370 vss.n16779 vss.n16268 4.587
R16371 vss.n16797 vss.n16267 4.587
R16372 vss.n8248 vss.n8243 4.581
R16373 vss.n14995 vss.n14993 4.577
R16374 vss.n11689 vss.n11688 4.577
R16375 vss.n10538 vss.n10537 4.577
R16376 vss.n13151 vss.n13150 4.577
R16377 vss.n13150 vss.n13149 4.577
R16378 vss.n13109 vss.n13108 4.577
R16379 vss.n13108 vss.n13107 4.577
R16380 vss.n10685 vss.n10684 4.577
R16381 vss.n10684 vss.n10683 4.577
R16382 vss.n12333 vss.n12332 4.577
R16383 vss.n12332 vss.n12331 4.577
R16384 vss.n12263 vss.n12262 4.577
R16385 vss.n12262 vss.n12261 4.577
R16386 vss.n14087 vss.n14086 4.577
R16387 vss.n14086 vss.n14085 4.577
R16388 vss.n13660 vss.n13659 4.577
R16389 vss.n13659 vss.n13658 4.577
R16390 vss.n11494 vss.n11493 4.577
R16391 vss.n11493 vss.n11492 4.577
R16392 vss.n11847 vss.n11846 4.577
R16393 vss.n11846 vss.n11845 4.577
R16394 vss.n11939 vss.n11938 4.577
R16395 vss.n11938 vss.n11937 4.577
R16396 vss.n13948 vss.n13944 4.577
R16397 vss.n13949 vss.n13948 4.577
R16398 vss.n11688 vss.n11687 4.577
R16399 vss.n14722 vss.n14721 4.577
R16400 vss.n14721 vss.n14720 4.577
R16401 vss.n14586 vss.n14585 4.577
R16402 vss.n14585 vss.n14584 4.577
R16403 vss.n14496 vss.n14495 4.562
R16404 vss.n13333 vss.n13332 4.562
R16405 vss.n13231 vss.n13230 4.562
R16406 vss.n13190 vss.n13189 4.562
R16407 vss.n12830 vss.n12829 4.562
R16408 vss.n14362 vss.n14361 4.562
R16409 vss.n13857 vss.n13856 4.562
R16410 vss.n11765 vss.n11764 4.562
R16411 vss.n12084 vss.n12083 4.562
R16412 vss.n12531 vss.n12530 4.562
R16413 vss.n10945 vss.n10944 4.562
R16414 vss.n11016 vss.n11015 4.562
R16415 vss.n20654 vss.n17528 4.558
R16416 vss.n12248 vss.n12056 4.558
R16417 vss.n12265 vss.n12046 4.558
R16418 vss.n11219 vss.n10975 4.558
R16419 vss.n11218 vss.n10985 4.558
R16420 vss.n11134 vss.n11120 4.558
R16421 vss.n11133 vss.n11130 4.558
R16422 vss.n13951 vss.n13828 4.558
R16423 vss.n13935 vss.n13838 4.558
R16424 vss.n14724 vss.n13369 4.558
R16425 vss.n14703 vss.n13389 4.558
R16426 vss.n14443 vss.n14201 4.558
R16427 vss.n14442 vss.n14211 4.558
R16428 vss.n7264 vss.n4138 4.558
R16429 vss.n1875 vss.n1650 4.558
R16430 vss.n1876 vss.n1638 4.558
R16431 vss.n2120 vss.n1623 4.558
R16432 vss.n2121 vss.n1611 4.558
R16433 vss.n2364 vss.n1598 4.558
R16434 vss.n2365 vss.n1586 4.558
R16435 vss.n2608 vss.n1573 4.558
R16436 vss.n2610 vss.n1560 4.558
R16437 vss.n2847 vss.n1543 4.558
R16438 vss.n2848 vss.n1528 4.558
R16439 vss.n3091 vss.n1515 4.558
R16440 vss.n3092 vss.n1503 4.558
R16441 vss.n3336 vss.n1488 4.558
R16442 vss.n3337 vss.n1476 4.558
R16443 vss.n336 vss.n111 4.558
R16444 vss.n337 vss.n99 4.558
R16445 vss.n581 vss.n84 4.558
R16446 vss.n582 vss.n72 4.558
R16447 vss.n825 vss.n59 4.558
R16448 vss.n826 vss.n47 4.558
R16449 vss.n1069 vss.n34 4.558
R16450 vss.n1071 vss.n21 4.558
R16451 vss.n23409 vss.n1323 4.558
R16452 vss.n23408 vss.n1335 4.558
R16453 vss.n23166 vss.n1349 4.558
R16454 vss.n23165 vss.n1361 4.558
R16455 vss.n22921 vss.n1376 4.558
R16456 vss.n22920 vss.n1388 4.558
R16457 vss.n12953 vss.n12951 4.557
R16458 vss.n13183 vss.n13164 4.557
R16459 vss.n12994 vss.n12992 4.557
R16460 vss.n12994 vss.n12982 4.557
R16461 vss.n12393 vss.n12365 4.557
R16462 vss.n12393 vss.n12392 4.557
R16463 vss.n10724 vss.n10706 4.557
R16464 vss.n10724 vss.n10696 4.557
R16465 vss.n10792 vss.n10791 4.557
R16466 vss.n13420 vss.n13419 4.557
R16467 vss.n13499 vss.n13498 4.557
R16468 vss.n12300 vss.n12299 4.557
R16469 vss.n13798 vss.n13797 4.557
R16470 vss.n13798 vss.n13786 4.557
R16471 vss.n11554 vss.n11553 4.557
R16472 vss.n11524 vss.n11522 4.557
R16473 vss.n21750 vss.n21705 4.551
R16474 vss.n3699 vss.n3654 4.551
R16475 vss.n12240 vss.n12085 4.527
R16476 vss.n12727 vss.n10510 4.527
R16477 vss.n12007 vss.n10829 4.527
R16478 vss.n11954 vss.n10903 4.527
R16479 vss.n11201 vss.n11017 4.527
R16480 vss.n11274 vss.n10955 4.527
R16481 vss.n14364 vss.n14363 4.527
R16482 vss.n13927 vss.n13867 4.527
R16483 vss.n11653 vss.n11577 4.527
R16484 vss.n11767 vss.n11766 4.527
R16485 vss.n14029 vss.n13982 4.527
R16486 vss.n14732 vss.n13343 4.527
R16487 vss.n14667 vss.n14666 4.527
R16488 vss.n14602 vss.n13584 4.527
R16489 vss.n14498 vss.n14497 4.527
R16490 vss.n15307 vss.n15249 4.526
R16491 vss.n16768 vss.n16767 4.526
R16492 vss.n12661 vss.n12437 4.521
R16493 vss.n14364 vss.n14351 4.521
R16494 vss.n14667 vss.n14655 4.521
R16495 vss.n14498 vss.n14485 4.521
R16496 vss.n20445 vss.n20444 4.517
R16497 vss.n20627 vss.n20626 4.517
R16498 vss.n20675 vss.n20674 4.517
R16499 vss.n20851 vss.n20850 4.517
R16500 vss.n21740 vss.n21714 4.517
R16501 vss.n21648 vss.n21643 4.517
R16502 vss.n12221 vss.n12220 4.517
R16503 vss.n12015 vss.n12014 4.517
R16504 vss.n11251 vss.n11250 4.517
R16505 vss.n11191 vss.n11190 4.517
R16506 vss.n13908 vss.n13907 4.517
R16507 vss.n14046 vss.n14045 4.517
R16508 vss.n11741 vss.n11740 4.517
R16509 vss.n11068 vss.n11067 4.517
R16510 vss.n14735 vss.n14734 4.517
R16511 vss.n14676 vss.n14675 4.517
R16512 vss.n14463 vss.n14462 4.517
R16513 vss.n14245 vss.n14244 4.517
R16514 vss.n12858 vss.n12848 4.517
R16515 vss.n12850 vss.n12849 4.517
R16516 vss.n12658 vss.n12648 4.517
R16517 vss.n12650 vss.n12649 4.517
R16518 vss.n3689 vss.n3663 4.517
R16519 vss.n3597 vss.n3592 4.517
R16520 vss.n7055 vss.n7054 4.517
R16521 vss.n7237 vss.n7236 4.517
R16522 vss.n7285 vss.n7284 4.517
R16523 vss.n7461 vss.n7460 4.517
R16524 vss.n1848 vss.n1847 4.517
R16525 vss.n1897 vss.n1896 4.517
R16526 vss.n2090 vss.n2089 4.517
R16527 vss.n2141 vss.n2140 4.517
R16528 vss.n2335 vss.n2334 4.517
R16529 vss.n2385 vss.n2384 4.517
R16530 vss.n2579 vss.n2578 4.517
R16531 vss.n2630 vss.n2629 4.517
R16532 vss.n2868 vss.n2867 4.517
R16533 vss.n3062 vss.n3061 4.517
R16534 vss.n3113 vss.n3112 4.517
R16535 vss.n3306 vss.n3305 4.517
R16536 vss.n3356 vss.n3355 4.517
R16537 vss.n309 vss.n308 4.517
R16538 vss.n358 vss.n357 4.517
R16539 vss.n551 vss.n550 4.517
R16540 vss.n602 vss.n601 4.517
R16541 vss.n796 vss.n795 4.517
R16542 vss.n846 vss.n845 4.517
R16543 vss.n1040 vss.n1039 4.517
R16544 vss.n1091 vss.n1090 4.517
R16545 vss.n1285 vss.n1284 4.517
R16546 vss.n23379 vss.n23378 4.517
R16547 vss.n23186 vss.n23185 4.517
R16548 vss.n23135 vss.n23134 4.517
R16549 vss.n22942 vss.n22941 4.517
R16550 vss.n22893 vss.n22892 4.517
R16551 vss.n21753 vss.n21705 4.514
R16552 vss.n3702 vss.n3654 4.514
R16553 vss.n21605 vss.n21590 4.513
R16554 vss.n20402 vss.n20401 4.5
R16555 vss.n20400 vss.n17551 4.5
R16556 vss.n20399 vss.n20398 4.5
R16557 vss.n17563 vss.n17558 4.5
R16558 vss.n17562 vss.n17558 4.5
R16559 vss.n20381 vss.n17558 4.5
R16560 vss.n17579 vss.n17576 4.5
R16561 vss.n20380 vss.n20379 4.5
R16562 vss.n20371 vss.n20370 4.5
R16563 vss.n20370 vss.n20369 4.5
R16564 vss.n20362 vss.n17583 4.5
R16565 vss.n17588 vss.n17583 4.5
R16566 vss.n20365 vss.n17580 4.5
R16567 vss.n19614 vss.n19613 4.5
R16568 vss.n19613 vss.n19612 4.5
R16569 vss.n20361 vss.n20360 4.5
R16570 vss.n19617 vss.n19588 4.5
R16571 vss.n19618 vss.n19617 4.5
R16572 vss.n19622 vss.n19621 4.5
R16573 vss.n19621 vss.n19620 4.5
R16574 vss.n20396 vss.n17557 4.5
R16575 vss.n20393 vss.n20392 4.5
R16576 vss.n20375 vss.n17574 4.5
R16577 vss.n17571 vss.n17570 4.5
R16578 vss.n20387 vss.n20386 4.5
R16579 vss.n17570 vss.n17565 4.5
R16580 vss.n17570 vss.n17569 4.5
R16581 vss.n20392 vss.n17560 4.5
R16582 vss.n20392 vss.n20391 4.5
R16583 vss.n17559 vss.n17557 4.5
R16584 vss.n20403 vss.n20402 4.5
R16585 vss.n20404 vss.n17550 4.5
R16586 vss.n21644 vss.n21641 4.5
R16587 vss.n21801 vss.n21641 4.5
R16588 vss.n21757 vss.n21756 4.5
R16589 vss.n21751 vss.n21750 4.5
R16590 vss.n21750 vss.n21749 4.5
R16591 vss.n21800 vss.n21644 4.5
R16592 vss.n21801 vss.n21800 4.5
R16593 vss.n21757 vss.n21755 4.5
R16594 vss.n21757 vss.n21702 4.5
R16595 vss.n21946 vss.n21945 4.5
R16596 vss.n21901 vss.n21900 4.5
R16597 vss.n21892 vss.n21891 4.5
R16598 vss.n21806 vss.n21805 4.5
R16599 vss.n9000 vss.n8984 4.5
R16600 vss.n9030 vss.n9014 4.5
R16601 vss.n9061 vss.n9045 4.5
R16602 vss.n9092 vss.n9076 4.5
R16603 vss.n9112 vss.n9096 4.5
R16604 vss.n14840 vss.n14839 4.5
R16605 vss.n14855 vss.n14854 4.5
R16606 vss.n14911 vss.n14910 4.5
R16607 vss.n14896 vss.n14895 4.5
R16608 vss.n14881 vss.n14880 4.5
R16609 vss.n12844 vss.n12843 4.5
R16610 vss.n12859 vss.n12858 4.5
R16611 vss.n12874 vss.n12873 4.5
R16612 vss.n12895 vss.n12894 4.5
R16613 vss.n12923 vss.n12922 4.5
R16614 vss.n12818 vss.n12817 4.5
R16615 vss.n12775 vss.n12774 4.5
R16616 vss.n15059 vss.n15058 4.5
R16617 vss.n12708 vss.n12707 4.5
R16618 vss.n12692 vss.n12691 4.5
R16619 vss.n12675 vss.n12674 4.5
R16620 vss.n12659 vss.n12658 4.5
R16621 vss.n12510 vss.n12509 4.5
R16622 vss.n12562 vss.n12561 4.5
R16623 vss.n12541 vss.n12540 4.5
R16624 vss.n3593 vss.n3590 4.5
R16625 vss.n3750 vss.n3590 4.5
R16626 vss.n3706 vss.n3705 4.5
R16627 vss.n3700 vss.n3699 4.5
R16628 vss.n3699 vss.n3698 4.5
R16629 vss.n3749 vss.n3593 4.5
R16630 vss.n3750 vss.n3749 4.5
R16631 vss.n3706 vss.n3704 4.5
R16632 vss.n3706 vss.n3651 4.5
R16633 vss.n3895 vss.n3894 4.5
R16634 vss.n3850 vss.n3849 4.5
R16635 vss.n3841 vss.n3840 4.5
R16636 vss.n3755 vss.n3754 4.5
R16637 vss.n7012 vss.n7011 4.5
R16638 vss.n7010 vss.n4161 4.5
R16639 vss.n7009 vss.n7008 4.5
R16640 vss.n4173 vss.n4168 4.5
R16641 vss.n4172 vss.n4168 4.5
R16642 vss.n6991 vss.n4168 4.5
R16643 vss.n4189 vss.n4186 4.5
R16644 vss.n6990 vss.n6989 4.5
R16645 vss.n6981 vss.n6980 4.5
R16646 vss.n6980 vss.n6979 4.5
R16647 vss.n6972 vss.n4193 4.5
R16648 vss.n4198 vss.n4193 4.5
R16649 vss.n6975 vss.n4190 4.5
R16650 vss.n6224 vss.n6223 4.5
R16651 vss.n6223 vss.n6222 4.5
R16652 vss.n6971 vss.n6970 4.5
R16653 vss.n6227 vss.n6198 4.5
R16654 vss.n6228 vss.n6227 4.5
R16655 vss.n6232 vss.n6231 4.5
R16656 vss.n6231 vss.n6230 4.5
R16657 vss.n7006 vss.n4167 4.5
R16658 vss.n7003 vss.n7002 4.5
R16659 vss.n6985 vss.n4184 4.5
R16660 vss.n4181 vss.n4180 4.5
R16661 vss.n6997 vss.n6996 4.5
R16662 vss.n4180 vss.n4175 4.5
R16663 vss.n4180 vss.n4179 4.5
R16664 vss.n7002 vss.n4170 4.5
R16665 vss.n7002 vss.n7001 4.5
R16666 vss.n4169 vss.n4167 4.5
R16667 vss.n7013 vss.n7012 4.5
R16668 vss.n7014 vss.n4160 4.5
R16669 vss.n10536 vss.n10535 4.498
R16670 vss.n14992 vss.n14991 4.498
R16671 vss.n13183 vss.n13165 4.483
R16672 vss.n13013 vss.n12996 4.483
R16673 vss.n13013 vss.n12995 4.483
R16674 vss.n12355 vss.n12353 4.483
R16675 vss.n12355 vss.n12354 4.483
R16676 vss.n10570 vss.n10569 4.483
R16677 vss.n10570 vss.n10568 4.483
R16678 vss.n10792 vss.n10781 4.483
R16679 vss.n13420 vss.n13409 4.483
R16680 vss.n13499 vss.n13469 4.483
R16681 vss.n12300 vss.n12269 4.483
R16682 vss.n13818 vss.n13799 4.483
R16683 vss.n13818 vss.n13817 4.483
R16684 vss.n11554 vss.n11525 4.483
R16685 vss.n16494 vss.n16482 4.48
R16686 vss.n16783 vss.n16782 4.48
R16687 vss.n17016 vss.n17015 4.48
R16688 vss.n17252 vss.n17251 4.48
R16689 vss.n16073 vss.n16061 4.48
R16690 vss.n15322 vss.n15312 4.48
R16691 vss.n15547 vss.n15535 4.48
R16692 vss.n15781 vss.n15771 4.48
R16693 vss.n20764 vss.n17502 4.47
R16694 vss.n20769 vss.n17501 4.47
R16695 vss.n21895 vss.n21861 4.47
R16696 vss.n21820 vss.n21817 4.47
R16697 vss.n11966 vss.n11957 4.47
R16698 vss.n11951 vss.n10926 4.47
R16699 vss.n11656 vss.n11566 4.47
R16700 vss.n11641 vss.n11640 4.47
R16701 vss.n14376 vss.n14281 4.47
R16702 vss.n14411 vss.n14269 4.47
R16703 vss.n14599 vss.n14598 4.47
R16704 vss.n14605 vss.n13565 4.47
R16705 vss.n3844 vss.n3810 4.47
R16706 vss.n3769 vss.n3766 4.47
R16707 vss.n7374 vss.n4112 4.47
R16708 vss.n7379 vss.n4111 4.47
R16709 vss.n1766 vss.n1651 4.47
R16710 vss.n1761 vss.n1652 4.47
R16711 vss.n15190 vss.n3428 4.47
R16712 vss.n15195 vss.n3427 4.47
R16713 vss.n227 vss.n112 4.47
R16714 vss.n222 vss.n113 4.47
R16715 vss.n22824 vss.n1403 4.47
R16716 vss.n22829 vss.n1402 4.47
R16717 vss.n12731 vss.n10480 4.468
R16718 vss.n11994 vss.n10848 4.468
R16719 vss.n11966 vss.n10892 4.468
R16720 vss.n14026 vss.n14003 4.468
R16721 vss.n11641 vss.n11595 4.468
R16722 vss.n14644 vss.n14643 4.468
R16723 vss.n14605 vss.n13564 4.468
R16724 vss.n17317 vss.n17286 4.466
R16725 vss.n11848 vss.n11838 4.453
R16726 vss.n14092 vss.n14080 4.453
R16727 vss.n13110 vss.n13100 4.453
R16728 vss.n13110 vss.n13102 4.453
R16729 vss.n12713 vss.n10540 4.453
R16730 vss.n12334 vss.n12320 4.453
R16731 vss.n10686 vss.n10678 4.453
R16732 vss.n11848 vss.n11840 4.453
R16733 vss.n12264 vss.n12250 4.453
R16734 vss.n11940 vss.n11926 4.453
R16735 vss.n14092 vss.n14091 4.453
R16736 vss.n13950 vss.n13937 4.453
R16737 vss.n11667 vss.n11558 4.453
R16738 vss.n14699 vss.n14688 4.453
R16739 vss.n14532 vss.n14166 4.453
R16740 vss.n14973 vss.n14970 4.453
R16741 vss.n8976 vss.n8975 4.451
R16742 vss.n11848 vss.n11836 4.425
R16743 vss.n14092 vss.n13639 4.425
R16744 vss.n13110 vss.n13015 4.425
R16745 vss.n13110 vss.n13098 4.425
R16746 vss.n12713 vss.n10529 4.425
R16747 vss.n12334 vss.n10729 4.425
R16748 vss.n12334 vss.n10727 4.425
R16749 vss.n11848 vss.n11834 4.425
R16750 vss.n12264 vss.n12252 4.425
R16751 vss.n11940 vss.n11928 4.425
R16752 vss.n14092 vss.n14089 4.425
R16753 vss.n13950 vss.n13939 4.425
R16754 vss.n11667 vss.n11556 4.425
R16755 vss.n14699 vss.n13501 4.425
R16756 vss.n14532 vss.n14531 4.425
R16757 vss.n14973 vss.n14972 4.425
R16758 vss.n21814 vss.n21813 4.387
R16759 vss.n3763 vss.n3762 4.387
R16760 vss.n21670 vss.n21669 4.385
R16761 vss.n3619 vss.n3618 4.385
R16762 vss.n12243 vss.n12073 4.384
R16763 vss.n12036 vss.n10802 4.384
R16764 vss.n11203 vss.n11005 4.384
R16765 vss.n11222 vss.n10965 4.384
R16766 vss.n11723 vss.n11722 4.384
R16767 vss.n14077 vss.n14076 4.384
R16768 vss.n13930 vss.n13855 4.384
R16769 vss.n14729 vss.n13353 4.384
R16770 vss.n14699 vss.n14698 4.384
R16771 vss.n14446 vss.n14191 4.384
R16772 vss.n10182 vss.n10179 4.37
R16773 vss.n11086 vss.n11085 4.327
R16774 vss.n12644 vss.n12457 4.326
R16775 vss.n9110 vss.n9109 4.307
R16776 vss.n20316 vss.n17558 4.302
R16777 vss.n22049 vss.n21984 4.302
R16778 vss.n21614 vss.n21613 4.302
R16779 vss.n11968 vss.n10872 4.302
R16780 vss.n11940 vss.n10927 4.302
R16781 vss.n11667 vss.n11559 4.302
R16782 vss.n11629 vss.n11604 4.302
R16783 vss.n14341 vss.n14282 4.302
R16784 vss.n14607 vss.n13535 4.302
R16785 vss.n14587 vss.n13598 4.302
R16786 vss.n3998 vss.n3933 4.302
R16787 vss.n3563 vss.n3562 4.302
R16788 vss.n6926 vss.n4168 4.302
R16789 vss.n17329 vss.n15210 4.266
R16790 vss.n14263 vss.n14262 4.238
R16791 vss.n12006 vss.n12005 4.201
R16792 vss.n13992 vss.n13991 4.201
R16793 vss.n13517 vss.n13516 4.201
R16794 vss.n21898 vss.n21897 4.191
R16795 vss.n3847 vss.n3846 4.191
R16796 vss.n21860 vss.n21857 4.162
R16797 vss.n3809 vss.n3806 4.162
R16798 vss.n15174 vss.n3477 4.147
R16799 vss.n22808 vss.n1452 4.147
R16800 vss.n20499 vss.n20491 4.141
R16801 vss.n20590 vss.n20582 4.141
R16802 vss.n20728 vss.n20720 4.141
R16803 vss.n20813 vss.n20805 4.141
R16804 vss.n21873 vss.n21869 4.141
R16805 vss.n21782 vss.n21775 4.141
R16806 vss.n12173 vss.n12166 4.141
R16807 vss.n11991 vss.n11984 4.141
R16808 vss.n11325 vss.n11318 4.141
R16809 vss.n14313 vss.n14306 4.141
R16810 vss.n11613 vss.n11606 4.141
R16811 vss.n11826 vss.n11819 4.141
R16812 vss.n14803 vss.n14796 4.141
R16813 vss.n14630 vss.n14623 4.141
R16814 vss.n14541 vss.n14534 4.141
R16815 vss.n14262 vss.n14255 4.141
R16816 vss.n14895 vss.n14894 4.141
R16817 vss.n14894 vss.n14887 4.141
R16818 vss.n15056 vss.n15043 4.141
R16819 vss.n15058 vss.n15056 4.141
R16820 vss.n12707 vss.n12706 4.141
R16821 vss.n12706 vss.n12699 4.141
R16822 vss.n3822 vss.n3818 4.141
R16823 vss.n3731 vss.n3724 4.141
R16824 vss.n7109 vss.n7101 4.141
R16825 vss.n7200 vss.n7192 4.141
R16826 vss.n7338 vss.n7330 4.141
R16827 vss.n7423 vss.n7415 4.141
R16828 vss.n1722 vss.n1714 4.141
R16829 vss.n1811 vss.n1803 4.141
R16830 vss.n1954 vss.n1945 4.141
R16831 vss.n2051 vss.n2042 4.141
R16832 vss.n2199 vss.n2190 4.141
R16833 vss.n2295 vss.n2286 4.141
R16834 vss.n2443 vss.n2434 4.141
R16835 vss.n2540 vss.n2531 4.141
R16836 vss.n2687 vss.n2678 4.141
R16837 vss.n2784 vss.n2775 4.141
R16838 vss.n2926 vss.n2917 4.141
R16839 vss.n3023 vss.n3014 4.141
R16840 vss.n3170 vss.n3161 4.141
R16841 vss.n3267 vss.n3258 4.141
R16842 vss.n3409 vss.n3401 4.141
R16843 vss.n3476 vss.n3468 4.141
R16844 vss.n183 vss.n175 4.141
R16845 vss.n272 vss.n264 4.141
R16846 vss.n415 vss.n406 4.141
R16847 vss.n512 vss.n503 4.141
R16848 vss.n660 vss.n651 4.141
R16849 vss.n756 vss.n747 4.141
R16850 vss.n904 vss.n895 4.141
R16851 vss.n1001 vss.n992 4.141
R16852 vss.n1148 vss.n1139 4.141
R16853 vss.n1245 vss.n1236 4.141
R16854 vss.n23340 vss.n23331 4.141
R16855 vss.n23243 vss.n23234 4.141
R16856 vss.n23096 vss.n23087 4.141
R16857 vss.n22999 vss.n22990 4.141
R16858 vss.n22856 vss.n22848 4.141
R16859 vss.n1451 vss.n1443 4.141
R16860 vss.n8925 vss.n8924 4.101
R16861 vss.n15156 vss.n3489 4.073
R16862 vss.n22790 vss.n1464 4.073
R16863 vss.n10770 vss.n10768 4.034
R16864 vss.n13397 vss.n13396 4.034
R16865 vss.n13173 vss.n13171 4.034
R16866 vss.n10721 vss.n10712 4.034
R16867 vss.n10560 vss.n10559 4.034
R16868 vss.n13011 vss.n13002 4.034
R16869 vss.n12380 vss.n12371 4.034
R16870 vss.n12345 vss.n12344 4.034
R16871 vss.n13769 vss.n13768 4.034
R16872 vss.n13814 vss.n13812 4.034
R16873 vss.n11540 vss.n11531 4.034
R16874 vss.n11505 vss.n11504 4.034
R16875 vss.n20413 vss.n20412 4.023
R16876 vss.n7023 vss.n7022 4.023
R16877 vss.n11994 vss.n10858 4.003
R16878 vss.n14026 vss.n14013 4.003
R16879 vss.n14644 vss.n13534 4.003
R16880 vss.n10770 vss.n10769 4.001
R16881 vss.n12932 vss.n12931 4.001
R16882 vss.n12963 vss.n12962 4.001
R16883 vss.n9672 vss.n9668 4
R16884 vss.n8927 vss.n8926 3.974
R16885 vss.n19020 vss.n17633 3.94
R16886 vss.n19008 vss.n17637 3.94
R16887 vss.n18893 vss.n17728 3.94
R16888 vss.n18884 vss.n17740 3.94
R16889 vss.n18773 vss.n17838 3.94
R16890 vss.n18763 vss.n17846 3.94
R16891 vss.n18652 vss.n17941 3.94
R16892 vss.n18643 vss.n17953 3.94
R16893 vss.n18532 vss.n18051 3.94
R16894 vss.n18522 vss.n18059 3.94
R16895 vss.n18411 vss.n18154 3.94
R16896 vss.n18402 vss.n18166 3.94
R16897 vss.n18291 vss.n18264 3.94
R16898 vss.n18281 vss.n18272 3.94
R16899 vss.n20285 vss.n17620 3.94
R16900 vss.n20277 vss.n19039 3.94
R16901 vss.n20166 vss.n19138 3.94
R16902 vss.n20154 vss.n19144 3.94
R16903 vss.n20039 vss.n19235 3.94
R16904 vss.n20030 vss.n19247 3.94
R16905 vss.n19919 vss.n19345 3.94
R16906 vss.n19907 vss.n19351 3.94
R16907 vss.n19792 vss.n19442 3.94
R16908 vss.n19783 vss.n19454 3.94
R16909 vss.n19672 vss.n19552 3.94
R16910 vss.n19660 vss.n19558 3.94
R16911 vss.n17611 vss.n17607 3.94
R16912 vss.n20302 vss.n20301 3.94
R16913 vss.n5630 vss.n4243 3.94
R16914 vss.n5618 vss.n4247 3.94
R16915 vss.n5503 vss.n4338 3.94
R16916 vss.n5494 vss.n4350 3.94
R16917 vss.n5383 vss.n4448 3.94
R16918 vss.n5373 vss.n4456 3.94
R16919 vss.n5262 vss.n4551 3.94
R16920 vss.n5253 vss.n4563 3.94
R16921 vss.n5142 vss.n4661 3.94
R16922 vss.n5132 vss.n4669 3.94
R16923 vss.n5021 vss.n4764 3.94
R16924 vss.n5012 vss.n4776 3.94
R16925 vss.n4901 vss.n4874 3.94
R16926 vss.n4891 vss.n4882 3.94
R16927 vss.n6895 vss.n4230 3.94
R16928 vss.n6887 vss.n5649 3.94
R16929 vss.n6776 vss.n5748 3.94
R16930 vss.n6764 vss.n5754 3.94
R16931 vss.n6649 vss.n5845 3.94
R16932 vss.n6640 vss.n5857 3.94
R16933 vss.n6529 vss.n5955 3.94
R16934 vss.n6517 vss.n5961 3.94
R16935 vss.n6402 vss.n6052 3.94
R16936 vss.n6393 vss.n6064 3.94
R16937 vss.n6282 vss.n6162 3.94
R16938 vss.n6270 vss.n6168 3.94
R16939 vss.n4221 vss.n4217 3.94
R16940 vss.n6912 vss.n6911 3.94
R16941 vss.n16682 vss.n16679 3.94
R16942 vss.n16887 vss.n16883 3.94
R16943 vss.n16910 vss.n16906 3.94
R16944 vss.n17123 vss.n17119 3.94
R16945 vss.n17146 vss.n17142 3.94
R16946 vss.n16263 vss.n16260 3.94
R16947 vss.n15933 vss.n15929 3.94
R16948 vss.n15957 vss.n15953 3.94
R16949 vss.n16169 vss.n16165 3.94
R16950 vss.n16193 vss.n16189 3.94
R16951 vss.n16291 vss.n16288 3.94
R16952 vss.n15409 vss.n15405 3.94
R16953 vss.n15430 vss.n15426 3.94
R16954 vss.n15645 vss.n15641 3.94
R16955 vss.n15666 vss.n15662 3.94
R16956 vss.n15871 vss.n15868 3.94
R16957 vss.n16356 vss.n16352 3.94
R16958 vss.n16377 vss.n16373 3.94
R16959 vss.n16592 vss.n16588 3.94
R16960 vss.n16613 vss.n16609 3.94
R16961 vss.n10301 vss.n10299 3.917
R16962 vss.n12416 vss.n12415 3.9
R16963 vss.n12528 vss.n12524 3.9
R16964 vss.n13119 vss.n13115 3.9
R16965 vss.n13668 vss.n13664 3.9
R16966 vss.n14169 vss.n14168 3.9
R16967 vss.n13504 vss.n13503 3.9
R16968 vss.n13595 vss.n13594 3.9
R16969 vss.n12827 vss.n12826 3.9
R16970 vss.n13356 vss.n13355 3.9
R16971 vss.n13228 vss.n13224 3.9
R16972 vss.n14984 vss.n14980 3.9
R16973 vss.n13146 vss.n13142 3.9
R16974 vss.n14277 vss.n14273 3.9
R16975 vss.n13655 vss.n13651 3.9
R16976 vss.n14064 vss.n14060 3.9
R16977 vss.n11563 vss.n11562 3.9
R16978 vss.n11479 vss.n11475 3.9
R16979 vss.n11697 vss.n11693 3.9
R16980 vss.n11702 vss.n11701 3.9
R16981 vss.n11042 vss.n11038 3.9
R16982 vss.n10815 vss.n10814 3.9
R16983 vss.n10940 vss.n10939 3.9
R16984 vss.n14565 vss.n14561 3.9
R16985 vss.n14102 vss.n14098 3.9
R16986 vss.n13752 vss.n13748 3.9
R16987 vss.n11449 vss.n11445 3.9
R16988 vss.n11858 vss.n11854 3.9
R16989 vss.n10935 vss.n10931 3.9
R16990 vss.n12411 vss.n12407 3.9
R16991 vss.n10674 vss.n10670 3.9
R16992 vss.n12328 vss.n12324 3.9
R16993 vss.n11489 vss.n11485 3.9
R16994 vss.n13377 vss.n13373 3.9
R16995 vss.n13460 vss.n13456 3.9
R16996 vss.n13091 vss.n13087 3.9
R16997 vss.n10644 vss.n10640 3.9
R16998 vss.n12313 vss.n12309 3.9
R16999 vss.n10810 vss.n10806 3.9
R17000 vss.n12007 vss.n12006 3.868
R17001 vss.n14029 vss.n13992 3.868
R17002 vss.n14667 vss.n13517 3.868
R17003 vss.n22702 vss.n22699 3.862
R17004 vss.n22685 vss.n22682 3.862
R17005 vss.n22494 vss.n22491 3.862
R17006 vss.n22477 vss.n22474 3.862
R17007 vss.n22286 vss.n22283 3.862
R17008 vss.n22269 vss.n22266 3.862
R17009 vss.n22076 vss.n22073 3.862
R17010 vss.n21599 vss.n21596 3.862
R17011 vss.n21422 vss.n21419 3.862
R17012 vss.n21405 vss.n21402 3.862
R17013 vss.n21214 vss.n21211 3.862
R17014 vss.n21197 vss.n21194 3.862
R17015 vss.n21006 vss.n21003 3.862
R17016 vss.n20989 vss.n20986 3.862
R17017 vss.n8865 vss.n8862 3.862
R17018 vss.n8848 vss.n8845 3.862
R17019 vss.n8657 vss.n8654 3.862
R17020 vss.n8640 vss.n8637 3.862
R17021 vss.n8449 vss.n8446 3.862
R17022 vss.n8432 vss.n8429 3.862
R17023 vss.n8236 vss.n8233 3.862
R17024 vss.n8225 vss.n8222 3.862
R17025 vss.n8033 vss.n8030 3.862
R17026 vss.n8016 vss.n8013 3.862
R17027 vss.n7824 vss.n7821 3.862
R17028 vss.n7807 vss.n7804 3.862
R17029 vss.n7616 vss.n7613 3.862
R17030 vss.n7599 vss.n7596 3.862
R17031 vss.n12488 vss.n12487 3.852
R17032 vss.n12821 vss.n12820 3.852
R17033 vss.n10450 vss.n10449 3.846
R17034 vss.n14389 vss.n14387 3.814
R17035 vss.n10524 vss.n10523 3.814
R17036 vss.n13287 vss.n13285 3.814
R17037 vss.n13186 vss.n13185 3.814
R17038 vss.n13841 vss.n13840 3.814
R17039 vss.n13967 vss.n13966 3.814
R17040 vss.n10921 vss.n10920 3.814
R17041 vss.n11030 vss.n11029 3.814
R17042 vss.n12566 vss.n12565 3.814
R17043 vss.n12059 vss.n12058 3.814
R17044 vss.n20307 vss.n20303 3.772
R17045 vss.n6917 vss.n6913 3.772
R17046 vss.n8964 vss.n8962 3.772
R17047 vss.n20461 vss.n20460 3.764
R17048 vss.n20612 vss.n20611 3.764
R17049 vss.n20690 vss.n20689 3.764
R17050 vss.n20835 vss.n20834 3.764
R17051 vss.n21746 vss.n21745 3.764
R17052 vss.n21694 vss.n21686 3.764
R17053 vss.n21797 vss.n21646 3.764
R17054 vss.n21655 vss.n21654 3.764
R17055 vss.n12546 vss.n12545 3.764
R17056 vss.n12561 vss.n12560 3.764
R17057 vss.n12194 vss.n12193 3.764
R17058 vss.n11998 vss.n11997 3.764
R17059 vss.n11277 vss.n11276 3.764
R17060 vss.n11175 vss.n11174 3.764
R17061 vss.n13874 vss.n13873 3.764
R17062 vss.n13984 vss.n13983 3.764
R17063 vss.n11778 vss.n11777 3.764
R17064 vss.n11088 vss.n11087 3.764
R17065 vss.n14768 vss.n14767 3.764
R17066 vss.n13509 vss.n13508 3.764
R17067 vss.n14501 vss.n14500 3.764
R17068 vss.n14215 vss.n14214 3.764
R17069 vss.n12843 vss.n12833 3.764
R17070 vss.n12835 vss.n12834 3.764
R17071 vss.n12802 vss.n12801 3.764
R17072 vss.n12817 vss.n12816 3.764
R17073 vss.n12674 vss.n12664 3.764
R17074 vss.n12666 vss.n12665 3.764
R17075 vss.n3695 vss.n3694 3.764
R17076 vss.n3643 vss.n3635 3.764
R17077 vss.n3746 vss.n3595 3.764
R17078 vss.n3604 vss.n3603 3.764
R17079 vss.n7071 vss.n7070 3.764
R17080 vss.n7222 vss.n7221 3.764
R17081 vss.n7300 vss.n7299 3.764
R17082 vss.n7445 vss.n7444 3.764
R17083 vss.n1684 vss.n1683 3.764
R17084 vss.n1833 vss.n1832 3.764
R17085 vss.n1913 vss.n1912 3.764
R17086 vss.n2074 vss.n2073 3.764
R17087 vss.n2157 vss.n2156 3.764
R17088 vss.n2319 vss.n2318 3.764
R17089 vss.n2402 vss.n2401 3.764
R17090 vss.n2563 vss.n2562 3.764
R17091 vss.n2646 vss.n2645 3.764
R17092 vss.n2807 vss.n2806 3.764
R17093 vss.n2884 vss.n2883 3.764
R17094 vss.n3046 vss.n3045 3.764
R17095 vss.n3129 vss.n3128 3.764
R17096 vss.n3290 vss.n3289 3.764
R17097 vss.n3371 vss.n3370 3.764
R17098 vss.n3480 vss.n3479 3.764
R17099 vss.n145 vss.n144 3.764
R17100 vss.n294 vss.n293 3.764
R17101 vss.n374 vss.n373 3.764
R17102 vss.n535 vss.n534 3.764
R17103 vss.n618 vss.n617 3.764
R17104 vss.n780 vss.n779 3.764
R17105 vss.n863 vss.n862 3.764
R17106 vss.n1024 vss.n1023 3.764
R17107 vss.n1107 vss.n1106 3.764
R17108 vss.n1268 vss.n1267 3.764
R17109 vss.n23363 vss.n23362 3.764
R17110 vss.n23202 vss.n23201 3.764
R17111 vss.n23119 vss.n23118 3.764
R17112 vss.n22958 vss.n22957 3.764
R17113 vss.n22878 vss.n22877 3.764
R17114 vss.n1455 vss.n1454 3.764
R17115 vss.n13698 vss.n13697 3.681
R17116 vss.t328 vss.n9162 3.56
R17117 vss.n21671 vss.n21670 3.544
R17118 vss.n3620 vss.n3619 3.544
R17119 vss.n3455 vss.n3454 3.53
R17120 vss.n1430 vss.n1429 3.53
R17121 vss.n19024 vss.n17629 3.419
R17122 vss.n5634 vss.n4239 3.419
R17123 vss.n20484 vss.n20476 3.388
R17124 vss.n20605 vss.n20597 3.388
R17125 vss.n20713 vss.n20705 3.388
R17126 vss.n20828 vss.n20820 3.388
R17127 vss.n21884 vss.n21880 3.388
R17128 vss.n21899 vss.n21898 3.388
R17129 vss.n21779 vss.n21778 3.388
R17130 vss.n12187 vss.n12180 3.388
R17131 vss.n10857 vss.n10850 3.388
R17132 vss.n11300 vss.n11293 3.388
R17133 vss.n11161 vss.n11154 3.388
R17134 vss.n14299 vss.n14292 3.388
R17135 vss.n14012 vss.n14005 3.388
R17136 vss.n11801 vss.n11794 3.388
R17137 vss.n11085 vss.n11078 3.388
R17138 vss.n14789 vss.n14782 3.388
R17139 vss.n13533 vss.n13526 3.388
R17140 vss.n14524 vss.n14517 3.388
R17141 vss.n14242 vss.n14235 3.388
R17142 vss.n14880 vss.n14879 3.388
R17143 vss.n14879 vss.n14872 3.388
R17144 vss.n12691 vss.n12690 3.388
R17145 vss.n12690 vss.n12683 3.388
R17146 vss.n3833 vss.n3829 3.388
R17147 vss.n3848 vss.n3847 3.388
R17148 vss.n3728 vss.n3727 3.388
R17149 vss.n7094 vss.n7086 3.388
R17150 vss.n7215 vss.n7207 3.388
R17151 vss.n7323 vss.n7315 3.388
R17152 vss.n7438 vss.n7430 3.388
R17153 vss.n1707 vss.n1699 3.388
R17154 vss.n1826 vss.n1818 3.388
R17155 vss.n1938 vss.n1929 3.388
R17156 vss.n2067 vss.n2058 3.388
R17157 vss.n2182 vss.n2173 3.388
R17158 vss.n2312 vss.n2303 3.388
R17159 vss.n2427 vss.n2418 3.388
R17160 vss.n2556 vss.n2547 3.388
R17161 vss.n2671 vss.n2662 3.388
R17162 vss.n2800 vss.n2791 3.388
R17163 vss.n2909 vss.n2900 3.388
R17164 vss.n3039 vss.n3030 3.388
R17165 vss.n3154 vss.n3145 3.388
R17166 vss.n3283 vss.n3274 3.388
R17167 vss.n3394 vss.n3386 3.388
R17168 vss.n15167 vss.n15159 3.388
R17169 vss.n168 vss.n160 3.388
R17170 vss.n287 vss.n279 3.388
R17171 vss.n399 vss.n390 3.388
R17172 vss.n528 vss.n519 3.388
R17173 vss.n643 vss.n634 3.388
R17174 vss.n773 vss.n764 3.388
R17175 vss.n888 vss.n879 3.388
R17176 vss.n1017 vss.n1008 3.388
R17177 vss.n1132 vss.n1123 3.388
R17178 vss.n1261 vss.n1252 3.388
R17179 vss.n23356 vss.n23347 3.388
R17180 vss.n23227 vss.n23218 3.388
R17181 vss.n23112 vss.n23103 3.388
R17182 vss.n22983 vss.n22974 3.388
R17183 vss.n22871 vss.n22863 3.388
R17184 vss.n22801 vss.n22793 3.388
R17185 vss.n14038 vss.n14030 3.377
R17186 vss.n11775 vss.n11768 3.377
R17187 vss.n10750 vss.n10749 3.377
R17188 vss.n13036 vss.n13035 3.377
R17189 vss.n11361 vss.n11360 3.377
R17190 vss.n13703 vss.n13702 3.377
R17191 vss.n19031 vss.n19030 3.364
R17192 vss.n19032 vss.n17618 3.364
R17193 vss.n5641 vss.n5640 3.364
R17194 vss.n5642 vss.n4228 3.364
R17195 vss.n11776 vss.n11775 3.335
R17196 vss.n14039 vss.n14038 3.335
R17197 vss.n14349 vss.n14348 3.333
R17198 vss.n14482 vss.n14481 3.333
R17199 vss.n11773 vss.n11772 3.333
R17200 vss.n11350 vss.n11349 3.333
R17201 vss.n11358 vss.n11357 3.333
R17202 vss.n10759 vss.n10757 3.333
R17203 vss.n10747 vss.n10746 3.333
R17204 vss.n12435 vss.n12434 3.333
R17205 vss.n13033 vss.n13032 3.333
R17206 vss.n12796 vss.n12794 3.333
R17207 vss.n13571 vss.n13570 3.333
R17208 vss.n14652 vss.n14651 3.333
R17209 vss.n13045 vss.n13043 3.333
R17210 vss.n13710 vss.n13709 3.333
R17211 vss.n13698 vss.n13696 3.333
R17212 vss.n21993 vss.n21992 3.306
R17213 vss.n21992 vss.t141 3.306
R17214 vss.n21996 vss.t357 3.306
R17215 vss.n21996 vss.n21993 3.306
R17216 vss.n21789 vss.n21691 3.306
R17217 vss.n21789 vss.n21647 3.306
R17218 vss.n21796 vss.n21647 3.306
R17219 vss.n21796 vss.t323 3.306
R17220 vss.n21618 vss.t322 3.306
R17221 vss.n21618 vss.t358 3.306
R17222 vss.n3942 vss.n3941 3.306
R17223 vss.n3941 vss.t150 3.306
R17224 vss.n3945 vss.t4 3.306
R17225 vss.n3945 vss.n3942 3.306
R17226 vss.n3738 vss.n3640 3.306
R17227 vss.n3738 vss.n3596 3.306
R17228 vss.n3745 vss.n3596 3.306
R17229 vss.n3745 vss.t6 3.306
R17230 vss.n3567 vss.t7 3.306
R17231 vss.n3567 vss.t5 3.306
R17232 vss.n17526 vss.n17520 3.293
R17233 vss.n17513 vss.n17508 3.293
R17234 vss.n4136 vss.n4130 3.293
R17235 vss.n4123 vss.n4118 3.293
R17236 vss.n1648 vss.n1642 3.293
R17237 vss.n1636 vss.n1630 3.293
R17238 vss.n1621 vss.n1615 3.293
R17239 vss.n1609 vss.n1603 3.293
R17240 vss.n1596 vss.n1590 3.293
R17241 vss.n1584 vss.n1578 3.293
R17242 vss.n1571 vss.n1565 3.293
R17243 vss.n1558 vss.n1552 3.293
R17244 vss.n1541 vss.n1532 3.293
R17245 vss.n1526 vss.n1520 3.293
R17246 vss.n1513 vss.n1507 3.293
R17247 vss.n1501 vss.n1495 3.293
R17248 vss.n1486 vss.n1480 3.293
R17249 vss.n1474 vss.n1468 3.293
R17250 vss.n109 vss.n103 3.293
R17251 vss.n97 vss.n91 3.293
R17252 vss.n82 vss.n76 3.293
R17253 vss.n70 vss.n64 3.293
R17254 vss.n57 vss.n51 3.293
R17255 vss.n45 vss.n39 3.293
R17256 vss.n32 vss.n26 3.293
R17257 vss.n19 vss.n13 3.293
R17258 vss.n1321 vss.n1315 3.293
R17259 vss.n1333 vss.n1327 3.293
R17260 vss.n1347 vss.n1341 3.293
R17261 vss.n1359 vss.n1353 3.293
R17262 vss.n1374 vss.n1368 3.293
R17263 vss.n1386 vss.n1380 3.293
R17264 vss.n12240 vss.n12239 3.27
R17265 vss.n11954 vss.n10918 3.27
R17266 vss.n12007 vss.n10837 3.269
R17267 vss.n11201 vss.n11026 3.269
R17268 vss.n11274 vss.n11273 3.269
R17269 vss.n13109 vss.n13105 3.231
R17270 vss.n10685 vss.n10681 3.231
R17271 vss.n14087 vss.n14083 3.231
R17272 vss.n11847 vss.n11843 3.231
R17273 vss.n14732 vss.n13331 3.217
R17274 vss.n14602 vss.n13573 3.217
R17275 vss.n19026 vss.n19025 3.2
R17276 vss.n19003 vss.n19002 3.2
R17277 vss.n18995 vss.n17646 3.2
R17278 vss.n17658 vss.n17655 3.2
R17279 vss.n18982 vss.n18981 3.2
R17280 vss.n17667 vss.n17665 3.2
R17281 vss.n17677 vss.n17675 3.2
R17282 vss.n18959 vss.n18958 3.2
R17283 vss.n18941 vss.n18940 3.2
R17284 vss.n18935 vss.n17693 3.2
R17285 vss.n18927 vss.n18926 3.2
R17286 vss.n17710 vss.n17706 3.2
R17287 vss.n18912 vss.n17715 3.2
R17288 vss.n18904 vss.n18903 3.2
R17289 vss.n17729 vss.n17725 3.2
R17290 vss.n17747 vss.n17741 3.2
R17291 vss.n17755 vss.n17753 3.2
R17292 vss.n18866 vss.n18865 3.2
R17293 vss.n17764 vss.n17762 3.2
R17294 vss.n17774 vss.n17772 3.2
R17295 vss.n18843 vss.n18842 3.2
R17296 vss.n17783 vss.n17781 3.2
R17297 vss.n18822 vss.n17796 3.2
R17298 vss.n18814 vss.n18813 3.2
R17299 vss.n17810 vss.n17806 3.2
R17300 vss.n18799 vss.n17815 3.2
R17301 vss.n18791 vss.n18790 3.2
R17302 vss.n17829 vss.n17825 3.2
R17303 vss.n18776 vss.n17834 3.2
R17304 vss.n17855 vss.n17853 3.2
R17305 vss.n18753 vss.n18752 3.2
R17306 vss.n17864 vss.n17862 3.2
R17307 vss.n17874 vss.n17872 3.2
R17308 vss.n18730 vss.n18729 3.2
R17309 vss.n17883 vss.n17881 3.2
R17310 vss.n17893 vss.n17891 3.2
R17311 vss.n18700 vss.n18699 3.2
R17312 vss.n18694 vss.n17906 3.2
R17313 vss.n18686 vss.n18685 3.2
R17314 vss.n17923 vss.n17919 3.2
R17315 vss.n18671 vss.n17928 3.2
R17316 vss.n18663 vss.n18662 3.2
R17317 vss.n17942 vss.n17938 3.2
R17318 vss.n17960 vss.n17954 3.2
R17319 vss.n17968 vss.n17966 3.2
R17320 vss.n18625 vss.n18624 3.2
R17321 vss.n17977 vss.n17975 3.2
R17322 vss.n17987 vss.n17985 3.2
R17323 vss.n18602 vss.n18601 3.2
R17324 vss.n17996 vss.n17994 3.2
R17325 vss.n18581 vss.n18009 3.2
R17326 vss.n18573 vss.n18572 3.2
R17327 vss.n18023 vss.n18019 3.2
R17328 vss.n18558 vss.n18028 3.2
R17329 vss.n18550 vss.n18549 3.2
R17330 vss.n18042 vss.n18038 3.2
R17331 vss.n18535 vss.n18047 3.2
R17332 vss.n18068 vss.n18066 3.2
R17333 vss.n18512 vss.n18511 3.2
R17334 vss.n18077 vss.n18075 3.2
R17335 vss.n18087 vss.n18085 3.2
R17336 vss.n18489 vss.n18488 3.2
R17337 vss.n18096 vss.n18094 3.2
R17338 vss.n18106 vss.n18104 3.2
R17339 vss.n18459 vss.n18458 3.2
R17340 vss.n18453 vss.n18119 3.2
R17341 vss.n18445 vss.n18444 3.2
R17342 vss.n18136 vss.n18132 3.2
R17343 vss.n18430 vss.n18141 3.2
R17344 vss.n18422 vss.n18421 3.2
R17345 vss.n18155 vss.n18151 3.2
R17346 vss.n18173 vss.n18167 3.2
R17347 vss.n18181 vss.n18179 3.2
R17348 vss.n18384 vss.n18383 3.2
R17349 vss.n18190 vss.n18188 3.2
R17350 vss.n18200 vss.n18198 3.2
R17351 vss.n18361 vss.n18360 3.2
R17352 vss.n18209 vss.n18207 3.2
R17353 vss.n18340 vss.n18222 3.2
R17354 vss.n18332 vss.n18331 3.2
R17355 vss.n18236 vss.n18232 3.2
R17356 vss.n18317 vss.n18241 3.2
R17357 vss.n18309 vss.n18308 3.2
R17358 vss.n18255 vss.n18251 3.2
R17359 vss.n18294 vss.n18260 3.2
R17360 vss.n18274 vss.n18273 3.2
R17361 vss.n20292 vss.n20291 3.2
R17362 vss.n20272 vss.n19042 3.2
R17363 vss.n19055 vss.n19052 3.2
R17364 vss.n20259 vss.n20258 3.2
R17365 vss.n19064 vss.n19062 3.2
R17366 vss.n19074 vss.n19072 3.2
R17367 vss.n20236 vss.n20235 3.2
R17368 vss.n19083 vss.n19081 3.2
R17369 vss.n20215 vss.n19096 3.2
R17370 vss.n20207 vss.n20206 3.2
R17371 vss.n19110 vss.n19106 3.2
R17372 vss.n20192 vss.n19115 3.2
R17373 vss.n20184 vss.n20183 3.2
R17374 vss.n19129 vss.n19125 3.2
R17375 vss.n20169 vss.n19134 3.2
R17376 vss.n20149 vss.n20148 3.2
R17377 vss.n20141 vss.n19153 3.2
R17378 vss.n19165 vss.n19162 3.2
R17379 vss.n20128 vss.n20127 3.2
R17380 vss.n19174 vss.n19172 3.2
R17381 vss.n19184 vss.n19182 3.2
R17382 vss.n20105 vss.n20104 3.2
R17383 vss.n20087 vss.n20086 3.2
R17384 vss.n20081 vss.n19200 3.2
R17385 vss.n20073 vss.n20072 3.2
R17386 vss.n19217 vss.n19213 3.2
R17387 vss.n20058 vss.n19222 3.2
R17388 vss.n20050 vss.n20049 3.2
R17389 vss.n19236 vss.n19232 3.2
R17390 vss.n19254 vss.n19248 3.2
R17391 vss.n19262 vss.n19260 3.2
R17392 vss.n20012 vss.n20011 3.2
R17393 vss.n19271 vss.n19269 3.2
R17394 vss.n19281 vss.n19279 3.2
R17395 vss.n19989 vss.n19988 3.2
R17396 vss.n19290 vss.n19288 3.2
R17397 vss.n19968 vss.n19303 3.2
R17398 vss.n19960 vss.n19959 3.2
R17399 vss.n19317 vss.n19313 3.2
R17400 vss.n19945 vss.n19322 3.2
R17401 vss.n19937 vss.n19936 3.2
R17402 vss.n19336 vss.n19332 3.2
R17403 vss.n19922 vss.n19341 3.2
R17404 vss.n19902 vss.n19901 3.2
R17405 vss.n19894 vss.n19360 3.2
R17406 vss.n19372 vss.n19369 3.2
R17407 vss.n19881 vss.n19880 3.2
R17408 vss.n19381 vss.n19379 3.2
R17409 vss.n19391 vss.n19389 3.2
R17410 vss.n19858 vss.n19857 3.2
R17411 vss.n19840 vss.n19839 3.2
R17412 vss.n19834 vss.n19407 3.2
R17413 vss.n19826 vss.n19825 3.2
R17414 vss.n19424 vss.n19420 3.2
R17415 vss.n19811 vss.n19429 3.2
R17416 vss.n19803 vss.n19802 3.2
R17417 vss.n19443 vss.n19439 3.2
R17418 vss.n19461 vss.n19455 3.2
R17419 vss.n19469 vss.n19467 3.2
R17420 vss.n19765 vss.n19764 3.2
R17421 vss.n19478 vss.n19476 3.2
R17422 vss.n19488 vss.n19486 3.2
R17423 vss.n19742 vss.n19741 3.2
R17424 vss.n19497 vss.n19495 3.2
R17425 vss.n19721 vss.n19510 3.2
R17426 vss.n19713 vss.n19712 3.2
R17427 vss.n19524 vss.n19520 3.2
R17428 vss.n19698 vss.n19529 3.2
R17429 vss.n19690 vss.n19689 3.2
R17430 vss.n19543 vss.n19539 3.2
R17431 vss.n19675 vss.n19548 3.2
R17432 vss.n19655 vss.n19654 3.2
R17433 vss.n19647 vss.n19567 3.2
R17434 vss.n19579 vss.n19576 3.2
R17435 vss.n19634 vss.n19633 3.2
R17436 vss.n19597 vss.n19586 3.2
R17437 vss.n5636 vss.n5635 3.2
R17438 vss.n5613 vss.n5612 3.2
R17439 vss.n5605 vss.n4256 3.2
R17440 vss.n4268 vss.n4265 3.2
R17441 vss.n5592 vss.n5591 3.2
R17442 vss.n4277 vss.n4275 3.2
R17443 vss.n4287 vss.n4285 3.2
R17444 vss.n5569 vss.n5568 3.2
R17445 vss.n5551 vss.n5550 3.2
R17446 vss.n5545 vss.n4303 3.2
R17447 vss.n5537 vss.n5536 3.2
R17448 vss.n4320 vss.n4316 3.2
R17449 vss.n5522 vss.n4325 3.2
R17450 vss.n5514 vss.n5513 3.2
R17451 vss.n4339 vss.n4335 3.2
R17452 vss.n4357 vss.n4351 3.2
R17453 vss.n4365 vss.n4363 3.2
R17454 vss.n5476 vss.n5475 3.2
R17455 vss.n4374 vss.n4372 3.2
R17456 vss.n4384 vss.n4382 3.2
R17457 vss.n5453 vss.n5452 3.2
R17458 vss.n4393 vss.n4391 3.2
R17459 vss.n5432 vss.n4406 3.2
R17460 vss.n5424 vss.n5423 3.2
R17461 vss.n4420 vss.n4416 3.2
R17462 vss.n5409 vss.n4425 3.2
R17463 vss.n5401 vss.n5400 3.2
R17464 vss.n4439 vss.n4435 3.2
R17465 vss.n5386 vss.n4444 3.2
R17466 vss.n4465 vss.n4463 3.2
R17467 vss.n5363 vss.n5362 3.2
R17468 vss.n4474 vss.n4472 3.2
R17469 vss.n4484 vss.n4482 3.2
R17470 vss.n5340 vss.n5339 3.2
R17471 vss.n4493 vss.n4491 3.2
R17472 vss.n4503 vss.n4501 3.2
R17473 vss.n5310 vss.n5309 3.2
R17474 vss.n5304 vss.n4516 3.2
R17475 vss.n5296 vss.n5295 3.2
R17476 vss.n4533 vss.n4529 3.2
R17477 vss.n5281 vss.n4538 3.2
R17478 vss.n5273 vss.n5272 3.2
R17479 vss.n4552 vss.n4548 3.2
R17480 vss.n4570 vss.n4564 3.2
R17481 vss.n4578 vss.n4576 3.2
R17482 vss.n5235 vss.n5234 3.2
R17483 vss.n4587 vss.n4585 3.2
R17484 vss.n4597 vss.n4595 3.2
R17485 vss.n5212 vss.n5211 3.2
R17486 vss.n4606 vss.n4604 3.2
R17487 vss.n5191 vss.n4619 3.2
R17488 vss.n5183 vss.n5182 3.2
R17489 vss.n4633 vss.n4629 3.2
R17490 vss.n5168 vss.n4638 3.2
R17491 vss.n5160 vss.n5159 3.2
R17492 vss.n4652 vss.n4648 3.2
R17493 vss.n5145 vss.n4657 3.2
R17494 vss.n4678 vss.n4676 3.2
R17495 vss.n5122 vss.n5121 3.2
R17496 vss.n4687 vss.n4685 3.2
R17497 vss.n4697 vss.n4695 3.2
R17498 vss.n5099 vss.n5098 3.2
R17499 vss.n4706 vss.n4704 3.2
R17500 vss.n4716 vss.n4714 3.2
R17501 vss.n5069 vss.n5068 3.2
R17502 vss.n5063 vss.n4729 3.2
R17503 vss.n5055 vss.n5054 3.2
R17504 vss.n4746 vss.n4742 3.2
R17505 vss.n5040 vss.n4751 3.2
R17506 vss.n5032 vss.n5031 3.2
R17507 vss.n4765 vss.n4761 3.2
R17508 vss.n4783 vss.n4777 3.2
R17509 vss.n4791 vss.n4789 3.2
R17510 vss.n4994 vss.n4993 3.2
R17511 vss.n4800 vss.n4798 3.2
R17512 vss.n4810 vss.n4808 3.2
R17513 vss.n4971 vss.n4970 3.2
R17514 vss.n4819 vss.n4817 3.2
R17515 vss.n4950 vss.n4832 3.2
R17516 vss.n4942 vss.n4941 3.2
R17517 vss.n4846 vss.n4842 3.2
R17518 vss.n4927 vss.n4851 3.2
R17519 vss.n4919 vss.n4918 3.2
R17520 vss.n4865 vss.n4861 3.2
R17521 vss.n4904 vss.n4870 3.2
R17522 vss.n4884 vss.n4883 3.2
R17523 vss.n6902 vss.n6901 3.2
R17524 vss.n6882 vss.n5652 3.2
R17525 vss.n5665 vss.n5662 3.2
R17526 vss.n6869 vss.n6868 3.2
R17527 vss.n5674 vss.n5672 3.2
R17528 vss.n5684 vss.n5682 3.2
R17529 vss.n6846 vss.n6845 3.2
R17530 vss.n5693 vss.n5691 3.2
R17531 vss.n6825 vss.n5706 3.2
R17532 vss.n6817 vss.n6816 3.2
R17533 vss.n5720 vss.n5716 3.2
R17534 vss.n6802 vss.n5725 3.2
R17535 vss.n6794 vss.n6793 3.2
R17536 vss.n5739 vss.n5735 3.2
R17537 vss.n6779 vss.n5744 3.2
R17538 vss.n6759 vss.n6758 3.2
R17539 vss.n6751 vss.n5763 3.2
R17540 vss.n5775 vss.n5772 3.2
R17541 vss.n6738 vss.n6737 3.2
R17542 vss.n5784 vss.n5782 3.2
R17543 vss.n5794 vss.n5792 3.2
R17544 vss.n6715 vss.n6714 3.2
R17545 vss.n6697 vss.n6696 3.2
R17546 vss.n6691 vss.n5810 3.2
R17547 vss.n6683 vss.n6682 3.2
R17548 vss.n5827 vss.n5823 3.2
R17549 vss.n6668 vss.n5832 3.2
R17550 vss.n6660 vss.n6659 3.2
R17551 vss.n5846 vss.n5842 3.2
R17552 vss.n5864 vss.n5858 3.2
R17553 vss.n5872 vss.n5870 3.2
R17554 vss.n6622 vss.n6621 3.2
R17555 vss.n5881 vss.n5879 3.2
R17556 vss.n5891 vss.n5889 3.2
R17557 vss.n6599 vss.n6598 3.2
R17558 vss.n5900 vss.n5898 3.2
R17559 vss.n6578 vss.n5913 3.2
R17560 vss.n6570 vss.n6569 3.2
R17561 vss.n5927 vss.n5923 3.2
R17562 vss.n6555 vss.n5932 3.2
R17563 vss.n6547 vss.n6546 3.2
R17564 vss.n5946 vss.n5942 3.2
R17565 vss.n6532 vss.n5951 3.2
R17566 vss.n6512 vss.n6511 3.2
R17567 vss.n6504 vss.n5970 3.2
R17568 vss.n5982 vss.n5979 3.2
R17569 vss.n6491 vss.n6490 3.2
R17570 vss.n5991 vss.n5989 3.2
R17571 vss.n6001 vss.n5999 3.2
R17572 vss.n6468 vss.n6467 3.2
R17573 vss.n6450 vss.n6449 3.2
R17574 vss.n6444 vss.n6017 3.2
R17575 vss.n6436 vss.n6435 3.2
R17576 vss.n6034 vss.n6030 3.2
R17577 vss.n6421 vss.n6039 3.2
R17578 vss.n6413 vss.n6412 3.2
R17579 vss.n6053 vss.n6049 3.2
R17580 vss.n6071 vss.n6065 3.2
R17581 vss.n6079 vss.n6077 3.2
R17582 vss.n6375 vss.n6374 3.2
R17583 vss.n6088 vss.n6086 3.2
R17584 vss.n6098 vss.n6096 3.2
R17585 vss.n6352 vss.n6351 3.2
R17586 vss.n6107 vss.n6105 3.2
R17587 vss.n6331 vss.n6120 3.2
R17588 vss.n6323 vss.n6322 3.2
R17589 vss.n6134 vss.n6130 3.2
R17590 vss.n6308 vss.n6139 3.2
R17591 vss.n6300 vss.n6299 3.2
R17592 vss.n6153 vss.n6149 3.2
R17593 vss.n6285 vss.n6158 3.2
R17594 vss.n6265 vss.n6264 3.2
R17595 vss.n6257 vss.n6177 3.2
R17596 vss.n6189 vss.n6186 3.2
R17597 vss.n6244 vss.n6243 3.2
R17598 vss.n6207 vss.n6196 3.2
R17599 vss.n18951 vss.n17684 3.155
R17600 vss.n17685 vss.n17684 3.155
R17601 vss.n17791 vss.n17785 3.155
R17602 vss.n17792 vss.n17791 3.155
R17603 vss.n17898 vss.n17892 3.155
R17604 vss.n17898 vss.n17895 3.155
R17605 vss.n18004 vss.n17998 3.155
R17606 vss.n18005 vss.n18004 3.155
R17607 vss.n18111 vss.n18105 3.155
R17608 vss.n18111 vss.n18108 3.155
R17609 vss.n18217 vss.n18211 3.155
R17610 vss.n18218 vss.n18217 3.155
R17611 vss.n19091 vss.n19085 3.155
R17612 vss.n19092 vss.n19091 3.155
R17613 vss.n20097 vss.n19191 3.155
R17614 vss.n19192 vss.n19191 3.155
R17615 vss.n19298 vss.n19292 3.155
R17616 vss.n19299 vss.n19298 3.155
R17617 vss.n19850 vss.n19397 3.155
R17618 vss.n19398 vss.n19397 3.155
R17619 vss.n19505 vss.n19499 3.155
R17620 vss.n19506 vss.n19505 3.155
R17621 vss.n5561 vss.n4294 3.155
R17622 vss.n4295 vss.n4294 3.155
R17623 vss.n4401 vss.n4395 3.155
R17624 vss.n4402 vss.n4401 3.155
R17625 vss.n4508 vss.n4502 3.155
R17626 vss.n4508 vss.n4505 3.155
R17627 vss.n4614 vss.n4608 3.155
R17628 vss.n4615 vss.n4614 3.155
R17629 vss.n4721 vss.n4715 3.155
R17630 vss.n4721 vss.n4718 3.155
R17631 vss.n4827 vss.n4821 3.155
R17632 vss.n4828 vss.n4827 3.155
R17633 vss.n5701 vss.n5695 3.155
R17634 vss.n5702 vss.n5701 3.155
R17635 vss.n6707 vss.n5801 3.155
R17636 vss.n5802 vss.n5801 3.155
R17637 vss.n5908 vss.n5902 3.155
R17638 vss.n5909 vss.n5908 3.155
R17639 vss.n6460 vss.n6007 3.155
R17640 vss.n6008 vss.n6007 3.155
R17641 vss.n6115 vss.n6109 3.155
R17642 vss.n6116 vss.n6115 3.155
R17643 vss.n15881 vss.n15880 3.105
R17644 vss.n9640 vss.n9639 3.1
R17645 vss.n9655 vss.n9654 3.1
R17646 vss.n12630 vss.n12629 3.1
R17647 vss.n12206 vss.n12094 3.1
R17648 vss.n11966 vss.n11965 3.1
R17649 vss.n11215 vss.n10994 3.1
R17650 vss.n11900 vss.n11891 3.1
R17651 vss.n11424 vss.n11415 3.1
R17652 vss.n14139 vss.n14130 3.1
R17653 vss.n14139 vss.n14138 3.1
R17654 vss.n11900 vss.n11899 3.1
R17655 vss.n10619 vss.n10610 3.1
R17656 vss.n10619 vss.n10618 3.1
R17657 vss.n12731 vss.n10469 3.1
R17658 vss.n11424 vss.n11423 3.1
R17659 vss.n11138 vss.n11109 3.1
R17660 vss.n13893 vss.n13892 3.1
R17661 vss.n11641 vss.n11603 3.1
R17662 vss.n14764 vss.n14763 3.1
R17663 vss.n14605 vss.n13553 3.1
R17664 vss.n14439 vss.n14438 3.1
R17665 vss.n14938 vss.n14937 3.1
R17666 vss.n16074 vss.n16073 3.1
R17667 vss.n13406 vss.n13405 3.099
R17668 vss.n20894 vss.n17485 3.069
R17669 vss.n21101 vss.n17474 3.069
R17670 vss.n21102 vss.n17463 3.069
R17671 vss.n21309 vss.n17452 3.069
R17672 vss.n21310 vss.n17441 3.069
R17673 vss.n21517 vss.n17430 3.069
R17674 vss.n21518 vss.n17419 3.069
R17675 vss.n7504 vss.n4095 3.069
R17676 vss.n7711 vss.n4084 3.069
R17677 vss.n7712 vss.n4073 3.069
R17678 vss.n7920 vss.n4062 3.069
R17679 vss.n7921 vss.n4051 3.069
R17680 vss.n8128 vss.n4040 3.069
R17681 vss.n8129 vss.n4029 3.069
R17682 vss.n8336 vss.n3555 3.069
R17683 vss.n8337 vss.n3544 3.069
R17684 vss.n8544 vss.n3533 3.069
R17685 vss.n8545 vss.n3522 3.069
R17686 vss.n8752 vss.n3511 3.069
R17687 vss.n8753 vss.n3500 3.069
R17688 vss.n22173 vss.n17397 3.069
R17689 vss.n22174 vss.n17386 3.069
R17690 vss.n22381 vss.n17375 3.069
R17691 vss.n22382 vss.n17364 3.069
R17692 vss.n22589 vss.n17353 3.069
R17693 vss.n22590 vss.n17342 3.069
R17694 vss.n9069 vss.n9067 3.067
R17695 vss.n12160 vss.n12102 3.062
R17696 vss.n11879 vss.n11337 3.062
R17697 vss.n12644 vss.n12447 3.062
R17698 vss.n14320 vss.n14289 3.062
R17699 vss.n11729 vss.n11712 3.062
R17700 vss.n13320 vss.n13283 3.062
R17701 vss.n15038 vss.n12788 3.062
R17702 vss.n14925 vss.n13211 3.062
R17703 vss.n11994 vss.n10871 3.062
R17704 vss.n11239 vss.n11237 3.062
R17705 vss.n13727 vss.n13724 3.062
R17706 vss.n11879 vss.n11344 3.062
R17707 vss.n14151 vss.n14150 3.062
R17708 vss.n14151 vss.n13605 3.062
R17709 vss.n13727 vss.n13718 3.062
R17710 vss.n13066 vss.n13063 3.062
R17711 vss.n13066 vss.n13053 3.062
R17712 vss.n14026 vss.n14024 3.062
R17713 vss.n14451 vss.n14180 3.062
R17714 vss.n14644 vss.n13524 3.062
R17715 vss.n22085 vss.n22082 3.04
R17716 vss.n21655 vss.n21641 3.033
R17717 vss.n21800 vss.n21643 3.033
R17718 vss.n10417 vss.n10416 3.033
R17719 vss.n14823 vss.n14822 3.033
R17720 vss.n14826 vss.n14825 3.033
R17721 vss.n14850 vss.n14849 3.033
R17722 vss.n12727 vss.n12726 3.033
R17723 vss.n12104 vss.n12103 3.033
R17724 vss.n12108 vss.n12107 3.033
R17725 vss.n3604 vss.n3590 3.033
R17726 vss.n3749 vss.n3592 3.033
R17727 vss.n20378 vss.n17575 3.032
R17728 vss.n6988 vss.n4185 3.032
R17729 vss.n14107 vss.n13615 3.024
R17730 vss.n13465 vss.n13429 3.024
R17731 vss.n12727 vss.n10499 3.024
R17732 vss.n14954 vss.n13200 3.024
R17733 vss.n12605 vss.n12520 3.024
R17734 vss.n11440 vss.n11404 3.024
R17735 vss.n11440 vss.n11396 3.024
R17736 vss.n14107 vss.n13625 3.024
R17737 vss.n10635 vss.n10591 3.024
R17738 vss.n13465 vss.n13438 3.024
R17739 vss.n10635 vss.n10599 3.024
R17740 vss.n11653 vss.n11652 3.024
R17741 vss.n13927 vss.n13926 3.024
R17742 vss.n13811 vss.n13807 3.022
R17743 vss.n13716 vss.n13713 3.022
R17744 vss.n11423 vss.n11418 3.022
R17745 vss.n14178 vss.n14173 3.022
R17746 vss.n14438 vss.n14433 3.022
R17747 vss.n14287 vss.n14283 3.022
R17748 vss.n13892 vss.n13887 3.022
R17749 vss.n13774 vss.n13773 3.022
R17750 vss.n13604 vss.n13600 3.022
R17751 vss.n14138 vss.n14137 3.022
R17752 vss.n11530 vss.n11526 3.022
R17753 vss.n11710 vss.n11706 3.022
R17754 vss.n11109 vss.n11108 3.022
R17755 vss.n11236 vss.n11235 3.022
R17756 vss.n10994 vss.n10988 3.022
R17757 vss.n11335 vss.n11331 3.022
R17758 vss.n11899 vss.n11898 3.022
R17759 vss.n12370 vss.n12369 3.022
R17760 vss.n10869 vss.n10859 3.022
R17761 vss.n11965 vss.n11960 3.022
R17762 vss.n12286 vss.n12282 3.022
R17763 vss.n12279 vss.n12278 3.022
R17764 vss.n10766 vss.n10762 3.022
R17765 vss.n12101 vss.n12100 3.022
R17766 vss.n12094 vss.n12093 3.022
R17767 vss.n12445 vss.n12438 3.022
R17768 vss.n12629 vss.n12628 3.022
R17769 vss.n12786 vss.n12779 3.022
R17770 vss.n10469 vss.n10468 3.022
R17771 vss.n13170 vss.n13166 3.022
R17772 vss.n13209 vss.n13201 3.022
R17773 vss.n14937 vss.n14936 3.022
R17774 vss.n13282 vss.n13279 3.022
R17775 vss.n14763 vss.n14758 3.022
R17776 vss.n13523 vss.n13519 3.022
R17777 vss.n13553 vss.n13547 3.022
R17778 vss.n14148 vss.n14144 3.022
R17779 vss.n14130 vss.n14125 3.022
R17780 vss.n12960 vss.n12959 3.022
R17781 vss.n13485 vss.n13481 3.022
R17782 vss.n13478 vss.n13477 3.022
R17783 vss.n13394 vss.n13390 3.022
R17784 vss.n13405 vss.n13400 3.022
R17785 vss.n12929 vss.n12928 3.022
R17786 vss.n11342 vss.n11338 3.022
R17787 vss.n11891 vss.n11886 3.022
R17788 vss.n10711 vss.n10707 3.022
R17789 vss.n13062 vss.n13055 3.022
R17790 vss.n10610 vss.n10609 3.022
R17791 vss.n13001 vss.n13000 3.022
R17792 vss.n13723 vss.n13720 3.022
R17793 vss.n11415 vss.n11410 3.022
R17794 vss.n10565 vss.n10564 3.022
R17795 vss.n13051 vss.n13048 3.022
R17796 vss.n10618 vss.n10613 3.022
R17797 vss.n12350 vss.n12349 3.022
R17798 vss.n14023 vss.n14015 3.022
R17799 vss.n11603 vss.n11598 3.022
R17800 vss.n11510 vss.n11509 3.022
R17801 vss.n20476 vss.n20475 3.011
R17802 vss.n20597 vss.n20596 3.011
R17803 vss.n20705 vss.n20704 3.011
R17804 vss.n20820 vss.n20819 3.011
R17805 vss.n21880 vss.n21879 3.011
R17806 vss.n21780 vss.n21779 3.011
R17807 vss.n12538 vss.n12537 3.011
R17808 vss.n12540 vss.n12539 3.011
R17809 vss.n12180 vss.n12179 3.011
R17810 vss.n10850 vss.n10849 3.011
R17811 vss.n11293 vss.n11292 3.011
R17812 vss.n11154 vss.n11153 3.011
R17813 vss.n14292 vss.n14291 3.011
R17814 vss.n14005 vss.n14004 3.011
R17815 vss.n11794 vss.n11793 3.011
R17816 vss.n11078 vss.n11077 3.011
R17817 vss.n14782 vss.n14781 3.011
R17818 vss.n13526 vss.n13525 3.011
R17819 vss.n14517 vss.n14516 3.011
R17820 vss.n14235 vss.n14234 3.011
R17821 vss.n14880 vss.n14870 3.011
R17822 vss.n14872 vss.n14871 3.011
R17823 vss.n12772 vss.n12771 3.011
R17824 vss.n12774 vss.n12773 3.011
R17825 vss.n12691 vss.n12681 3.011
R17826 vss.n12683 vss.n12682 3.011
R17827 vss.n3829 vss.n3828 3.011
R17828 vss.n3729 vss.n3728 3.011
R17829 vss.n7086 vss.n7085 3.011
R17830 vss.n7207 vss.n7206 3.011
R17831 vss.n7315 vss.n7314 3.011
R17832 vss.n7430 vss.n7429 3.011
R17833 vss.n1699 vss.n1698 3.011
R17834 vss.n1818 vss.n1817 3.011
R17835 vss.n1929 vss.n1928 3.011
R17836 vss.n2058 vss.n2057 3.011
R17837 vss.n2173 vss.n2172 3.011
R17838 vss.n2303 vss.n2302 3.011
R17839 vss.n2418 vss.n2417 3.011
R17840 vss.n2547 vss.n2546 3.011
R17841 vss.n2662 vss.n2661 3.011
R17842 vss.n2791 vss.n2790 3.011
R17843 vss.n2900 vss.n2899 3.011
R17844 vss.n3030 vss.n3029 3.011
R17845 vss.n3145 vss.n3144 3.011
R17846 vss.n3274 vss.n3273 3.011
R17847 vss.n3386 vss.n3385 3.011
R17848 vss.n15159 vss.n15158 3.011
R17849 vss.n160 vss.n159 3.011
R17850 vss.n279 vss.n278 3.011
R17851 vss.n390 vss.n389 3.011
R17852 vss.n519 vss.n518 3.011
R17853 vss.n634 vss.n633 3.011
R17854 vss.n764 vss.n763 3.011
R17855 vss.n879 vss.n878 3.011
R17856 vss.n1008 vss.n1007 3.011
R17857 vss.n1123 vss.n1122 3.011
R17858 vss.n1252 vss.n1251 3.011
R17859 vss.n23347 vss.n23346 3.011
R17860 vss.n23218 vss.n23217 3.011
R17861 vss.n23103 vss.n23102 3.011
R17862 vss.n22974 vss.n22973 3.011
R17863 vss.n22863 vss.n22862 3.011
R17864 vss.n22793 vss.n22792 3.011
R17865 vss.n21817 vss.n21816 2.992
R17866 vss.n3766 vss.n3765 2.992
R17867 vss.n11863 vss.n11353 2.987
R17868 vss.n13743 vss.n13701 2.986
R17869 vss.n13743 vss.n13712 2.986
R17870 vss.n11863 vss.n11362 2.986
R17871 vss.n13082 vss.n13047 2.986
R17872 vss.n12304 vss.n10761 2.986
R17873 vss.n12304 vss.n10751 2.986
R17874 vss.n13082 vss.n13037 2.986
R17875 vss.n15022 vss.n12798 2.986
R17876 vss.n13247 vss.n13220 2.986
R17877 vss.n21812 vss.n21811 2.975
R17878 vss.n3761 vss.n3760 2.975
R17879 vss.n9639 vss.n9636 2.965
R17880 vss.n12102 vss.n12096 2.962
R17881 vss.n13283 vss.n13278 2.962
R17882 vss.n14180 vss.n14179 2.961
R17883 vss.n11237 vss.n11227 2.961
R17884 vss.n10871 vss.n10870 2.961
R17885 vss.n13524 vss.n13518 2.961
R17886 vss.n20316 vss.n20315 2.955
R17887 vss.n6926 vss.n6925 2.955
R17888 vss.n12639 vss.n12485 2.953
R17889 vss.n20346 vss.n20345 2.941
R17890 vss.n20345 vss.n20344 2.941
R17891 vss.n6956 vss.n6955 2.941
R17892 vss.n6955 vss.n6954 2.941
R17893 vss.n21984 vss.n21981 2.94
R17894 vss.n21613 vss.n21610 2.94
R17895 vss.n3933 vss.n3930 2.94
R17896 vss.n3562 vss.n3559 2.94
R17897 vss.n15213 vss.t359 2.935
R17898 vss.n13217 vss.n13216 2.933
R17899 vss.n13328 vss.n13327 2.933
R17900 vss.n14035 vss.n14034 2.933
R17901 vss.n13132 vss.n13131 2.925
R17902 vss.n13673 vss.n13672 2.925
R17903 vss.n10652 vss.n10651 2.925
R17904 vss.n11457 vss.n11456 2.925
R17905 vss.n12277 vss.n12276 2.907
R17906 vss.n10617 vss.n10616 2.907
R17907 vss.n10467 vss.n10466 2.907
R17908 vss.n10608 vss.n10607 2.907
R17909 vss.n11414 vss.n11413 2.907
R17910 vss.n11890 vss.n11889 2.907
R17911 vss.n14289 vss.n14288 2.903
R17912 vss.n11712 vss.n11711 2.903
R17913 vss.n11337 vss.n11336 2.903
R17914 vss.n12447 vss.n12446 2.903
R17915 vss.n12788 vss.n12787 2.903
R17916 vss.n13211 vss.n13210 2.903
R17917 vss.n13718 vss.n13717 2.903
R17918 vss.n13605 vss.n13599 2.903
R17919 vss.n14150 vss.n14149 2.903
R17920 vss.n11344 vss.n11343 2.903
R17921 vss.n13063 vss.n13054 2.903
R17922 vss.n13724 vss.n13719 2.903
R17923 vss.n13053 vss.n13052 2.903
R17924 vss.n14024 vss.n14014 2.903
R17925 vss.n21820 vss.n21814 2.876
R17926 vss.n12716 vss.n10520 2.876
R17927 vss.n12731 vss.n10490 2.876
R17928 vss.n3769 vss.n3763 2.876
R17929 vss.n13801 vss.n13800 2.844
R17930 vss.n11417 vss.n11416 2.844
R17931 vss.n14432 vss.n14431 2.844
R17932 vss.n13886 vss.n13885 2.844
R17933 vss.n13760 vss.n13759 2.844
R17934 vss.n14132 vss.n14131 2.844
R17935 vss.n11533 vss.n11532 2.844
R17936 vss.n11103 vss.n11102 2.844
R17937 vss.n10987 vss.n10986 2.844
R17938 vss.n11893 vss.n11892 2.844
R17939 vss.n12373 vss.n12372 2.844
R17940 vss.n11959 vss.n11958 2.844
R17941 vss.n12287 vss.n12281 2.844
R17942 vss.n12272 vss.n12271 2.844
R17943 vss.n10772 vss.n10771 2.844
R17944 vss.n12087 vss.n12086 2.844
R17945 vss.n12623 vss.n12622 2.844
R17946 vss.n10462 vss.n10461 2.844
R17947 vss.n13175 vss.n13174 2.844
R17948 vss.n14931 vss.n14930 2.844
R17949 vss.n14757 vss.n14756 2.844
R17950 vss.n13546 vss.n13545 2.844
R17951 vss.n14124 vss.n14123 2.844
R17952 vss.n12965 vss.n12964 2.844
R17953 vss.n13486 vss.n13480 2.844
R17954 vss.n13472 vss.n13471 2.844
R17955 vss.n13399 vss.n13398 2.844
R17956 vss.n12934 vss.n12933 2.844
R17957 vss.n11885 vss.n11884 2.844
R17958 vss.n10714 vss.n10713 2.844
R17959 vss.n10603 vss.n10602 2.844
R17960 vss.n13004 vss.n13003 2.844
R17961 vss.n11409 vss.n11408 2.844
R17962 vss.n10552 vss.n10551 2.844
R17963 vss.n10612 vss.n10611 2.844
R17964 vss.n12336 vss.n12335 2.844
R17965 vss.n11597 vss.n11596 2.844
R17966 vss.n11497 vss.n11496 2.844
R17967 vss.n12953 vss.n12952 2.835
R17968 vss.n12994 vss.n12993 2.835
R17969 vss.n12393 vss.n12382 2.835
R17970 vss.n10724 vss.n10723 2.835
R17971 vss.n13798 vss.n13787 2.835
R17972 vss.n11524 vss.n11523 2.835
R17973 vss.n12122 vss.n12121 2.826
R17974 vss.n13276 vss.n13275 2.826
R17975 vss.n12135 vss.n12131 2.826
R17976 vss.n13263 vss.n13259 2.826
R17977 vss.n12642 vss.n12468 2.804
R17978 vss.n9666 vss.n9663 2.8
R17979 vss.n9139 vss.n9138 2.782
R17980 vss.n10228 vss.n10227 2.742
R17981 vss.n12734 vss.n10460 2.735
R17982 vss.n12713 vss.n10550 2.735
R17983 vss.n12146 vss.n12145 2.709
R17984 vss.n14818 vss.n14817 2.709
R17985 vss.n3425 vss.n3424 2.709
R17986 vss.n3466 vss.n3465 2.709
R17987 vss.n22840 vss.n22839 2.709
R17988 vss.n1441 vss.n1440 2.709
R17989 vss.n11169 vss.n11044 2.682
R17990 vss.n14410 vss.n14392 2.682
R17991 vss.n12588 vss.n12569 2.682
R17992 vss.n13308 vss.n13290 2.682
R17993 vss.n11169 vss.n11056 2.679
R17994 vss.n14410 vss.n14404 2.679
R17995 vss.n12588 vss.n12587 2.679
R17996 vss.n12661 vss.n12429 2.679
R17997 vss.n13308 vss.n13302 2.679
R17998 vss.n15816 vss.n15795 2.678
R17999 vss.n17317 vss.n17296 2.678
R18000 vss.n17317 vss.n17275 2.676
R18001 vss.n15816 vss.n15805 2.675
R18002 vss.n17317 vss.n17306 2.675
R18003 vss.n15816 vss.n15815 2.673
R18004 vss.n17317 vss.n17316 2.672
R18005 vss.n17317 vss.n17285 2.672
R18006 vss.n21796 vss.n21658 2.671
R18007 vss.n3745 vss.n3607 2.671
R18008 vss.n21983 vss.n21982 2.67
R18009 vss.n21742 vss.n21712 2.67
R18010 vss.n21612 vss.n21611 2.67
R18011 vss.n3932 vss.n3931 2.67
R18012 vss.n3691 vss.n3661 2.67
R18013 vss.n3561 vss.n3560 2.67
R18014 vss.n17588 vss.n17582 2.666
R18015 vss.n13693 vss.n13692 2.666
R18016 vss.n14344 vss.n14343 2.666
R18017 vss.n14478 vss.n14477 2.666
R18018 vss.n11770 vss.n11769 2.666
R18019 vss.n11346 vss.n11345 2.666
R18020 vss.n10754 vss.n10753 2.666
R18021 vss.n10743 vss.n10742 2.666
R18022 vss.n12432 vss.n12431 2.666
R18023 vss.n12791 vss.n12790 2.666
R18024 vss.n13214 vss.n13213 2.666
R18025 vss.n13568 vss.n13567 2.666
R18026 vss.n14648 vss.n14647 2.666
R18027 vss.n13325 vss.n13324 2.666
R18028 vss.n11355 vss.n11354 2.666
R18029 vss.n13040 vss.n13039 2.666
R18030 vss.n13705 vss.n13704 2.666
R18031 vss.n13029 vss.n13028 2.666
R18032 vss.n14032 vss.n14031 2.666
R18033 vss.n4198 vss.n4192 2.666
R18034 vss.n11709 vss.n11707 2.65
R18035 vss.n11334 vss.n11332 2.65
R18036 vss.n11341 vss.n11339 2.65
R18037 vss.n10765 vss.n10763 2.65
R18038 vss.n12444 vss.n12442 2.65
R18039 vss.n14147 vss.n14145 2.65
R18040 vss.n13484 vss.n13482 2.65
R18041 vss.n13393 vss.n13392 2.65
R18042 vss.n14022 vss.n14020 2.65
R18043 vss.n22016 vss.n22015 2.648
R18044 vss.n3965 vss.n3964 2.648
R18045 vss.n20469 vss.n20461 2.635
R18046 vss.n20620 vss.n20612 2.635
R18047 vss.n20698 vss.n20690 2.635
R18048 vss.n20843 vss.n20835 2.635
R18049 vss.n21791 vss.n21686 2.635
R18050 vss.n21657 vss.n21655 2.635
R18051 vss.n12559 vss.n12546 2.635
R18052 vss.n12561 vss.n12559 2.635
R18053 vss.n12201 vss.n12194 2.635
R18054 vss.n12005 vss.n11998 2.635
R18055 vss.n11284 vss.n11277 2.635
R18056 vss.n11182 vss.n11175 2.635
R18057 vss.n13881 vss.n13874 2.635
R18058 vss.n13991 vss.n13984 2.635
R18059 vss.n11785 vss.n11778 2.635
R18060 vss.n11095 vss.n11088 2.635
R18061 vss.n14775 vss.n14768 2.635
R18062 vss.n13516 vss.n13509 2.635
R18063 vss.n14508 vss.n14501 2.635
R18064 vss.n14222 vss.n14215 2.635
R18065 vss.n12843 vss.n12842 2.635
R18066 vss.n12842 vss.n12835 2.635
R18067 vss.n12815 vss.n12802 2.635
R18068 vss.n12817 vss.n12815 2.635
R18069 vss.n12674 vss.n12673 2.635
R18070 vss.n12673 vss.n12666 2.635
R18071 vss.n3740 vss.n3635 2.635
R18072 vss.n3606 vss.n3604 2.635
R18073 vss.n7079 vss.n7071 2.635
R18074 vss.n7230 vss.n7222 2.635
R18075 vss.n7308 vss.n7300 2.635
R18076 vss.n7453 vss.n7445 2.635
R18077 vss.n1692 vss.n1684 2.635
R18078 vss.n1841 vss.n1833 2.635
R18079 vss.n1922 vss.n1913 2.635
R18080 vss.n2083 vss.n2074 2.635
R18081 vss.n2166 vss.n2157 2.635
R18082 vss.n2328 vss.n2319 2.635
R18083 vss.n2411 vss.n2402 2.635
R18084 vss.n2572 vss.n2563 2.635
R18085 vss.n2655 vss.n2646 2.635
R18086 vss.n2815 vss.n2807 2.635
R18087 vss.n2893 vss.n2884 2.635
R18088 vss.n3055 vss.n3046 2.635
R18089 vss.n3138 vss.n3129 2.635
R18090 vss.n3299 vss.n3290 2.635
R18091 vss.n3379 vss.n3371 2.635
R18092 vss.n3488 vss.n3480 2.635
R18093 vss.n153 vss.n145 2.635
R18094 vss.n302 vss.n294 2.635
R18095 vss.n383 vss.n374 2.635
R18096 vss.n544 vss.n535 2.635
R18097 vss.n627 vss.n618 2.635
R18098 vss.n789 vss.n780 2.635
R18099 vss.n872 vss.n863 2.635
R18100 vss.n1033 vss.n1024 2.635
R18101 vss.n1116 vss.n1107 2.635
R18102 vss.n1277 vss.n1268 2.635
R18103 vss.n23372 vss.n23363 2.635
R18104 vss.n23211 vss.n23202 2.635
R18105 vss.n23128 vss.n23119 2.635
R18106 vss.n22967 vss.n22958 2.635
R18107 vss.n22886 vss.n22878 2.635
R18108 vss.n1463 vss.n1455 2.635
R18109 vss.n22045 vss.n22044 2.599
R18110 vss.n3994 vss.n3993 2.599
R18111 vss.n19612 vss.n19611 2.577
R18112 vss.n6222 vss.n6221 2.577
R18113 vss.n10560 vss.n10558 2.549
R18114 vss.n12345 vss.n12343 2.549
R18115 vss.n13769 vss.n13767 2.549
R18116 vss.n11505 vss.n11503 2.549
R18117 vss.n12932 vss.n12930 2.545
R18118 vss.n12963 vss.n12961 2.545
R18119 vss.n11389 vss.n11388 2.488
R18120 vss.n13920 vss.n13919 2.488
R18121 vss.n13607 vss.n13606 2.488
R18122 vss.n11019 vss.n11018 2.488
R18123 vss.n11266 vss.n11265 2.488
R18124 vss.n10832 vss.n10831 2.488
R18125 vss.n12232 vss.n12231 2.488
R18126 vss.n12513 vss.n12512 2.488
R18127 vss.n10492 vss.n10491 2.488
R18128 vss.n13193 vss.n13192 2.488
R18129 vss.n13617 vss.n13616 2.488
R18130 vss.n13422 vss.n13421 2.488
R18131 vss.n13431 vss.n13430 2.488
R18132 vss.n10912 vss.n10911 2.488
R18133 vss.n10585 vss.n10584 2.488
R18134 vss.n11399 vss.n11398 2.488
R18135 vss.n10594 vss.n10593 2.488
R18136 vss.n11646 vss.n11645 2.488
R18137 vss.n9713 vss.n9699 2.479
R18138 vss.n9709 vss.n9708 2.479
R18139 vss.n10214 vss.n10213 2.479
R18140 vss.n21649 vss.n21646 2.476
R18141 vss.n3598 vss.n3595 2.476
R18142 vss.n20893 vss.n20892 2.471
R18143 vss.n16674 vss.n16673 2.444
R18144 vss.n7503 vss.n7502 2.442
R18145 vss.n14243 vss.n14242 2.423
R18146 vss.n22028 vss.n22027 2.422
R18147 vss.n3977 vss.n3976 2.422
R18148 vss.n21788 vss.n21689 2.422
R18149 vss.n3737 vss.n3638 2.422
R18150 vss.n19618 vss.n19591 2.4
R18151 vss.n6228 vss.n6201 2.4
R18152 vss.n14652 vss.n14649 2.376
R18153 vss.n22051 vss.n22050 2.356
R18154 vss.n4000 vss.n3999 2.356
R18155 vss.n10303 vss.n10301 2.349
R18156 vss.n10362 vss.n10360 2.349
R18157 vss.n21789 vss.n21772 2.344
R18158 vss.n3738 vss.n3721 2.344
R18159 vss.n14349 vss.n14345 2.332
R18160 vss.n13612 vss.n13611 2.332
R18161 vss.n12518 vss.n12517 2.332
R18162 vss.n13152 vss.n13151 2.325
R18163 vss.n13110 vss.n13109 2.325
R18164 vss.n10686 vss.n10685 2.325
R18165 vss.n12334 vss.n12333 2.325
R18166 vss.n13758 vss.n13660 2.325
R18167 vss.n14092 vss.n14087 2.325
R18168 vss.n11495 vss.n11494 2.325
R18169 vss.n11848 vss.n11847 2.325
R18170 vss.n17342 vss.n17341 2.323
R18171 vss.n17353 vss.n17352 2.323
R18172 vss.n17364 vss.n17363 2.323
R18173 vss.n17375 vss.n17374 2.323
R18174 vss.n17386 vss.n17385 2.323
R18175 vss.n17397 vss.n17396 2.323
R18176 vss.n17419 vss.n17418 2.323
R18177 vss.n17430 vss.n17429 2.323
R18178 vss.n17441 vss.n17440 2.323
R18179 vss.n17452 vss.n17451 2.323
R18180 vss.n17463 vss.n17462 2.323
R18181 vss.n17474 vss.n17473 2.323
R18182 vss.n17485 vss.n17484 2.323
R18183 vss.n3500 vss.n3499 2.323
R18184 vss.n3511 vss.n3510 2.323
R18185 vss.n3522 vss.n3521 2.323
R18186 vss.n3533 vss.n3532 2.323
R18187 vss.n3544 vss.n3543 2.323
R18188 vss.n3555 vss.n3554 2.323
R18189 vss.n4029 vss.n4028 2.323
R18190 vss.n4040 vss.n4039 2.323
R18191 vss.n4051 vss.n4050 2.323
R18192 vss.n4062 vss.n4061 2.323
R18193 vss.n4073 vss.n4072 2.323
R18194 vss.n4084 vss.n4083 2.323
R18195 vss.n4095 vss.n4094 2.323
R18196 vss.n8934 vss.n8923 2.317
R18197 vss.n8952 vss.n8948 2.317
R18198 vss.n10264 vss.n10254 2.315
R18199 vss.n10306 vss.n10297 2.315
R18200 vss.n10386 vss.n10357 2.315
R18201 vss.n15214 ldomc_0.vdm_0.vss 2.314
R18202 vss.n10283 vss.n10278 2.313
R18203 vss.n13451 vss.n13450 2.295
R18204 vss.n13096 vss.n13027 2.295
R18205 vss.n10649 vss.n10582 2.295
R18206 vss.n12318 vss.n10741 2.295
R18207 vss.n14093 vss.n13637 2.295
R18208 vss.n13757 vss.n13691 2.295
R18209 vss.n11454 vss.n11386 2.295
R18210 vss.n11849 vss.n11374 2.295
R18211 vss.n20308 vss.n20307 2.293
R18212 vss.n6918 vss.n6917 2.293
R18213 vss.n13440 vss.n13439 2.281
R18214 vss.n13026 vss.n13025 2.281
R18215 vss.n10572 vss.n10571 2.281
R18216 vss.n10740 vss.n10739 2.281
R18217 vss.n13627 vss.n13626 2.281
R18218 vss.n13690 vss.n13689 2.281
R18219 vss.n11376 vss.n11375 2.281
R18220 vss.n11373 vss.n11372 2.281
R18221 vss.n21753 vss.n21752 2.276
R18222 vss.n3702 vss.n3701 2.276
R18223 vss.n17333 vss.n17332 2.275
R18224 vss.n17344 vss.n17343 2.275
R18225 vss.n17355 vss.n17354 2.275
R18226 vss.n17366 vss.n17365 2.275
R18227 vss.n17377 vss.n17376 2.275
R18228 vss.n17388 vss.n17387 2.275
R18229 vss.n17410 vss.n17409 2.275
R18230 vss.n17421 vss.n17420 2.275
R18231 vss.n17432 vss.n17431 2.275
R18232 vss.n17443 vss.n17442 2.275
R18233 vss.n17454 vss.n17453 2.275
R18234 vss.n17465 vss.n17464 2.275
R18235 vss.n17476 vss.n17475 2.275
R18236 vss.n3491 vss.n3490 2.275
R18237 vss.n3502 vss.n3501 2.275
R18238 vss.n3513 vss.n3512 2.275
R18239 vss.n3524 vss.n3523 2.275
R18240 vss.n3535 vss.n3534 2.275
R18241 vss.n3546 vss.n3545 2.275
R18242 vss.n4020 vss.n4019 2.275
R18243 vss.n4031 vss.n4030 2.275
R18244 vss.n4042 vss.n4041 2.275
R18245 vss.n4053 vss.n4052 2.275
R18246 vss.n4064 vss.n4063 2.275
R18247 vss.n4075 vss.n4074 2.275
R18248 vss.n4086 vss.n4085 2.275
R18249 vss.n20318 vss.n20317 2.273
R18250 vss.n6928 vss.n6927 2.273
R18251 vss.n20491 vss.n20490 2.258
R18252 vss.n20582 vss.n20581 2.258
R18253 vss.n20720 vss.n20719 2.258
R18254 vss.n20805 vss.n20804 2.258
R18255 vss.n21869 vss.n21868 2.258
R18256 vss.n21945 vss.n21944 2.258
R18257 vss.n21786 vss.n21775 2.258
R18258 vss.n12166 vss.n12165 2.258
R18259 vss.n11984 vss.n11983 2.258
R18260 vss.n11318 vss.n11317 2.258
R18261 vss.n14306 vss.n14305 2.258
R18262 vss.n11606 vss.n11605 2.258
R18263 vss.n11819 vss.n11818 2.258
R18264 vss.n14796 vss.n14795 2.258
R18265 vss.n14623 vss.n14622 2.258
R18266 vss.n14534 vss.n14533 2.258
R18267 vss.n14255 vss.n14254 2.258
R18268 vss.n14895 vss.n14885 2.258
R18269 vss.n14887 vss.n14886 2.258
R18270 vss.n15043 vss.n15042 2.258
R18271 vss.n15058 vss.n15057 2.258
R18272 vss.n12707 vss.n12697 2.258
R18273 vss.n12699 vss.n12698 2.258
R18274 vss.n3818 vss.n3817 2.258
R18275 vss.n3894 vss.n3893 2.258
R18276 vss.n3735 vss.n3724 2.258
R18277 vss.n7101 vss.n7100 2.258
R18278 vss.n7192 vss.n7191 2.258
R18279 vss.n7330 vss.n7329 2.258
R18280 vss.n7415 vss.n7414 2.258
R18281 vss.n1714 vss.n1713 2.258
R18282 vss.n1803 vss.n1802 2.258
R18283 vss.n1945 vss.n1944 2.258
R18284 vss.n2042 vss.n2041 2.258
R18285 vss.n2190 vss.n2189 2.258
R18286 vss.n2286 vss.n2285 2.258
R18287 vss.n2434 vss.n2433 2.258
R18288 vss.n2531 vss.n2530 2.258
R18289 vss.n2678 vss.n2677 2.258
R18290 vss.n2775 vss.n2774 2.258
R18291 vss.n2917 vss.n2916 2.258
R18292 vss.n3014 vss.n3013 2.258
R18293 vss.n3161 vss.n3160 2.258
R18294 vss.n3258 vss.n3257 2.258
R18295 vss.n3401 vss.n3400 2.258
R18296 vss.n3468 vss.n3467 2.258
R18297 vss.n175 vss.n174 2.258
R18298 vss.n264 vss.n263 2.258
R18299 vss.n406 vss.n405 2.258
R18300 vss.n503 vss.n502 2.258
R18301 vss.n651 vss.n650 2.258
R18302 vss.n747 vss.n746 2.258
R18303 vss.n895 vss.n894 2.258
R18304 vss.n992 vss.n991 2.258
R18305 vss.n1139 vss.n1138 2.258
R18306 vss.n1236 vss.n1235 2.258
R18307 vss.n23331 vss.n23330 2.258
R18308 vss.n23234 vss.n23233 2.258
R18309 vss.n23087 vss.n23086 2.258
R18310 vss.n22990 vss.n22989 2.258
R18311 vss.n22848 vss.n22847 2.258
R18312 vss.n1443 vss.n1442 2.258
R18313 vss.n22758 vss.n17331 2.255
R18314 vss.n17567 vss.n17558 2.251
R18315 vss.n4177 vss.n4168 2.251
R18316 vss.n11096 vss.n11095 2.25
R18317 vss.n14223 vss.n14222 2.25
R18318 vss.n20377 vss.n17574 2.25
R18319 vss.n21759 vss.n21758 2.25
R18320 vss.n21919 vss.n21821 2.25
R18321 vss.n21918 vss.n21917 2.25
R18322 vss.n21709 vss.n21704 2.25
R18323 vss.n21758 vss.n21698 2.25
R18324 vss.n21707 vss.n21704 2.25
R18325 vss.n10275 vss.n10274 2.25
R18326 vss.n10264 vss.n10263 2.25
R18327 vss.n10283 vss.n10282 2.25
R18328 vss.n10294 vss.n10293 2.25
R18329 vss.n10306 vss.n10305 2.25
R18330 vss.n10319 vss.n10318 2.25
R18331 vss.n10386 vss.n10385 2.25
R18332 vss.n8946 vss.n8945 2.25
R18333 vss.n8934 vss.n8933 2.25
R18334 vss.n8971 vss.n8970 2.25
R18335 vss.n8952 vss.n8951 2.25
R18336 vss.n3708 vss.n3707 2.25
R18337 vss.n3868 vss.n3770 2.25
R18338 vss.n3867 vss.n3866 2.25
R18339 vss.n3658 vss.n3653 2.25
R18340 vss.n3707 vss.n3647 2.25
R18341 vss.n3656 vss.n3653 2.25
R18342 vss.n6987 vss.n4184 2.25
R18343 vss.n15216 vss.n15215 2.25
R18344 vss.n21947 vss.n21946 2.248
R18345 vss.n22053 vss.n22052 2.248
R18346 vss.n3896 vss.n3895 2.248
R18347 vss.n4002 vss.n4001 2.248
R18348 vss.n17554 vss.n17550 2.247
R18349 vss.n21710 vss.n21704 2.247
R18350 vss.n3659 vss.n3653 2.247
R18351 vss.n4164 vss.n4160 2.247
R18352 vss.n21650 vss.n21645 2.246
R18353 vss.n3599 vss.n3594 2.246
R18354 vss.n20406 vss.n20405 2.246
R18355 vss.n7016 vss.n7015 2.246
R18356 vss.n17566 vss.n17558 2.246
R18357 vss.n4176 vss.n4168 2.246
R18358 vss.n21918 vss.n21913 2.245
R18359 vss.n3867 vss.n3862 2.245
R18360 vss.n20405 vss.n17555 2.245
R18361 vss.n7015 vss.n4165 2.245
R18362 vss.n21651 vss.n21650 2.244
R18363 vss.n3600 vss.n3599 2.244
R18364 vss.n20383 vss.n20382 2.241
R18365 vss.n6993 vss.n6992 2.241
R18366 vss.n20386 vss.n20385 2.241
R18367 vss.n6996 vss.n6995 2.241
R18368 vss.n21943 vss.n21942 2.24
R18369 vss.n3892 vss.n3891 2.24
R18370 vss.n22082 vss.n22081 2.227
R18371 vss.n9145 vss.n9143 2.2
R18372 vss.n16368 vss.n16363 2.176
R18373 vss.n16494 vss.n16493 2.176
R18374 vss.n16604 vss.n16599 2.176
R18375 vss.n16901 vss.n16900 2.176
R18376 vss.n17137 vss.n17136 2.176
R18377 vss.n15945 vss.n15940 2.176
R18378 vss.n16073 vss.n16072 2.176
R18379 vss.n16181 vss.n16176 2.176
R18380 vss.n15322 vss.n15321 2.176
R18381 vss.n15421 vss.n15416 2.176
R18382 vss.n15547 vss.n15546 2.176
R18383 vss.n15657 vss.n15652 2.176
R18384 vss.n15781 vss.n15780 2.176
R18385 ldomc_0.otaldom_0.ncsm_0.vss vss.n21801 2.172
R18386 bandgapmd_0.otam_1.ncsm_0.vss vss.n3750 2.172
R18387 vss.n22030 vss.n22029 2.172
R18388 vss.n21692 vss.n21690 2.172
R18389 vss.n3979 vss.n3978 2.172
R18390 vss.n3641 vss.n3639 2.172
R18391 vss.n1745 vss.n1744 2.169
R18392 vss.n206 vss.n205 2.169
R18393 vss.n22707 vss.n22698 2.133
R18394 vss.n22709 vss.n22707 2.133
R18395 vss.n22689 vss.n22688 2.133
R18396 vss.n22688 vss.n22679 2.133
R18397 vss.n22499 vss.n22490 2.133
R18398 vss.n22501 vss.n22499 2.133
R18399 vss.n22481 vss.n22480 2.133
R18400 vss.n22480 vss.n22471 2.133
R18401 vss.n22291 vss.n22282 2.133
R18402 vss.n22293 vss.n22291 2.133
R18403 vss.n22273 vss.n22272 2.133
R18404 vss.n22272 vss.n22263 2.133
R18405 vss.n22081 vss.n22072 2.133
R18406 vss.n21603 vss.n21602 2.133
R18407 vss.n21602 vss.n21593 2.133
R18408 vss.n21427 vss.n21418 2.133
R18409 vss.n21429 vss.n21427 2.133
R18410 vss.n21409 vss.n21408 2.133
R18411 vss.n21408 vss.n21399 2.133
R18412 vss.n21219 vss.n21210 2.133
R18413 vss.n21221 vss.n21219 2.133
R18414 vss.n21201 vss.n21200 2.133
R18415 vss.n21200 vss.n21191 2.133
R18416 vss.n21011 vss.n21002 2.133
R18417 vss.n21013 vss.n21011 2.133
R18418 vss.n20993 vss.n20992 2.133
R18419 vss.n20992 vss.n20983 2.133
R18420 vss.n8870 vss.n8861 2.133
R18421 vss.n8872 vss.n8870 2.133
R18422 vss.n8852 vss.n8851 2.133
R18423 vss.n8851 vss.n8842 2.133
R18424 vss.n8662 vss.n8653 2.133
R18425 vss.n8664 vss.n8662 2.133
R18426 vss.n8644 vss.n8643 2.133
R18427 vss.n8643 vss.n8634 2.133
R18428 vss.n8454 vss.n8445 2.133
R18429 vss.n8456 vss.n8454 2.133
R18430 vss.n8436 vss.n8435 2.133
R18431 vss.n8435 vss.n8426 2.133
R18432 vss.n8241 vss.n8232 2.133
R18433 vss.n8242 vss.n8241 2.133
R18434 vss.n8229 vss.n8228 2.133
R18435 vss.n8228 vss.n8219 2.133
R18436 vss.n8038 vss.n8029 2.133
R18437 vss.n8040 vss.n8038 2.133
R18438 vss.n8020 vss.n8019 2.133
R18439 vss.n8019 vss.n8010 2.133
R18440 vss.n7829 vss.n7820 2.133
R18441 vss.n7831 vss.n7829 2.133
R18442 vss.n7811 vss.n7810 2.133
R18443 vss.n7810 vss.n7801 2.133
R18444 vss.n7621 vss.n7612 2.133
R18445 vss.n7623 vss.n7621 2.133
R18446 vss.n7603 vss.n7602 2.133
R18447 vss.n7602 vss.n7593 2.133
R18448 vss.n8966 vss.n8964 2.111
R18449 vss.n12147 vss.n12122 2.102
R18450 vss.n14820 vss.n13276 2.102
R18451 vss.n12147 vss.n12135 2.102
R18452 vss.n14820 vss.n13263 2.102
R18453 vss.n22031 vss.n22030 2.093
R18454 vss.n21792 vss.n21690 2.093
R18455 vss.n3980 vss.n3979 2.093
R18456 vss.n3741 vss.n3639 2.093
R18457 vss.n11097 vss.n11066 2.093
R18458 vss.n14264 vss.n14233 2.093
R18459 vss.n12147 vss.n12146 2.085
R18460 vss.n14820 vss.n14818 2.085
R18461 vss.n3426 vss.n3425 2.085
R18462 vss.n15175 vss.n3466 2.085
R18463 vss.n22841 vss.n22840 2.085
R18464 vss.n22809 vss.n1441 2.085
R18465 vss.n21792 vss.n21689 2.079
R18466 vss.n3741 vss.n3638 2.079
R18467 vss.n22031 vss.n22028 2.079
R18468 vss.n11097 vss.n11076 2.079
R18469 vss.n14264 vss.n14253 2.079
R18470 vss.n3980 vss.n3977 2.079
R18471 vss.n22031 vss.n22016 2.072
R18472 vss.n11097 vss.n11096 2.072
R18473 vss.n14264 vss.n14223 2.072
R18474 vss.n3980 vss.n3965 2.072
R18475 vss.n14264 vss.n14243 2.07
R18476 vss.n11076 vss.n11075 2.056
R18477 vss.n14253 vss.n14252 2.056
R18478 vss.n16476 vss.n16469 2.048
R18479 vss.n16493 vss.n16484 2.048
R18480 vss.n16664 vss.n16663 2.048
R18481 vss.n16677 vss.n16676 2.048
R18482 vss.n16777 vss.n16770 2.048
R18483 vss.n16795 vss.n16786 2.048
R18484 vss.n16895 vss.n16894 2.048
R18485 vss.n16912 vss.n16911 2.048
R18486 vss.n17011 vss.n17002 2.048
R18487 vss.n17028 vss.n17027 2.048
R18488 vss.n17131 vss.n17130 2.048
R18489 vss.n17148 vss.n17147 2.048
R18490 vss.n17247 vss.n17238 2.048
R18491 vss.n17264 vss.n17255 2.048
R18492 vss.n15946 vss.n15939 2.048
R18493 vss.n15960 vss.n15959 2.048
R18494 vss.n16056 vss.n16049 2.048
R18495 vss.n16072 vss.n16063 2.048
R18496 vss.n16182 vss.n16175 2.048
R18497 vss.n16196 vss.n16195 2.048
R18498 vss.n16296 vss.n16295 2.048
R18499 vss.n15238 vss.n15229 2.048
R18500 vss.n15321 vss.n15314 2.048
R18501 vss.n15529 vss.n15522 2.048
R18502 vss.n15546 vss.n15537 2.048
R18503 vss.n15765 vss.n15758 2.048
R18504 vss.n15875 vss.n15874 2.048
R18505 vss.n15239 vss.n15238 2.047
R18506 vss.n15227 vss.n15226 2.047
R18507 vss.n16242 vss.n16241 2.027
R18508 vss.n14172 vss.n14171 2.025
R18509 vss.n13507 vss.n13506 2.025
R18510 vss.n13597 vss.n13592 2.025
R18511 vss.n13359 vss.n13358 2.025
R18512 vss.n13232 vss.n13231 2.025
R18513 vss.n13191 vss.n13190 2.025
R18514 vss.n12831 vss.n12830 2.025
R18515 vss.n10527 vss.n10521 2.025
R18516 vss.n14280 vss.n14279 2.025
R18517 vss.n13845 vss.n13844 2.025
R18518 vss.n11705 vss.n11704 2.025
R18519 vss.n13971 vss.n13970 2.025
R18520 vss.n11565 vss.n11560 2.025
R18521 vss.n12063 vss.n12062 2.025
R18522 vss.n12419 vss.n12418 2.025
R18523 vss.n12532 vss.n12531 2.025
R18524 vss.n10818 vss.n10817 2.025
R18525 vss.n10925 vss.n10924 2.025
R18526 vss.n10943 vss.n10942 2.025
R18527 vss.n11034 vss.n11033 2.025
R18528 ldomc_0.otaldom_0.vss vss.n20413 1.999
R18529 bandgapmd_0.otam_1.vss vss.n7023 1.999
R18530 vss.n22603 vss.n22593 1.991
R18531 vss.n22595 vss.n22594 1.991
R18532 vss.n22576 vss.n22575 1.991
R18533 vss.n22585 vss.n22584 1.991
R18534 vss.n22395 vss.n22385 1.991
R18535 vss.n22387 vss.n22386 1.991
R18536 vss.n22368 vss.n22367 1.991
R18537 vss.n22377 vss.n22376 1.991
R18538 vss.n22187 vss.n22177 1.991
R18539 vss.n22179 vss.n22178 1.991
R18540 vss.n22160 vss.n22159 1.991
R18541 vss.n22169 vss.n22168 1.991
R18542 vss.n21531 vss.n21521 1.991
R18543 vss.n21523 vss.n21522 1.991
R18544 vss.n21504 vss.n21503 1.991
R18545 vss.n21513 vss.n21512 1.991
R18546 vss.n21323 vss.n21313 1.991
R18547 vss.n21315 vss.n21314 1.991
R18548 vss.n21296 vss.n21295 1.991
R18549 vss.n21305 vss.n21304 1.991
R18550 vss.n21115 vss.n21105 1.991
R18551 vss.n21107 vss.n21106 1.991
R18552 vss.n21088 vss.n21087 1.991
R18553 vss.n21097 vss.n21096 1.991
R18554 vss.n20907 vss.n20897 1.991
R18555 vss.n20899 vss.n20898 1.991
R18556 vss.n8766 vss.n8756 1.991
R18557 vss.n8758 vss.n8757 1.991
R18558 vss.n8739 vss.n8738 1.991
R18559 vss.n8748 vss.n8747 1.991
R18560 vss.n8558 vss.n8548 1.991
R18561 vss.n8550 vss.n8549 1.991
R18562 vss.n8531 vss.n8530 1.991
R18563 vss.n8540 vss.n8539 1.991
R18564 vss.n8350 vss.n8340 1.991
R18565 vss.n8342 vss.n8341 1.991
R18566 vss.n8323 vss.n8322 1.991
R18567 vss.n8332 vss.n8331 1.991
R18568 vss.n8142 vss.n8132 1.991
R18569 vss.n8134 vss.n8133 1.991
R18570 vss.n8115 vss.n8114 1.991
R18571 vss.n8124 vss.n8123 1.991
R18572 vss.n7934 vss.n7924 1.991
R18573 vss.n7926 vss.n7925 1.991
R18574 vss.n7907 vss.n7906 1.991
R18575 vss.n7916 vss.n7915 1.991
R18576 vss.n7725 vss.n7715 1.991
R18577 vss.n7717 vss.n7716 1.991
R18578 vss.n7698 vss.n7697 1.991
R18579 vss.n7707 vss.n7706 1.991
R18580 vss.n7517 vss.n7507 1.991
R18581 vss.n7509 vss.n7508 1.991
R18582 vss.n18957 vss.n17681 1.97
R18583 vss.n18942 vss.n17688 1.97
R18584 vss.n17786 vss.n17780 1.97
R18585 vss.n17799 vss.n17790 1.97
R18586 vss.n18713 vss.n17887 1.97
R18587 vss.n18701 vss.n17900 1.97
R18588 vss.n17999 vss.n17993 1.97
R18589 vss.n18012 vss.n18003 1.97
R18590 vss.n18472 vss.n18100 1.97
R18591 vss.n18460 vss.n18113 1.97
R18592 vss.n18212 vss.n18206 1.97
R18593 vss.n18225 vss.n18216 1.97
R18594 vss.n19086 vss.n19080 1.97
R18595 vss.n19099 vss.n19090 1.97
R18596 vss.n20103 vss.n19188 1.97
R18597 vss.n20088 vss.n19195 1.97
R18598 vss.n19293 vss.n19287 1.97
R18599 vss.n19306 vss.n19297 1.97
R18600 vss.n19856 vss.n19395 1.97
R18601 vss.n19841 vss.n19401 1.97
R18602 vss.n19500 vss.n19494 1.97
R18603 vss.n19513 vss.n19504 1.97
R18604 vss.n19610 vss.n17592 1.97
R18605 vss.n5567 vss.n4291 1.97
R18606 vss.n5552 vss.n4298 1.97
R18607 vss.n4396 vss.n4390 1.97
R18608 vss.n4409 vss.n4400 1.97
R18609 vss.n5323 vss.n4497 1.97
R18610 vss.n5311 vss.n4510 1.97
R18611 vss.n4609 vss.n4603 1.97
R18612 vss.n4622 vss.n4613 1.97
R18613 vss.n5082 vss.n4710 1.97
R18614 vss.n5070 vss.n4723 1.97
R18615 vss.n4822 vss.n4816 1.97
R18616 vss.n4835 vss.n4826 1.97
R18617 vss.n5696 vss.n5690 1.97
R18618 vss.n5709 vss.n5700 1.97
R18619 vss.n6713 vss.n5798 1.97
R18620 vss.n6698 vss.n5805 1.97
R18621 vss.n5903 vss.n5897 1.97
R18622 vss.n5916 vss.n5907 1.97
R18623 vss.n6466 vss.n6005 1.97
R18624 vss.n6451 vss.n6011 1.97
R18625 vss.n6110 vss.n6104 1.97
R18626 vss.n6123 vss.n6114 1.97
R18627 vss.n6220 vss.n4202 1.97
R18628 vss.n16772 vss.n16771 1.97
R18629 vss.n16790 vss.n16789 1.97
R18630 vss.n17004 vss.n17003 1.97
R18631 vss.n17021 vss.n17020 1.97
R18632 vss.n17240 vss.n17239 1.97
R18633 vss.n17259 vss.n17258 1.97
R18634 vss.n16053 vss.n16050 1.97
R18635 vss.n16069 vss.n16066 1.97
R18636 vss.n16245 vss.n16244 1.97
R18637 vss.n15231 vss.n15230 1.97
R18638 vss.n15316 vss.n15315 1.97
R18639 vss.n15524 vss.n15523 1.97
R18640 vss.n15541 vss.n15540 1.97
R18641 vss.n15760 vss.n15759 1.97
R18642 vss.n15775 vss.n15774 1.97
R18643 vss.n16471 vss.n16470 1.97
R18644 vss.n16488 vss.n16487 1.97
R18645 vss.n16668 vss.n16667 1.97
R18646 vss.n9109 vss.n9108 1.969
R18647 vss.n21833 vss.n21832 1.965
R18648 vss.n21840 vss.n21839 1.965
R18649 vss.n21727 vss.n21726 1.965
R18650 vss.n21734 vss.n21732 1.965
R18651 vss.n3782 vss.n3781 1.965
R18652 vss.n3789 vss.n3788 1.965
R18653 vss.n3676 vss.n3675 1.965
R18654 vss.n3683 vss.n3681 1.965
R18655 vss.n9646 vss.n9645 1.957
R18656 vss.n15003 vss.n14999 1.95
R18657 vss.n13961 vss.n13957 1.95
R18658 vss.n11814 vss.n11810 1.95
R18659 vss.n14575 vss.n14571 1.95
R18660 vss.n13635 vss.n13631 1.95
R18661 vss.n13687 vss.n13683 1.95
R18662 vss.n11384 vss.n11380 1.95
R18663 vss.n11370 vss.n11366 1.95
R18664 vss.n11313 vss.n11309 1.95
R18665 vss.n12401 vss.n12397 1.95
R18666 vss.n14711 vss.n14707 1.95
R18667 vss.n13448 vss.n13444 1.95
R18668 vss.n13023 vss.n13019 1.95
R18669 vss.n10580 vss.n10576 1.95
R18670 vss.n10737 vss.n10733 1.95
R18671 vss.n12033 vss.n12029 1.95
R18672 vss.n10250 vss.n10249 1.94
R18673 vss.n10354 vss.n10353 1.94
R18674 vss.n17339 vss.n17335 1.931
R18675 vss.n17350 vss.n17346 1.931
R18676 vss.n17361 vss.n17357 1.931
R18677 vss.n17372 vss.n17368 1.931
R18678 vss.n17383 vss.n17379 1.931
R18679 vss.n17394 vss.n17390 1.931
R18680 vss.n17416 vss.n17412 1.931
R18681 vss.n17427 vss.n17423 1.931
R18682 vss.n17438 vss.n17434 1.931
R18683 vss.n17449 vss.n17445 1.931
R18684 vss.n17460 vss.n17456 1.931
R18685 vss.n17471 vss.n17467 1.931
R18686 vss.n17482 vss.n17478 1.931
R18687 vss.n3497 vss.n3493 1.931
R18688 vss.n3508 vss.n3504 1.931
R18689 vss.n3519 vss.n3515 1.931
R18690 vss.n3530 vss.n3526 1.931
R18691 vss.n3541 vss.n3537 1.931
R18692 vss.n3552 vss.n3548 1.931
R18693 vss.n4026 vss.n4022 1.931
R18694 vss.n4037 vss.n4033 1.931
R18695 vss.n4048 vss.n4044 1.931
R18696 vss.n4059 vss.n4055 1.931
R18697 vss.n4070 vss.n4066 1.931
R18698 vss.n4081 vss.n4077 1.931
R18699 vss.n4092 vss.n4088 1.931
R18700 vss.n21945 vss.n21943 1.925
R18701 vss.n3894 vss.n3892 1.925
R18702 vss.n16350 vss.n16349 1.92
R18703 vss.n16371 vss.n16370 1.92
R18704 vss.n16586 vss.n16585 1.92
R18705 vss.n16607 vss.n16606 1.92
R18706 vss.n16664 vss.n16662 1.92
R18707 vss.n16889 vss.n16888 1.92
R18708 vss.n16904 vss.n16903 1.92
R18709 vss.n17011 vss.n17010 1.92
R18710 vss.n17042 vss.n17033 1.92
R18711 vss.n17125 vss.n17124 1.92
R18712 vss.n17140 vss.n17139 1.92
R18713 vss.n17247 vss.n17246 1.92
R18714 vss.n15927 vss.n15926 1.92
R18715 vss.n15951 vss.n15950 1.92
R18716 vss.n16058 vss.n16056 1.92
R18717 vss.n16087 vss.n16086 1.92
R18718 vss.n16163 vss.n16162 1.92
R18719 vss.n16187 vss.n16186 1.92
R18720 vss.n16295 vss.n16294 1.92
R18721 vss.n15403 vss.n15402 1.92
R18722 vss.n15424 vss.n15423 1.92
R18723 vss.n15639 vss.n15638 1.92
R18724 vss.n15660 vss.n15659 1.92
R18725 vss.n15874 vss.n15873 1.92
R18726 vss.n13135 vss.n13134 1.914
R18727 vss.n13676 vss.n13675 1.914
R18728 vss.n13126 vss.n13125 1.914
R18729 vss.n11468 vss.n11467 1.914
R18730 vss.n10663 vss.n10662 1.914
R18731 vss.n11460 vss.n11459 1.914
R18732 vss.n10655 vss.n10654 1.914
R18733 vss.n13644 vss.n13643 1.914
R18734 vss.n15249 vss.n15248 1.914
R18735 vss.n13222 vss.n13221 1.9
R18736 vss.n14271 vss.n14270 1.9
R18737 vss.n11036 vss.n11035 1.9
R18738 vss.n12522 vss.n12521 1.9
R18739 vss.n16258 vss.n16257 1.9
R18740 vss.n14497 vss.n14496 1.894
R18741 vss.n14666 vss.n14665 1.894
R18742 vss.n13584 vss.n13574 1.894
R18743 vss.n13343 vss.n13333 1.894
R18744 vss.n10510 vss.n10500 1.894
R18745 vss.n14363 vss.n14362 1.894
R18746 vss.n13867 vss.n13857 1.894
R18747 vss.n11766 vss.n11765 1.894
R18748 vss.n13982 vss.n13972 1.894
R18749 vss.n11577 vss.n11567 1.894
R18750 vss.n12085 vss.n12084 1.894
R18751 vss.n10829 vss.n10828 1.894
R18752 vss.n10903 vss.n10902 1.894
R18753 vss.n10955 vss.n10945 1.894
R18754 vss.n11017 vss.n11016 1.894
R18755 vss.n20453 vss.n20445 1.882
R18756 vss.n20635 vss.n20627 1.882
R18757 vss.n20683 vss.n20675 1.882
R18758 vss.n20859 vss.n20851 1.882
R18759 vss.n21666 vss.n21660 1.882
R18760 vss.n21666 vss.n21659 1.882
R18761 vss.n21798 vss.n21643 1.882
R18762 vss.n12228 vss.n12221 1.882
R18763 vss.n12022 vss.n12015 1.882
R18764 vss.n11258 vss.n11251 1.882
R18765 vss.n11198 vss.n11191 1.882
R18766 vss.n13915 vss.n13908 1.882
R18767 vss.n14053 vss.n14046 1.882
R18768 vss.n11748 vss.n11741 1.882
R18769 vss.n11075 vss.n11068 1.882
R18770 vss.n14742 vss.n14735 1.882
R18771 vss.n14683 vss.n14676 1.882
R18772 vss.n14470 vss.n14463 1.882
R18773 vss.n14252 vss.n14245 1.882
R18774 vss.n12858 vss.n12857 1.882
R18775 vss.n12857 vss.n12850 1.882
R18776 vss.n12658 vss.n12657 1.882
R18777 vss.n12657 vss.n12650 1.882
R18778 vss.n3615 vss.n3609 1.882
R18779 vss.n3615 vss.n3608 1.882
R18780 vss.n3747 vss.n3592 1.882
R18781 vss.n7063 vss.n7055 1.882
R18782 vss.n7245 vss.n7237 1.882
R18783 vss.n7293 vss.n7285 1.882
R18784 vss.n7469 vss.n7461 1.882
R18785 vss.n1856 vss.n1848 1.882
R18786 vss.n1906 vss.n1897 1.882
R18787 vss.n2099 vss.n2090 1.882
R18788 vss.n2150 vss.n2141 1.882
R18789 vss.n2344 vss.n2335 1.882
R18790 vss.n2394 vss.n2385 1.882
R18791 vss.n2588 vss.n2579 1.882
R18792 vss.n2639 vss.n2630 1.882
R18793 vss.n2830 vss.n2822 1.882
R18794 vss.n2877 vss.n2868 1.882
R18795 vss.n3071 vss.n3062 1.882
R18796 vss.n3122 vss.n3113 1.882
R18797 vss.n3315 vss.n3306 1.882
R18798 vss.n3364 vss.n3356 1.882
R18799 vss.n317 vss.n309 1.882
R18800 vss.n367 vss.n358 1.882
R18801 vss.n560 vss.n551 1.882
R18802 vss.n611 vss.n602 1.882
R18803 vss.n805 vss.n796 1.882
R18804 vss.n855 vss.n846 1.882
R18805 vss.n1049 vss.n1040 1.882
R18806 vss.n1100 vss.n1091 1.882
R18807 vss.n1294 vss.n1285 1.882
R18808 vss.n23388 vss.n23379 1.882
R18809 vss.n23195 vss.n23186 1.882
R18810 vss.n23144 vss.n23135 1.882
R18811 vss.n22951 vss.n22942 1.882
R18812 vss.n22901 vss.n22893 1.882
R18813 vss.n20367 vss.n17582 1.866
R18814 vss.n6977 vss.n4192 1.866
R18815 vss.n21972 vss.n21971 1.864
R18816 vss.n21609 vss.n21608 1.864
R18817 vss.n3921 vss.n3920 1.864
R18818 vss.n3558 vss.n3557 1.864
R18819 vss.n22721 vss.n22714 1.848
R18820 vss.n22723 vss.n22721 1.848
R18821 vss.n22673 vss.n22672 1.848
R18822 vss.n22672 vss.n22665 1.848
R18823 vss.n22513 vss.n22506 1.848
R18824 vss.n22515 vss.n22513 1.848
R18825 vss.n22465 vss.n22464 1.848
R18826 vss.n22464 vss.n22457 1.848
R18827 vss.n22305 vss.n22298 1.848
R18828 vss.n22307 vss.n22305 1.848
R18829 vss.n22257 vss.n22256 1.848
R18830 vss.n22256 vss.n22249 1.848
R18831 vss.n22097 vss.n22090 1.848
R18832 vss.n22099 vss.n22097 1.848
R18833 vss.n21589 vss.n21588 1.848
R18834 vss.n21588 vss.n21581 1.848
R18835 vss.n21441 vss.n21434 1.848
R18836 vss.n21443 vss.n21441 1.848
R18837 vss.n21393 vss.n21392 1.848
R18838 vss.n21392 vss.n21385 1.848
R18839 vss.n21233 vss.n21226 1.848
R18840 vss.n21235 vss.n21233 1.848
R18841 vss.n21185 vss.n21184 1.848
R18842 vss.n21184 vss.n21177 1.848
R18843 vss.n21025 vss.n21018 1.848
R18844 vss.n21027 vss.n21025 1.848
R18845 vss.n20977 vss.n20976 1.848
R18846 vss.n20976 vss.n20969 1.848
R18847 vss.n8884 vss.n8877 1.848
R18848 vss.n8886 vss.n8884 1.848
R18849 vss.n8836 vss.n8835 1.848
R18850 vss.n8835 vss.n8828 1.848
R18851 vss.n8676 vss.n8669 1.848
R18852 vss.n8678 vss.n8676 1.848
R18853 vss.n8628 vss.n8627 1.848
R18854 vss.n8627 vss.n8620 1.848
R18855 vss.n8468 vss.n8461 1.848
R18856 vss.n8470 vss.n8468 1.848
R18857 vss.n8420 vss.n8419 1.848
R18858 vss.n8419 vss.n8412 1.848
R18859 vss.n8260 vss.n8253 1.848
R18860 vss.n8262 vss.n8260 1.848
R18861 vss.n8212 vss.n8211 1.848
R18862 vss.n8211 vss.n8204 1.848
R18863 vss.n8052 vss.n8045 1.848
R18864 vss.n8054 vss.n8052 1.848
R18865 vss.n8004 vss.n8003 1.848
R18866 vss.n8003 vss.n7996 1.848
R18867 vss.n7843 vss.n7836 1.848
R18868 vss.n7845 vss.n7843 1.848
R18869 vss.n7795 vss.n7794 1.848
R18870 vss.n7794 vss.n7787 1.848
R18871 vss.n7635 vss.n7628 1.848
R18872 vss.n7637 vss.n7635 1.848
R18873 vss.n7587 vss.n7586 1.848
R18874 vss.n7586 vss.n7579 1.848
R18875 vss.n11066 vss.n11065 1.839
R18876 vss.n14233 vss.n14232 1.839
R18877 vss.n20405 vss.n17556 1.836
R18878 vss.n7015 vss.n4166 1.836
R18879 vss.n21658 vss.n21651 1.82
R18880 vss.n3607 vss.n3600 1.82
R18881 vss.n16462 vss.n16455 1.792
R18882 vss.n16509 vss.n16502 1.792
R18883 vss.n16696 vss.n16695 1.792
R18884 vss.n16765 vss.n16758 1.792
R18885 vss.n16806 vss.n16799 1.792
R18886 vss.n16881 vss.n16880 1.792
R18887 vss.n16926 vss.n16925 1.792
R18888 vss.n16997 vss.n16988 1.792
R18889 vss.n17042 vss.n17041 1.792
R18890 vss.n17117 vss.n17116 1.792
R18891 vss.n17162 vss.n17161 1.792
R18892 vss.n17233 vss.n17224 1.792
R18893 vss.n17295 vss.n17288 1.792
R18894 vss.n15935 vss.n15925 1.792
R18895 vss.n15974 vss.n15973 1.792
R18896 vss.n16042 vss.n16035 1.792
R18897 vss.n16086 vss.n16079 1.792
R18898 vss.n16171 vss.n16161 1.792
R18899 vss.n16210 vss.n16209 1.792
R18900 vss.n15248 vss.n15241 1.792
R18901 vss.n15226 vss.n15219 1.792
R18902 vss.n15515 vss.n15508 1.792
R18903 vss.n15562 vss.n15555 1.792
R18904 vss.n15751 vss.n15744 1.792
R18905 vss.n15792 vss.n15785 1.792
R18906 vss.n16256 vss.n16255 1.774
R18907 vss.n14643 vss.n14642 1.76
R18908 vss.n13564 vss.n13554 1.76
R18909 vss.n10480 vss.n10470 1.76
R18910 vss.n14003 vss.n13993 1.76
R18911 vss.n11595 vss.n11585 1.76
R18912 vss.n10848 vss.n10838 1.76
R18913 vss.n10892 vss.n10882 1.76
R18914 vss.n16672 vss.n16668 1.732
R18915 vss.n16249 vss.n16245 1.732
R18916 vss.n17329 vss.n17328 1.728
R18917 vss.n8999 vss.n8998 1.724
R18918 vss.n22617 vss.n22607 1.706
R18919 vss.n22609 vss.n22608 1.706
R18920 vss.n22562 vss.n22561 1.706
R18921 vss.n22571 vss.n22570 1.706
R18922 vss.n22409 vss.n22399 1.706
R18923 vss.n22401 vss.n22400 1.706
R18924 vss.n22354 vss.n22353 1.706
R18925 vss.n22363 vss.n22362 1.706
R18926 vss.n22201 vss.n22191 1.706
R18927 vss.n22193 vss.n22192 1.706
R18928 vss.n22146 vss.n22145 1.706
R18929 vss.n22155 vss.n22154 1.706
R18930 vss.n21545 vss.n21535 1.706
R18931 vss.n21537 vss.n21536 1.706
R18932 vss.n21490 vss.n21489 1.706
R18933 vss.n21499 vss.n21498 1.706
R18934 vss.n21337 vss.n21327 1.706
R18935 vss.n21329 vss.n21328 1.706
R18936 vss.n21282 vss.n21281 1.706
R18937 vss.n21291 vss.n21290 1.706
R18938 vss.n21129 vss.n21119 1.706
R18939 vss.n21121 vss.n21120 1.706
R18940 vss.n21074 vss.n21073 1.706
R18941 vss.n21083 vss.n21082 1.706
R18942 vss.n20921 vss.n20911 1.706
R18943 vss.n20913 vss.n20912 1.706
R18944 vss.n8780 vss.n8770 1.706
R18945 vss.n8772 vss.n8771 1.706
R18946 vss.n8725 vss.n8724 1.706
R18947 vss.n8734 vss.n8733 1.706
R18948 vss.n8572 vss.n8562 1.706
R18949 vss.n8564 vss.n8563 1.706
R18950 vss.n8517 vss.n8516 1.706
R18951 vss.n8526 vss.n8525 1.706
R18952 vss.n8364 vss.n8354 1.706
R18953 vss.n8356 vss.n8355 1.706
R18954 vss.n8309 vss.n8308 1.706
R18955 vss.n8318 vss.n8317 1.706
R18956 vss.n8156 vss.n8146 1.706
R18957 vss.n8148 vss.n8147 1.706
R18958 vss.n8101 vss.n8100 1.706
R18959 vss.n8110 vss.n8109 1.706
R18960 vss.n7948 vss.n7938 1.706
R18961 vss.n7940 vss.n7939 1.706
R18962 vss.n7893 vss.n7892 1.706
R18963 vss.n7902 vss.n7901 1.706
R18964 vss.n7739 vss.n7729 1.706
R18965 vss.n7731 vss.n7730 1.706
R18966 vss.n7684 vss.n7683 1.706
R18967 vss.n7693 vss.n7692 1.706
R18968 vss.n7531 vss.n7521 1.706
R18969 vss.n7523 vss.n7522 1.706
R18970 vss.n19605 vss.n19604 1.688
R18971 vss.n6215 vss.n6214 1.688
R18972 vss.n13765 vss.n13763 1.666
R18973 vss.n14136 vss.n14135 1.666
R18974 vss.n10993 vss.n10991 1.666
R18975 vss.n11537 vss.n11536 1.666
R18976 vss.n11964 vss.n11962 1.666
R18977 vss.n11890 vss.n11888 1.666
R18978 vss.n10718 vss.n10717 1.666
R18979 vss.n12277 vss.n12275 1.666
R18980 vss.n12092 vss.n12090 1.666
R18981 vss.n12377 vss.n12376 1.666
R18982 vss.n12341 vss.n12339 1.666
R18983 vss.n10617 vss.n10615 1.666
R18984 vss.n13179 vss.n13178 1.666
R18985 vss.n10467 vss.n10465 1.666
R18986 vss.n12938 vss.n12937 1.666
R18987 vss.n12969 vss.n12968 1.666
R18988 vss.n13552 vss.n13550 1.666
R18989 vss.n13008 vss.n13007 1.666
R18990 vss.n10608 vss.n10606 1.666
R18991 vss.n10556 vss.n10555 1.666
R18992 vss.n11414 vss.n11412 1.666
R18993 vss.n11501 vss.n11500 1.666
R18994 vss.n16336 vss.n16335 1.664
R18995 vss.n16385 vss.n16384 1.664
R18996 vss.n16572 vss.n16571 1.664
R18997 vss.n16621 vss.n16620 1.664
R18998 vss.n16688 vss.n16687 1.664
R18999 vss.n16820 vss.n16811 1.664
R19000 vss.n16875 vss.n16874 1.664
R19001 vss.n16918 vss.n16917 1.664
R19002 vss.n16997 vss.n16996 1.664
R19003 vss.n17056 vss.n17047 1.664
R19004 vss.n17111 vss.n17110 1.664
R19005 vss.n17154 vss.n17153 1.664
R19006 vss.n17233 vss.n17232 1.664
R19007 vss.n15913 vss.n15912 1.664
R19008 vss.n15965 vss.n15964 1.664
R19009 vss.n16044 vss.n16042 1.664
R19010 vss.n16101 vss.n16100 1.664
R19011 vss.n16149 vss.n16148 1.664
R19012 vss.n16201 vss.n16200 1.664
R19013 vss.n16274 vss.n16273 1.664
R19014 vss.n15389 vss.n15388 1.664
R19015 vss.n15438 vss.n15437 1.664
R19016 vss.n15625 vss.n15624 1.664
R19017 vss.n15674 vss.n15673 1.664
R19018 vss.n15853 vss.n15852 1.664
R19019 vss.n14487 vss.n14486 1.647
R19020 vss.n14394 vss.n14393 1.647
R19021 vss.n14657 vss.n14656 1.647
R19022 vss.n13576 vss.n13575 1.647
R19023 vss.n13294 vss.n13293 1.647
R19024 vss.n13335 vss.n13334 1.647
R19025 vss.n10502 vss.n10501 1.647
R19026 vss.n14353 vss.n14352 1.647
R19027 vss.n13859 vss.n13858 1.647
R19028 vss.n11756 vss.n11755 1.647
R19029 vss.n11046 vss.n11045 1.647
R19030 vss.n13974 vss.n13973 1.647
R19031 vss.n11569 vss.n11568 1.647
R19032 vss.n12579 vss.n12578 1.647
R19033 vss.n12075 vss.n12074 1.647
R19034 vss.n12421 vss.n12420 1.647
R19035 vss.n10820 vss.n10819 1.647
R19036 vss.n10894 vss.n10893 1.647
R19037 vss.n10947 vss.n10946 1.647
R19038 vss.n11007 vss.n11006 1.647
R19039 vss.n17273 vss.n17272 1.647
R19040 vss.n15817 vss.t229 1.641
R19041 vss.n15211 vss.t310 1.64
R19042 vss.n20407 vss.n17549 1.618
R19043 vss.n7017 vss.n4159 1.618
R19044 vss.n9154 vss.n9153 1.603
R19045 vss.n21992 vss.n21991 1.601
R19046 vss.n21789 vss.n21696 1.601
R19047 vss.n21796 vss.n21663 1.601
R19048 vss.n3941 vss.n3940 1.601
R19049 vss.n3738 vss.n3645 1.601
R19050 vss.n3745 vss.n3612 1.601
R19051 vss.n21996 vss.n21995 1.601
R19052 vss.n3945 vss.n3944 1.601
R19053 vss.n13804 vss.n13803 1.577
R19054 vss.n14761 vss.n14760 1.577
R19055 vss.n14436 vss.n14435 1.573
R19056 vss.t2 vss.n10184 1.569
R19057 vss.n10418 vss.n10395 1.567
R19058 vss.n22735 vss.n22728 1.564
R19059 vss.n22737 vss.n22735 1.564
R19060 vss.n22659 vss.n22658 1.564
R19061 vss.n22658 vss.n22651 1.564
R19062 vss.n22527 vss.n22520 1.564
R19063 vss.n22529 vss.n22527 1.564
R19064 vss.n22451 vss.n22450 1.564
R19065 vss.n22450 vss.n22443 1.564
R19066 vss.n22319 vss.n22312 1.564
R19067 vss.n22321 vss.n22319 1.564
R19068 vss.n22243 vss.n22242 1.564
R19069 vss.n22242 vss.n22235 1.564
R19070 vss.n22111 vss.n22104 1.564
R19071 vss.n22113 vss.n22111 1.564
R19072 vss.n17408 vss.n17407 1.564
R19073 vss.n17407 vss.n17400 1.564
R19074 vss.n21455 vss.n21448 1.564
R19075 vss.n21457 vss.n21455 1.564
R19076 vss.n21379 vss.n21378 1.564
R19077 vss.n21378 vss.n21371 1.564
R19078 vss.n21247 vss.n21240 1.564
R19079 vss.n21249 vss.n21247 1.564
R19080 vss.n21171 vss.n21170 1.564
R19081 vss.n21170 vss.n21163 1.564
R19082 vss.n21039 vss.n21032 1.564
R19083 vss.n21041 vss.n21039 1.564
R19084 vss.n20963 vss.n20962 1.564
R19085 vss.n20962 vss.n20955 1.564
R19086 vss.n8898 vss.n8891 1.564
R19087 vss.n8900 vss.n8898 1.564
R19088 vss.n8822 vss.n8821 1.564
R19089 vss.n8821 vss.n8814 1.564
R19090 vss.n8690 vss.n8683 1.564
R19091 vss.n8692 vss.n8690 1.564
R19092 vss.n8614 vss.n8613 1.564
R19093 vss.n8613 vss.n8606 1.564
R19094 vss.n8482 vss.n8475 1.564
R19095 vss.n8484 vss.n8482 1.564
R19096 vss.n8406 vss.n8405 1.564
R19097 vss.n8405 vss.n8398 1.564
R19098 vss.n8274 vss.n8267 1.564
R19099 vss.n8276 vss.n8274 1.564
R19100 vss.n8198 vss.n8197 1.564
R19101 vss.n8197 vss.n8190 1.564
R19102 vss.n8066 vss.n8059 1.564
R19103 vss.n8068 vss.n8066 1.564
R19104 vss.n7990 vss.n7989 1.564
R19105 vss.n7989 vss.n7982 1.564
R19106 vss.n7858 vss.n7851 1.564
R19107 vss.n7860 vss.n7858 1.564
R19108 vss.n7781 vss.n7780 1.564
R19109 vss.n7780 vss.n7773 1.564
R19110 vss.n7649 vss.n7642 1.564
R19111 vss.n7651 vss.n7649 1.564
R19112 vss.n7573 vss.n7572 1.564
R19113 vss.n7572 vss.n7565 1.564
R19114 vss.n16448 vss.n16441 1.536
R19115 vss.n16523 vss.n16516 1.536
R19116 vss.n16710 vss.n16709 1.536
R19117 vss.n16753 vss.n16744 1.536
R19118 vss.n16820 vss.n16813 1.536
R19119 vss.n16867 vss.n16866 1.536
R19120 vss.n16940 vss.n16939 1.536
R19121 vss.n16983 vss.n16974 1.536
R19122 vss.n17056 vss.n17055 1.536
R19123 vss.n17103 vss.n17102 1.536
R19124 vss.n17176 vss.n17175 1.536
R19125 vss.n17219 vss.n17210 1.536
R19126 vss.n17305 vss.n17298 1.536
R19127 vss.n15921 vss.n15911 1.536
R19128 vss.n15988 vss.n15987 1.536
R19129 vss.n16028 vss.n16021 1.536
R19130 vss.n16100 vss.n16093 1.536
R19131 vss.n16157 vss.n16147 1.536
R19132 vss.n16224 vss.n16223 1.536
R19133 vss.n15300 vss.n15293 1.536
R19134 vss.n15339 vss.n15332 1.536
R19135 vss.n15501 vss.n15494 1.536
R19136 vss.n15576 vss.n15569 1.536
R19137 vss.n15737 vss.n15730 1.536
R19138 vss.n15804 vss.n15797 1.536
R19139 vss.n10301 vss.n10300 1.533
R19140 vss.n10360 vss.n10359 1.533
R19141 vss.n22050 vss.n22049 1.525
R19142 vss.n3999 vss.n3998 1.525
R19143 vss.n21760 vss.n21701 1.525
R19144 vss.n3709 vss.n3650 1.525
R19145 vss.n21906 vss.n21905 1.511
R19146 vss.n3855 vss.n3854 1.511
R19147 vss.n20507 vss.n20506 1.505
R19148 vss.n20567 vss.n20566 1.505
R19149 vss.n20735 vss.n20734 1.505
R19150 vss.n20789 vss.n20788 1.505
R19151 vss.n21805 vss.n21804 1.505
R19152 vss.n21667 vss.n21648 1.505
R19153 vss.n12138 vss.n12137 1.505
R19154 vss.n11970 vss.n11969 1.505
R19155 vss.n11916 vss.n11915 1.505
R19156 vss.n14332 vss.n14331 1.505
R19157 vss.n11620 vss.n11619 1.505
R19158 vss.n11669 vss.n11668 1.505
R19159 vss.n14810 vss.n14809 1.505
R19160 vss.n14609 vss.n14608 1.505
R19161 vss.n14549 vss.n14548 1.505
R19162 vss.n14910 vss.n14909 1.505
R19163 vss.n14900 vss.n14899 1.505
R19164 vss.n10459 vss.n10458 1.505
R19165 vss.n10542 vss.n10541 1.505
R19166 vss.n3754 vss.n3753 1.505
R19167 vss.n3616 vss.n3597 1.505
R19168 vss.n7117 vss.n7116 1.505
R19169 vss.n7177 vss.n7176 1.505
R19170 vss.n7345 vss.n7344 1.505
R19171 vss.n7399 vss.n7398 1.505
R19172 vss.n1729 vss.n1728 1.505
R19173 vss.n1788 vss.n1787 1.505
R19174 vss.n1961 vss.n1960 1.505
R19175 vss.n2026 vss.n2025 1.505
R19176 vss.n2206 vss.n2205 1.505
R19177 vss.n2270 vss.n2269 1.505
R19178 vss.n2450 vss.n2449 1.505
R19179 vss.n2515 vss.n2514 1.505
R19180 vss.n2694 vss.n2693 1.505
R19181 vss.n2759 vss.n2758 1.505
R19182 vss.n2933 vss.n2932 1.505
R19183 vss.n2997 vss.n2996 1.505
R19184 vss.n3177 vss.n3176 1.505
R19185 vss.n3242 vss.n3241 1.505
R19186 vss.n3416 vss.n3415 1.505
R19187 vss.n3457 vss.n3456 1.505
R19188 vss.n190 vss.n189 1.505
R19189 vss.n249 vss.n248 1.505
R19190 vss.n422 vss.n421 1.505
R19191 vss.n487 vss.n486 1.505
R19192 vss.n667 vss.n666 1.505
R19193 vss.n731 vss.n730 1.505
R19194 vss.n911 vss.n910 1.505
R19195 vss.n976 vss.n975 1.505
R19196 vss.n1155 vss.n1154 1.505
R19197 vss.n1220 vss.n1219 1.505
R19198 vss.n23315 vss.n23314 1.505
R19199 vss.n23251 vss.n23250 1.505
R19200 vss.n23071 vss.n23070 1.505
R19201 vss.n23006 vss.n23005 1.505
R19202 vss.n22831 vss.n22830 1.505
R19203 vss.n1432 vss.n1431 1.505
R19204 vss.n21953 vss.n21952 1.5
R19205 vss.n3902 vss.n3901 1.5
R19206 vss.n17585 vss.n17584 1.5
R19207 vss.n20364 vss.n20363 1.5
R19208 vss.n20372 vss.n17577 1.5
R19209 vss.n21758 vss.n21700 1.5
R19210 vss.n10418 vss.n10417 1.5
R19211 vss.n3707 vss.n3649 1.5
R19212 vss.n4195 vss.n4194 1.5
R19213 vss.n6974 vss.n6973 1.5
R19214 vss.n6982 vss.n4187 1.5
R19215 vss.n21926 vss.n21925 1.497
R19216 vss.n3875 vss.n3874 1.497
R19217 vss.n13890 vss.n13889 1.49
R19218 vss.n11106 vss.n11105 1.49
R19219 vss.n11896 vss.n11895 1.49
R19220 vss.n10775 vss.n10774 1.49
R19221 vss.n12626 vss.n12625 1.49
R19222 vss.n14934 vss.n14933 1.49
R19223 vss.n13403 vss.n13402 1.49
R19224 vss.n14128 vss.n14127 1.49
R19225 vss.n13475 vss.n13474 1.49
R19226 vss.n11421 vss.n11420 1.49
R19227 vss.n11601 vss.n11600 1.49
R19228 vss.n9647 vss.n9159 1.473
R19229 vss.n17331 ldomc_0.vss 1.472
R19230 vss.n18952 vss.n18951 1.466
R19231 vss.n18947 vss.n17685 1.466
R19232 vss.n18831 vss.n17785 1.466
R19233 vss.n18825 vss.n17792 1.466
R19234 vss.n18711 vss.n17892 1.466
R19235 vss.n18706 vss.n17895 1.466
R19236 vss.n18590 vss.n17998 1.466
R19237 vss.n18584 vss.n18005 1.466
R19238 vss.n18470 vss.n18105 1.466
R19239 vss.n18465 vss.n18108 1.466
R19240 vss.n18349 vss.n18211 1.466
R19241 vss.n18343 vss.n18218 1.466
R19242 vss.n20224 vss.n19085 1.466
R19243 vss.n20218 vss.n19092 1.466
R19244 vss.n20098 vss.n20097 1.466
R19245 vss.n20093 vss.n19192 1.466
R19246 vss.n19977 vss.n19292 1.466
R19247 vss.n19971 vss.n19299 1.466
R19248 vss.n19851 vss.n19850 1.466
R19249 vss.n19846 vss.n19398 1.466
R19250 vss.n19730 vss.n19499 1.466
R19251 vss.n19724 vss.n19506 1.466
R19252 vss.n5562 vss.n5561 1.466
R19253 vss.n5557 vss.n4295 1.466
R19254 vss.n5441 vss.n4395 1.466
R19255 vss.n5435 vss.n4402 1.466
R19256 vss.n5321 vss.n4502 1.466
R19257 vss.n5316 vss.n4505 1.466
R19258 vss.n5200 vss.n4608 1.466
R19259 vss.n5194 vss.n4615 1.466
R19260 vss.n5080 vss.n4715 1.466
R19261 vss.n5075 vss.n4718 1.466
R19262 vss.n4959 vss.n4821 1.466
R19263 vss.n4953 vss.n4828 1.466
R19264 vss.n6834 vss.n5695 1.466
R19265 vss.n6828 vss.n5702 1.466
R19266 vss.n6708 vss.n6707 1.466
R19267 vss.n6703 vss.n5802 1.466
R19268 vss.n6587 vss.n5902 1.466
R19269 vss.n6581 vss.n5909 1.466
R19270 vss.n6461 vss.n6460 1.466
R19271 vss.n6456 vss.n6008 1.466
R19272 vss.n6340 vss.n6109 1.466
R19273 vss.n6334 vss.n6116 1.466
R19274 vss.n22631 vss.n22621 1.422
R19275 vss.n22623 vss.n22622 1.422
R19276 vss.n22548 vss.n22547 1.422
R19277 vss.n22557 vss.n22556 1.422
R19278 vss.n22423 vss.n22413 1.422
R19279 vss.n22415 vss.n22414 1.422
R19280 vss.n22340 vss.n22339 1.422
R19281 vss.n22349 vss.n22348 1.422
R19282 vss.n22215 vss.n22205 1.422
R19283 vss.n22207 vss.n22206 1.422
R19284 vss.n22132 vss.n22131 1.422
R19285 vss.n22141 vss.n22140 1.422
R19286 vss.n21559 vss.n21549 1.422
R19287 vss.n21551 vss.n21550 1.422
R19288 vss.n21476 vss.n21475 1.422
R19289 vss.n21485 vss.n21484 1.422
R19290 vss.n21351 vss.n21341 1.422
R19291 vss.n21343 vss.n21342 1.422
R19292 vss.n21268 vss.n21267 1.422
R19293 vss.n21277 vss.n21276 1.422
R19294 vss.n21143 vss.n21133 1.422
R19295 vss.n21135 vss.n21134 1.422
R19296 vss.n21060 vss.n21059 1.422
R19297 vss.n21069 vss.n21068 1.422
R19298 vss.n20935 vss.n20925 1.422
R19299 vss.n20927 vss.n20926 1.422
R19300 vss.n18952 vss.n17680 1.422
R19301 vss.n18947 vss.n17687 1.422
R19302 vss.n18831 vss.n17784 1.422
R19303 vss.n18825 vss.n17793 1.422
R19304 vss.n18712 vss.n18711 1.422
R19305 vss.n18706 vss.n17897 1.422
R19306 vss.n18590 vss.n17997 1.422
R19307 vss.n18584 vss.n18006 1.422
R19308 vss.n18471 vss.n18470 1.422
R19309 vss.n18465 vss.n18110 1.422
R19310 vss.n18349 vss.n18210 1.422
R19311 vss.n18343 vss.n18219 1.422
R19312 vss.n20358 vss.n17587 1.422
R19313 vss.n20224 vss.n19084 1.422
R19314 vss.n20218 vss.n19093 1.422
R19315 vss.n20098 vss.n19187 1.422
R19316 vss.n20093 vss.n19194 1.422
R19317 vss.n19977 vss.n19291 1.422
R19318 vss.n19971 vss.n19300 1.422
R19319 vss.n19851 vss.n19394 1.422
R19320 vss.n19846 vss.n19400 1.422
R19321 vss.n19730 vss.n19498 1.422
R19322 vss.n19724 vss.n19507 1.422
R19323 vss.n5562 vss.n4290 1.422
R19324 vss.n5557 vss.n4297 1.422
R19325 vss.n5441 vss.n4394 1.422
R19326 vss.n5435 vss.n4403 1.422
R19327 vss.n5322 vss.n5321 1.422
R19328 vss.n5316 vss.n4507 1.422
R19329 vss.n5200 vss.n4607 1.422
R19330 vss.n5194 vss.n4616 1.422
R19331 vss.n5081 vss.n5080 1.422
R19332 vss.n5075 vss.n4720 1.422
R19333 vss.n4959 vss.n4820 1.422
R19334 vss.n4953 vss.n4829 1.422
R19335 vss.n6968 vss.n4197 1.422
R19336 vss.n6834 vss.n5694 1.422
R19337 vss.n6828 vss.n5703 1.422
R19338 vss.n6708 vss.n5797 1.422
R19339 vss.n6703 vss.n5804 1.422
R19340 vss.n6587 vss.n5901 1.422
R19341 vss.n6581 vss.n5910 1.422
R19342 vss.n6461 vss.n6004 1.422
R19343 vss.n6456 vss.n6010 1.422
R19344 vss.n6340 vss.n6108 1.422
R19345 vss.n6334 vss.n6117 1.422
R19346 vss.n8794 vss.n8784 1.422
R19347 vss.n8786 vss.n8785 1.422
R19348 vss.n8711 vss.n8710 1.422
R19349 vss.n8720 vss.n8719 1.422
R19350 vss.n8586 vss.n8576 1.422
R19351 vss.n8578 vss.n8577 1.422
R19352 vss.n8503 vss.n8502 1.422
R19353 vss.n8512 vss.n8511 1.422
R19354 vss.n8378 vss.n8368 1.422
R19355 vss.n8370 vss.n8369 1.422
R19356 vss.n8295 vss.n8294 1.422
R19357 vss.n8304 vss.n8303 1.422
R19358 vss.n8170 vss.n8160 1.422
R19359 vss.n8162 vss.n8161 1.422
R19360 vss.n8087 vss.n8086 1.422
R19361 vss.n8096 vss.n8095 1.422
R19362 vss.n7962 vss.n7952 1.422
R19363 vss.n7954 vss.n7953 1.422
R19364 vss.n7879 vss.n7878 1.422
R19365 vss.n7888 vss.n7887 1.422
R19366 vss.n7753 vss.n7743 1.422
R19367 vss.n7745 vss.n7744 1.422
R19368 vss.n7670 vss.n7669 1.422
R19369 vss.n7679 vss.n7678 1.422
R19370 vss.n7545 vss.n7535 1.422
R19371 vss.n7537 vss.n7536 1.422
R19372 vss.n10451 vss.n10450 1.418
R19373 vss.n13812 vss.n13811 1.411
R19374 vss.n11531 vss.n11530 1.411
R19375 vss.n12371 vss.n12370 1.411
R19376 vss.n13171 vss.n13170 1.411
R19377 vss.n10712 vss.n10711 1.411
R19378 vss.n13002 vss.n13001 1.411
R19379 vss.n12457 vss.n12456 1.409
R19380 vss.n16322 vss.n16321 1.408
R19381 vss.n16399 vss.n16398 1.408
R19382 vss.n16558 vss.n16557 1.408
R19383 vss.n16635 vss.n16634 1.408
R19384 vss.n16702 vss.n16701 1.408
R19385 vss.n16753 vss.n16752 1.408
R19386 vss.n16834 vss.n16825 1.408
R19387 vss.n16861 vss.n16860 1.408
R19388 vss.n16932 vss.n16931 1.408
R19389 vss.n16983 vss.n16982 1.408
R19390 vss.n17070 vss.n17061 1.408
R19391 vss.n17097 vss.n17096 1.408
R19392 vss.n17168 vss.n17167 1.408
R19393 vss.n17219 vss.n17218 1.408
R19394 vss.n17314 vss.n17313 1.408
R19395 vss.n15899 vss.n15898 1.408
R19396 vss.n15979 vss.n15978 1.408
R19397 vss.n16030 vss.n16028 1.408
R19398 vss.n16115 vss.n16114 1.408
R19399 vss.n16135 vss.n16134 1.408
R19400 vss.n16215 vss.n16214 1.408
R19401 vss.n15251 vss.n15250 1.408
R19402 vss.n15375 vss.n15374 1.408
R19403 vss.n15452 vss.n15451 1.408
R19404 vss.n15611 vss.n15610 1.408
R19405 vss.n15688 vss.n15687 1.408
R19406 vss.n15839 vss.n15838 1.408
R19407 vss.n21796 vss.n21795 1.4
R19408 vss.n3745 vss.n3744 1.4
R19409 vss.n21997 vss.n21996 1.396
R19410 vss.n3946 vss.n3945 1.396
R19411 vss.n14403 vss.n14402 1.394
R19412 vss.n14634 vss.n14633 1.394
R19413 vss.n13556 vss.n13555 1.394
R19414 vss.n13292 vss.n13291 1.394
R19415 vss.n14914 vss.n14913 1.394
R19416 vss.n14942 vss.n14941 1.394
R19417 vss.n15027 vss.n15026 1.394
R19418 vss.n10472 vss.n10471 1.394
R19419 vss.n11055 vss.n11054 1.394
R19420 vss.n13995 vss.n13994 1.394
R19421 vss.n11587 vss.n11586 1.394
R19422 vss.n12577 vss.n12576 1.394
R19423 vss.n12449 vss.n12448 1.394
R19424 vss.n12611 vss.n12610 1.394
R19425 vss.n10840 vss.n10839 1.394
R19426 vss.n10884 vss.n10883 1.394
R19427 vss.n20326 vss.n17604 1.39
R19428 vss.n6936 vss.n4214 1.39
R19429 vss.n9203 vss.t1 1.368
R19430 vss.n19025 vss.n17630 1.333
R19431 vss.n19015 vss.n17632 1.333
R19432 vss.n19013 vss.n17636 1.333
R19433 vss.n19003 vss.n17640 1.333
R19434 vss.n17730 vss.n17729 1.333
R19435 vss.n17734 vss.n17731 1.333
R19436 vss.n18883 vss.n17735 1.333
R19437 vss.n18881 vss.n17741 1.333
R19438 vss.n18776 vss.n18775 1.333
R19439 vss.n18768 vss.n17835 1.333
R19440 vss.n17844 vss.n17842 1.333
R19441 vss.n17855 vss.n17845 1.333
R19442 vss.n17943 vss.n17942 1.333
R19443 vss.n17947 vss.n17944 1.333
R19444 vss.n18642 vss.n17948 1.333
R19445 vss.n18640 vss.n17954 1.333
R19446 vss.n18535 vss.n18534 1.333
R19447 vss.n18527 vss.n18048 1.333
R19448 vss.n18057 vss.n18055 1.333
R19449 vss.n18068 vss.n18058 1.333
R19450 vss.n18156 vss.n18155 1.333
R19451 vss.n18160 vss.n18157 1.333
R19452 vss.n18401 vss.n18161 1.333
R19453 vss.n18399 vss.n18167 1.333
R19454 vss.n18294 vss.n18293 1.333
R19455 vss.n18286 vss.n18261 1.333
R19456 vss.n18270 vss.n18268 1.333
R19457 vss.n18273 vss.n18271 1.333
R19458 vss.n20291 vss.n17622 1.333
R19459 vss.n20286 vss.n19034 1.333
R19460 vss.n20279 vss.n20278 1.333
R19461 vss.n19045 vss.n19042 1.333
R19462 vss.n20169 vss.n20168 1.333
R19463 vss.n20161 vss.n19135 1.333
R19464 vss.n20159 vss.n19143 1.333
R19465 vss.n20149 vss.n19147 1.333
R19466 vss.n19237 vss.n19236 1.333
R19467 vss.n19241 vss.n19238 1.333
R19468 vss.n20029 vss.n19242 1.333
R19469 vss.n20027 vss.n19248 1.333
R19470 vss.n19922 vss.n19921 1.333
R19471 vss.n19914 vss.n19342 1.333
R19472 vss.n19912 vss.n19350 1.333
R19473 vss.n19902 vss.n19354 1.333
R19474 vss.n19444 vss.n19443 1.333
R19475 vss.n19448 vss.n19445 1.333
R19476 vss.n19782 vss.n19449 1.333
R19477 vss.n19780 vss.n19455 1.333
R19478 vss.n19675 vss.n19674 1.333
R19479 vss.n19667 vss.n19549 1.333
R19480 vss.n19665 vss.n19557 1.333
R19481 vss.n19655 vss.n19561 1.333
R19482 vss.n5635 vss.n4240 1.333
R19483 vss.n5625 vss.n4242 1.333
R19484 vss.n5623 vss.n4246 1.333
R19485 vss.n5613 vss.n4250 1.333
R19486 vss.n4340 vss.n4339 1.333
R19487 vss.n4344 vss.n4341 1.333
R19488 vss.n5493 vss.n4345 1.333
R19489 vss.n5491 vss.n4351 1.333
R19490 vss.n5386 vss.n5385 1.333
R19491 vss.n5378 vss.n4445 1.333
R19492 vss.n4454 vss.n4452 1.333
R19493 vss.n4465 vss.n4455 1.333
R19494 vss.n4553 vss.n4552 1.333
R19495 vss.n4557 vss.n4554 1.333
R19496 vss.n5252 vss.n4558 1.333
R19497 vss.n5250 vss.n4564 1.333
R19498 vss.n5145 vss.n5144 1.333
R19499 vss.n5137 vss.n4658 1.333
R19500 vss.n4667 vss.n4665 1.333
R19501 vss.n4678 vss.n4668 1.333
R19502 vss.n4766 vss.n4765 1.333
R19503 vss.n4770 vss.n4767 1.333
R19504 vss.n5011 vss.n4771 1.333
R19505 vss.n5009 vss.n4777 1.333
R19506 vss.n4904 vss.n4903 1.333
R19507 vss.n4896 vss.n4871 1.333
R19508 vss.n4880 vss.n4878 1.333
R19509 vss.n4883 vss.n4881 1.333
R19510 vss.n6901 vss.n4232 1.333
R19511 vss.n6896 vss.n5644 1.333
R19512 vss.n6889 vss.n6888 1.333
R19513 vss.n5655 vss.n5652 1.333
R19514 vss.n6779 vss.n6778 1.333
R19515 vss.n6771 vss.n5745 1.333
R19516 vss.n6769 vss.n5753 1.333
R19517 vss.n6759 vss.n5757 1.333
R19518 vss.n5847 vss.n5846 1.333
R19519 vss.n5851 vss.n5848 1.333
R19520 vss.n6639 vss.n5852 1.333
R19521 vss.n6637 vss.n5858 1.333
R19522 vss.n6532 vss.n6531 1.333
R19523 vss.n6524 vss.n5952 1.333
R19524 vss.n6522 vss.n5960 1.333
R19525 vss.n6512 vss.n5964 1.333
R19526 vss.n6054 vss.n6053 1.333
R19527 vss.n6058 vss.n6055 1.333
R19528 vss.n6392 vss.n6059 1.333
R19529 vss.n6390 vss.n6065 1.333
R19530 vss.n6285 vss.n6284 1.333
R19531 vss.n6277 vss.n6159 1.333
R19532 vss.n6275 vss.n6167 1.333
R19533 vss.n6265 vss.n6171 1.333
R19534 vss.n22749 vss.n22742 1.28
R19535 vss.n22751 vss.n22749 1.28
R19536 vss.n22645 vss.n22644 1.28
R19537 vss.n22644 vss.n22637 1.28
R19538 vss.n22541 vss.n22534 1.28
R19539 vss.n22543 vss.n22541 1.28
R19540 vss.n22437 vss.n22436 1.28
R19541 vss.n22436 vss.n22429 1.28
R19542 vss.n22333 vss.n22326 1.28
R19543 vss.n22335 vss.n22333 1.28
R19544 vss.n22229 vss.n22228 1.28
R19545 vss.n22228 vss.n22221 1.28
R19546 vss.n22125 vss.n22118 1.28
R19547 vss.n22127 vss.n22125 1.28
R19548 vss.n21573 vss.n21572 1.28
R19549 vss.n21572 vss.n21565 1.28
R19550 vss.n21469 vss.n21462 1.28
R19551 vss.n21471 vss.n21469 1.28
R19552 vss.n21365 vss.n21364 1.28
R19553 vss.n21364 vss.n21357 1.28
R19554 vss.n21261 vss.n21254 1.28
R19555 vss.n21263 vss.n21261 1.28
R19556 vss.n21157 vss.n21156 1.28
R19557 vss.n21156 vss.n21149 1.28
R19558 vss.n21053 vss.n21046 1.28
R19559 vss.n21055 vss.n21053 1.28
R19560 vss.n20949 vss.n20948 1.28
R19561 vss.n20948 vss.n20941 1.28
R19562 vss.n8912 vss.n8905 1.28
R19563 vss.n8914 vss.n8912 1.28
R19564 vss.n8808 vss.n8807 1.28
R19565 vss.n8807 vss.n8800 1.28
R19566 vss.n8704 vss.n8697 1.28
R19567 vss.n8706 vss.n8704 1.28
R19568 vss.n8600 vss.n8599 1.28
R19569 vss.n8599 vss.n8592 1.28
R19570 vss.n8496 vss.n8489 1.28
R19571 vss.n8498 vss.n8496 1.28
R19572 vss.n8392 vss.n8391 1.28
R19573 vss.n8391 vss.n8384 1.28
R19574 vss.n8288 vss.n8281 1.28
R19575 vss.n8290 vss.n8288 1.28
R19576 vss.n8184 vss.n8183 1.28
R19577 vss.n8183 vss.n8176 1.28
R19578 vss.n8080 vss.n8073 1.28
R19579 vss.n8082 vss.n8080 1.28
R19580 vss.n7976 vss.n7975 1.28
R19581 vss.n7975 vss.n7968 1.28
R19582 vss.n7872 vss.n7865 1.28
R19583 vss.n7874 vss.n7872 1.28
R19584 vss.n7767 vss.n7766 1.28
R19585 vss.n7766 vss.n7759 1.28
R19586 vss.n7663 vss.n7656 1.28
R19587 vss.n7665 vss.n7663 1.28
R19588 vss.n7559 vss.n7558 1.28
R19589 vss.n7558 vss.n7551 1.28
R19590 vss.n16434 vss.n16427 1.28
R19591 vss.n16537 vss.n16530 1.28
R19592 vss.n16724 vss.n16723 1.28
R19593 vss.n16739 vss.n16730 1.28
R19594 vss.n16834 vss.n16827 1.28
R19595 vss.n16853 vss.n16852 1.28
R19596 vss.n16954 vss.n16953 1.28
R19597 vss.n16969 vss.n16960 1.28
R19598 vss.n17070 vss.n17069 1.28
R19599 vss.n17089 vss.n17088 1.28
R19600 vss.n17190 vss.n17189 1.28
R19601 vss.n17205 vss.n17196 1.28
R19602 vss.n17326 vss.n17325 1.28
R19603 vss.n15907 vss.n15897 1.28
R19604 vss.n16002 vss.n16001 1.28
R19605 vss.n16014 vss.n16007 1.28
R19606 vss.n16114 vss.n16107 1.28
R19607 vss.n16143 vss.n16133 1.28
R19608 vss.n16238 vss.n16237 1.28
R19609 vss.n15286 vss.n15279 1.28
R19610 vss.n15353 vss.n15346 1.28
R19611 vss.n15487 vss.n15480 1.28
R19612 vss.n15590 vss.n15583 1.28
R19613 vss.n15723 vss.n15716 1.28
R19614 vss.n15814 vss.n15807 1.28
R19615 vss.n9117 vss.n9115 1.266
R19616 vss.n18964 vss.n18963 1.244
R19617 vss.n18963 vss.n17676 1.244
R19618 vss.n18939 vss.n17691 1.244
R19619 vss.n17698 vss.n17691 1.244
R19620 vss.n18836 vss.n17777 1.244
R19621 vss.n18836 vss.n18835 1.244
R19622 vss.n18821 vss.n18820 1.244
R19623 vss.n18820 vss.n17797 1.244
R19624 vss.n18718 vss.n17884 1.244
R19625 vss.n18718 vss.n17885 1.244
R19626 vss.n18698 vss.n17904 1.244
R19627 vss.n17911 vss.n17904 1.244
R19628 vss.n18595 vss.n17990 1.244
R19629 vss.n18595 vss.n18594 1.244
R19630 vss.n18580 vss.n18579 1.244
R19631 vss.n18579 vss.n18010 1.244
R19632 vss.n18477 vss.n18097 1.244
R19633 vss.n18477 vss.n18098 1.244
R19634 vss.n18457 vss.n18117 1.244
R19635 vss.n18124 vss.n18117 1.244
R19636 vss.n18354 vss.n18203 1.244
R19637 vss.n18354 vss.n18353 1.244
R19638 vss.n18339 vss.n18338 1.244
R19639 vss.n18338 vss.n18223 1.244
R19640 vss.n20368 vss.n20367 1.244
R19641 vss.n20229 vss.n19077 1.244
R19642 vss.n20229 vss.n20228 1.244
R19643 vss.n20214 vss.n20213 1.244
R19644 vss.n20213 vss.n19097 1.244
R19645 vss.n20110 vss.n20109 1.244
R19646 vss.n20109 vss.n19183 1.244
R19647 vss.n20085 vss.n19198 1.244
R19648 vss.n19205 vss.n19198 1.244
R19649 vss.n19982 vss.n19284 1.244
R19650 vss.n19982 vss.n19981 1.244
R19651 vss.n19967 vss.n19966 1.244
R19652 vss.n19966 vss.n19304 1.244
R19653 vss.n19863 vss.n19862 1.244
R19654 vss.n19862 vss.n19390 1.244
R19655 vss.n19838 vss.n19405 1.244
R19656 vss.n19412 vss.n19405 1.244
R19657 vss.n19735 vss.n19491 1.244
R19658 vss.n19735 vss.n19734 1.244
R19659 vss.n19720 vss.n19719 1.244
R19660 vss.n19719 vss.n19511 1.244
R19661 vss.n19620 vss.n19619 1.244
R19662 vss.n5574 vss.n5573 1.244
R19663 vss.n5573 vss.n4286 1.244
R19664 vss.n5549 vss.n4301 1.244
R19665 vss.n4308 vss.n4301 1.244
R19666 vss.n5446 vss.n4387 1.244
R19667 vss.n5446 vss.n5445 1.244
R19668 vss.n5431 vss.n5430 1.244
R19669 vss.n5430 vss.n4407 1.244
R19670 vss.n5328 vss.n4494 1.244
R19671 vss.n5328 vss.n4495 1.244
R19672 vss.n5308 vss.n4514 1.244
R19673 vss.n4521 vss.n4514 1.244
R19674 vss.n5205 vss.n4600 1.244
R19675 vss.n5205 vss.n5204 1.244
R19676 vss.n5190 vss.n5189 1.244
R19677 vss.n5189 vss.n4620 1.244
R19678 vss.n5087 vss.n4707 1.244
R19679 vss.n5087 vss.n4708 1.244
R19680 vss.n5067 vss.n4727 1.244
R19681 vss.n4734 vss.n4727 1.244
R19682 vss.n4964 vss.n4813 1.244
R19683 vss.n4964 vss.n4963 1.244
R19684 vss.n4949 vss.n4948 1.244
R19685 vss.n4948 vss.n4833 1.244
R19686 vss.n6978 vss.n6977 1.244
R19687 vss.n6839 vss.n5687 1.244
R19688 vss.n6839 vss.n6838 1.244
R19689 vss.n6824 vss.n6823 1.244
R19690 vss.n6823 vss.n5707 1.244
R19691 vss.n6720 vss.n6719 1.244
R19692 vss.n6719 vss.n5793 1.244
R19693 vss.n6695 vss.n5808 1.244
R19694 vss.n5815 vss.n5808 1.244
R19695 vss.n6592 vss.n5894 1.244
R19696 vss.n6592 vss.n6591 1.244
R19697 vss.n6577 vss.n6576 1.244
R19698 vss.n6576 vss.n5914 1.244
R19699 vss.n6473 vss.n6472 1.244
R19700 vss.n6472 vss.n6000 1.244
R19701 vss.n6448 vss.n6015 1.244
R19702 vss.n6022 vss.n6015 1.244
R19703 vss.n6345 vss.n6101 1.244
R19704 vss.n6345 vss.n6344 1.244
R19705 vss.n6330 vss.n6329 1.244
R19706 vss.n6329 vss.n6121 1.244
R19707 vss.n6230 vss.n6229 1.244
R19708 vss.n10768 vss.n10767 1.234
R19709 vss.n13396 vss.n13395 1.234
R19710 vss.n17296 vss.n17295 1.195
R19711 vss.n15795 vss.n15792 1.195
R19712 vss.n15121 vss.n15120 1.195
R19713 vss.n13810 vss.n13809 1.184
R19714 vss.n20407 vss.n20406 1.184
R19715 vss.n7017 vss.n7016 1.184
R19716 vss.n10456 bandgapmd_0.vss 1.183
R19717 vss.n21619 vss.n21618 1.181
R19718 vss.n3568 vss.n3567 1.181
R19719 vss.n8972 vss.n8946 1.17
R19720 vss.n8978 vss.n8976 1.165
R19721 vss.n19027 vss.n19026 1.155
R19722 vss.n19002 vss.n19001 1.155
R19723 vss.n17648 vss.n17646 1.155
R19724 vss.n18903 vss.n17723 1.155
R19725 vss.n18898 vss.n17725 1.155
R19726 vss.n17747 vss.n17743 1.155
R19727 vss.n17755 vss.n17744 1.155
R19728 vss.n17830 vss.n17829 1.155
R19729 vss.n17834 vss.n17831 1.155
R19730 vss.n18758 vss.n17853 1.155
R19731 vss.n18753 vss.n17854 1.155
R19732 vss.n18662 vss.n17936 1.155
R19733 vss.n18657 vss.n17938 1.155
R19734 vss.n17960 vss.n17956 1.155
R19735 vss.n17968 vss.n17957 1.155
R19736 vss.n18043 vss.n18042 1.155
R19737 vss.n18047 vss.n18044 1.155
R19738 vss.n18517 vss.n18066 1.155
R19739 vss.n18512 vss.n18067 1.155
R19740 vss.n18421 vss.n18149 1.155
R19741 vss.n18416 vss.n18151 1.155
R19742 vss.n18173 vss.n18169 1.155
R19743 vss.n18181 vss.n18170 1.155
R19744 vss.n18256 vss.n18255 1.155
R19745 vss.n18260 vss.n18257 1.155
R19746 vss.n18274 vss.n17624 1.155
R19747 vss.n20369 vss.n17575 1.155
R19748 vss.n20292 vss.n17621 1.155
R19749 vss.n20272 vss.n20271 1.155
R19750 vss.n19055 vss.n19043 1.155
R19751 vss.n19130 vss.n19129 1.155
R19752 vss.n19134 vss.n19131 1.155
R19753 vss.n20148 vss.n20147 1.155
R19754 vss.n19155 vss.n19153 1.155
R19755 vss.n20049 vss.n19230 1.155
R19756 vss.n20044 vss.n19232 1.155
R19757 vss.n19254 vss.n19250 1.155
R19758 vss.n19262 vss.n19251 1.155
R19759 vss.n19337 vss.n19336 1.155
R19760 vss.n19341 vss.n19338 1.155
R19761 vss.n19901 vss.n19900 1.155
R19762 vss.n19362 vss.n19360 1.155
R19763 vss.n19802 vss.n19437 1.155
R19764 vss.n19797 vss.n19439 1.155
R19765 vss.n19461 vss.n19457 1.155
R19766 vss.n19469 vss.n19458 1.155
R19767 vss.n19544 vss.n19543 1.155
R19768 vss.n19548 vss.n19545 1.155
R19769 vss.n19654 vss.n19653 1.155
R19770 vss.n19569 vss.n19567 1.155
R19771 vss.n5637 vss.n5636 1.155
R19772 vss.n5612 vss.n5611 1.155
R19773 vss.n4258 vss.n4256 1.155
R19774 vss.n5513 vss.n4333 1.155
R19775 vss.n5508 vss.n4335 1.155
R19776 vss.n4357 vss.n4353 1.155
R19777 vss.n4365 vss.n4354 1.155
R19778 vss.n4440 vss.n4439 1.155
R19779 vss.n4444 vss.n4441 1.155
R19780 vss.n5368 vss.n4463 1.155
R19781 vss.n5363 vss.n4464 1.155
R19782 vss.n5272 vss.n4546 1.155
R19783 vss.n5267 vss.n4548 1.155
R19784 vss.n4570 vss.n4566 1.155
R19785 vss.n4578 vss.n4567 1.155
R19786 vss.n4653 vss.n4652 1.155
R19787 vss.n4657 vss.n4654 1.155
R19788 vss.n5127 vss.n4676 1.155
R19789 vss.n5122 vss.n4677 1.155
R19790 vss.n5031 vss.n4759 1.155
R19791 vss.n5026 vss.n4761 1.155
R19792 vss.n4783 vss.n4779 1.155
R19793 vss.n4791 vss.n4780 1.155
R19794 vss.n4866 vss.n4865 1.155
R19795 vss.n4870 vss.n4867 1.155
R19796 vss.n4884 vss.n4234 1.155
R19797 vss.n6979 vss.n4185 1.155
R19798 vss.n6902 vss.n4231 1.155
R19799 vss.n6882 vss.n6881 1.155
R19800 vss.n5665 vss.n5653 1.155
R19801 vss.n5740 vss.n5739 1.155
R19802 vss.n5744 vss.n5741 1.155
R19803 vss.n6758 vss.n6757 1.155
R19804 vss.n5765 vss.n5763 1.155
R19805 vss.n6659 vss.n5840 1.155
R19806 vss.n6654 vss.n5842 1.155
R19807 vss.n5864 vss.n5860 1.155
R19808 vss.n5872 vss.n5861 1.155
R19809 vss.n5947 vss.n5946 1.155
R19810 vss.n5951 vss.n5948 1.155
R19811 vss.n6511 vss.n6510 1.155
R19812 vss.n5972 vss.n5970 1.155
R19813 vss.n6412 vss.n6047 1.155
R19814 vss.n6407 vss.n6049 1.155
R19815 vss.n6071 vss.n6067 1.155
R19816 vss.n6079 vss.n6068 1.155
R19817 vss.n6154 vss.n6153 1.155
R19818 vss.n6158 vss.n6155 1.155
R19819 vss.n6264 vss.n6263 1.155
R19820 vss.n6179 vss.n6177 1.155
R19821 vss.n3489 vss.n3488 1.155
R19822 vss.n1464 vss.n1463 1.155
R19823 vss.n16308 vss.n16307 1.152
R19824 vss.n16413 vss.n16412 1.152
R19825 vss.n16544 vss.n16543 1.152
R19826 vss.n16649 vss.n16648 1.152
R19827 vss.n16716 vss.n16715 1.152
R19828 vss.n16739 vss.n16738 1.152
R19829 vss.n16848 vss.n16839 1.152
R19830 vss.n16841 vss.n16840 1.152
R19831 vss.n16946 vss.n16945 1.152
R19832 vss.n16969 vss.n16968 1.152
R19833 vss.n17084 vss.n17075 1.152
R19834 vss.n17083 vss.n17082 1.152
R19835 vss.n17182 vss.n17181 1.152
R19836 vss.n17205 vss.n17204 1.152
R19837 vss.n17277 vss.n17276 1.152
R19838 vss.n15893 vss.n15892 1.152
R19839 vss.n15885 vss.n15884 1.152
R19840 vss.n15993 vss.n15992 1.152
R19841 vss.n16016 vss.n16014 1.152
R19842 vss.n16129 vss.n16128 1.152
R19843 vss.n16121 vss.n16120 1.152
R19844 vss.n16229 vss.n16228 1.152
R19845 vss.n15265 vss.n15264 1.152
R19846 vss.n15361 vss.n15360 1.152
R19847 vss.n15466 vss.n15465 1.152
R19848 vss.n15597 vss.n15596 1.152
R19849 vss.n15702 vss.n15701 1.152
R19850 vss.n15825 vss.n15824 1.152
R19851 vss.n9091 vss.n9090 1.148
R19852 vss.n21669 vss.n21640 1.146
R19853 vss.n3618 vss.n3589 1.146
R19854 vss.n19623 vss.n19622 1.142
R19855 vss.n6233 vss.n6232 1.142
R19856 vss.n10251 vss.n10228 1.137
R19857 vss.n22742 vss.n22741 1.137
R19858 vss.n22751 vss.n22750 1.137
R19859 vss.n22645 vss.n22635 1.137
R19860 vss.n22637 vss.n22636 1.137
R19861 vss.n22534 vss.n22533 1.137
R19862 vss.n22543 vss.n22542 1.137
R19863 vss.n22437 vss.n22427 1.137
R19864 vss.n22429 vss.n22428 1.137
R19865 vss.n22326 vss.n22325 1.137
R19866 vss.n22335 vss.n22334 1.137
R19867 vss.n22229 vss.n22219 1.137
R19868 vss.n22221 vss.n22220 1.137
R19869 vss.n22118 vss.n22117 1.137
R19870 vss.n22127 vss.n22126 1.137
R19871 vss.n21573 vss.n21563 1.137
R19872 vss.n21565 vss.n21564 1.137
R19873 vss.n21462 vss.n21461 1.137
R19874 vss.n21471 vss.n21470 1.137
R19875 vss.n21365 vss.n21355 1.137
R19876 vss.n21357 vss.n21356 1.137
R19877 vss.n21254 vss.n21253 1.137
R19878 vss.n21263 vss.n21262 1.137
R19879 vss.n21157 vss.n21147 1.137
R19880 vss.n21149 vss.n21148 1.137
R19881 vss.n21046 vss.n21045 1.137
R19882 vss.n21055 vss.n21054 1.137
R19883 vss.n20949 vss.n20939 1.137
R19884 vss.n20941 vss.n20940 1.137
R19885 vss.n8905 vss.n8904 1.137
R19886 vss.n8914 vss.n8913 1.137
R19887 vss.n8808 vss.n8798 1.137
R19888 vss.n8800 vss.n8799 1.137
R19889 vss.n8697 vss.n8696 1.137
R19890 vss.n8706 vss.n8705 1.137
R19891 vss.n8600 vss.n8590 1.137
R19892 vss.n8592 vss.n8591 1.137
R19893 vss.n8489 vss.n8488 1.137
R19894 vss.n8498 vss.n8497 1.137
R19895 vss.n8392 vss.n8382 1.137
R19896 vss.n8384 vss.n8383 1.137
R19897 vss.n8281 vss.n8280 1.137
R19898 vss.n8290 vss.n8289 1.137
R19899 vss.n8184 vss.n8174 1.137
R19900 vss.n8176 vss.n8175 1.137
R19901 vss.n8073 vss.n8072 1.137
R19902 vss.n8082 vss.n8081 1.137
R19903 vss.n7976 vss.n7966 1.137
R19904 vss.n7968 vss.n7967 1.137
R19905 vss.n7865 vss.n7864 1.137
R19906 vss.n7874 vss.n7873 1.137
R19907 vss.n7767 vss.n7757 1.137
R19908 vss.n7759 vss.n7758 1.137
R19909 vss.n7656 vss.n7655 1.137
R19910 vss.n7665 vss.n7664 1.137
R19911 vss.n7559 vss.n7549 1.137
R19912 vss.n7551 vss.n7550 1.137
R19913 vss.n17306 vss.n17305 1.131
R19914 vss.n15805 vss.n15804 1.131
R19915 vss.n13772 vss.n13771 1.13
R19916 vss.n12099 vss.n12098 1.13
R19917 vss.n13522 vss.n13521 1.13
R19918 vss.n20650 vss.n20642 1.129
R19919 vss.n20668 vss.n20660 1.129
R19920 vss.n21853 vss.n21848 1.129
R19921 vss.n21742 vss.n21741 1.129
R19922 vss.n10393 vss.n10391 1.129
R19923 vss.n12072 vss.n12065 1.129
R19924 vss.n10801 vss.n10794 1.129
R19925 vss.n10964 vss.n10957 1.129
R19926 vss.n11004 vss.n10997 1.129
R19927 vss.n13854 vss.n13847 1.129
R19928 vss.n14075 vss.n14068 1.129
R19929 vss.n11721 vss.n11714 1.129
R19930 vss.n11065 vss.n11058 1.129
R19931 vss.n13352 vss.n13345 1.129
R19932 vss.n14697 vss.n14690 1.129
R19933 vss.n14190 vss.n14183 1.129
R19934 vss.n14232 vss.n14225 1.129
R19935 vss.n12873 vss.n12872 1.129
R19936 vss.n12872 vss.n12865 1.129
R19937 vss.n12921 vss.n12908 1.129
R19938 vss.n12922 vss.n12921 1.129
R19939 vss.n12467 vss.n12460 1.129
R19940 vss.n12508 vss.n12495 1.129
R19941 vss.n12509 vss.n12508 1.129
R19942 vss.n3802 vss.n3797 1.129
R19943 vss.n3691 vss.n3690 1.129
R19944 vss.n7260 vss.n7252 1.129
R19945 vss.n7278 vss.n7270 1.129
R19946 vss.n1871 vss.n1863 1.129
R19947 vss.n1890 vss.n1881 1.129
R19948 vss.n2116 vss.n2107 1.129
R19949 vss.n2134 vss.n2125 1.129
R19950 vss.n2360 vss.n2351 1.129
R19951 vss.n2378 vss.n2369 1.129
R19952 vss.n2604 vss.n2595 1.129
R19953 vss.n2623 vss.n2614 1.129
R19954 vss.n2842 vss.n1546 1.129
R19955 vss.n2843 vss.n2842 1.129
R19956 vss.n2861 vss.n2852 1.129
R19957 vss.n3087 vss.n3078 1.129
R19958 vss.n3105 vss.n3096 1.129
R19959 vss.n3331 vss.n3322 1.129
R19960 vss.n3349 vss.n3341 1.129
R19961 vss.n332 vss.n324 1.129
R19962 vss.n351 vss.n342 1.129
R19963 vss.n577 vss.n568 1.129
R19964 vss.n595 vss.n586 1.129
R19965 vss.n821 vss.n812 1.129
R19966 vss.n839 vss.n830 1.129
R19967 vss.n1065 vss.n1056 1.129
R19968 vss.n1084 vss.n1075 1.129
R19969 vss.n1310 vss.n1301 1.129
R19970 vss.n23404 vss.n23395 1.129
R19971 vss.n23179 vss.n23170 1.129
R19972 vss.n23161 vss.n23152 1.129
R19973 vss.n22935 vss.n22926 1.129
R19974 vss.n22916 vss.n22908 1.129
R19975 vss.n19616 vss.n19615 1.125
R19976 vss.n6226 vss.n6225 1.125
R19977 vss.n15214 vss.n15213 1.117
R19978 vss.n14286 vss.n14285 1.08
R19979 vss.n13603 vss.n13602 1.08
R19980 vss.n12285 vss.n12284 1.08
R19981 vss.n12785 vss.n12784 1.08
R19982 vss.n13208 vss.n13207 1.08
R19983 vss.n13061 vss.n13060 1.08
R19984 vss.n21673 vss.n21661 1.069
R19985 vss.n3622 vss.n3610 1.069
R19986 vss.n15120 vss.n15119 1.069
R19987 vss.n18970 vss.n17668 1.066
R19988 vss.n18970 vss.n17669 1.066
R19989 vss.n18934 vss.n18933 1.066
R19990 vss.n18933 vss.n17694 1.066
R19991 vss.n18848 vss.n18847 1.066
R19992 vss.n18847 vss.n17773 1.066
R19993 vss.n18809 vss.n17804 1.066
R19994 vss.n18809 vss.n18808 1.066
R19995 vss.n18723 vss.n17877 1.066
R19996 vss.n18723 vss.n18722 1.066
R19997 vss.n18693 vss.n18692 1.066
R19998 vss.n18692 vss.n17907 1.066
R19999 vss.n18607 vss.n18606 1.066
R20000 vss.n18606 vss.n17986 1.066
R20001 vss.n18568 vss.n18017 1.066
R20002 vss.n18568 vss.n18567 1.066
R20003 vss.n18482 vss.n18090 1.066
R20004 vss.n18482 vss.n18481 1.066
R20005 vss.n18452 vss.n18451 1.066
R20006 vss.n18451 vss.n18120 1.066
R20007 vss.n18366 vss.n18365 1.066
R20008 vss.n18365 vss.n18199 1.066
R20009 vss.n18327 vss.n18230 1.066
R20010 vss.n18327 vss.n18326 1.066
R20011 vss.n17591 vss.n17590 1.066
R20012 vss.n20241 vss.n20240 1.066
R20013 vss.n20240 vss.n19073 1.066
R20014 vss.n20202 vss.n19104 1.066
R20015 vss.n20202 vss.n20201 1.066
R20016 vss.n20116 vss.n19175 1.066
R20017 vss.n20116 vss.n19176 1.066
R20018 vss.n20080 vss.n20079 1.066
R20019 vss.n20079 vss.n19201 1.066
R20020 vss.n19994 vss.n19993 1.066
R20021 vss.n19993 vss.n19280 1.066
R20022 vss.n19955 vss.n19311 1.066
R20023 vss.n19955 vss.n19954 1.066
R20024 vss.n19869 vss.n19382 1.066
R20025 vss.n19869 vss.n19383 1.066
R20026 vss.n19833 vss.n19832 1.066
R20027 vss.n19832 vss.n19408 1.066
R20028 vss.n19747 vss.n19746 1.066
R20029 vss.n19746 vss.n19487 1.066
R20030 vss.n19708 vss.n19518 1.066
R20031 vss.n19708 vss.n19707 1.066
R20032 vss.n19598 vss.n19590 1.066
R20033 vss.n5580 vss.n4278 1.066
R20034 vss.n5580 vss.n4279 1.066
R20035 vss.n5544 vss.n5543 1.066
R20036 vss.n5543 vss.n4304 1.066
R20037 vss.n5458 vss.n5457 1.066
R20038 vss.n5457 vss.n4383 1.066
R20039 vss.n5419 vss.n4414 1.066
R20040 vss.n5419 vss.n5418 1.066
R20041 vss.n5333 vss.n4487 1.066
R20042 vss.n5333 vss.n5332 1.066
R20043 vss.n5303 vss.n5302 1.066
R20044 vss.n5302 vss.n4517 1.066
R20045 vss.n5217 vss.n5216 1.066
R20046 vss.n5216 vss.n4596 1.066
R20047 vss.n5178 vss.n4627 1.066
R20048 vss.n5178 vss.n5177 1.066
R20049 vss.n5092 vss.n4700 1.066
R20050 vss.n5092 vss.n5091 1.066
R20051 vss.n5062 vss.n5061 1.066
R20052 vss.n5061 vss.n4730 1.066
R20053 vss.n4976 vss.n4975 1.066
R20054 vss.n4975 vss.n4809 1.066
R20055 vss.n4937 vss.n4840 1.066
R20056 vss.n4937 vss.n4936 1.066
R20057 vss.n4201 vss.n4200 1.066
R20058 vss.n6851 vss.n6850 1.066
R20059 vss.n6850 vss.n5683 1.066
R20060 vss.n6812 vss.n5714 1.066
R20061 vss.n6812 vss.n6811 1.066
R20062 vss.n6726 vss.n5785 1.066
R20063 vss.n6726 vss.n5786 1.066
R20064 vss.n6690 vss.n6689 1.066
R20065 vss.n6689 vss.n5811 1.066
R20066 vss.n6604 vss.n6603 1.066
R20067 vss.n6603 vss.n5890 1.066
R20068 vss.n6565 vss.n5921 1.066
R20069 vss.n6565 vss.n6564 1.066
R20070 vss.n6479 vss.n5992 1.066
R20071 vss.n6479 vss.n5993 1.066
R20072 vss.n6443 vss.n6442 1.066
R20073 vss.n6442 vss.n6018 1.066
R20074 vss.n6357 vss.n6356 1.066
R20075 vss.n6356 vss.n6097 1.066
R20076 vss.n6318 vss.n6128 1.066
R20077 vss.n6318 vss.n6317 1.066
R20078 vss.n6208 vss.n6200 1.066
R20079 vss.n15815 vss.n15814 1.064
R20080 vss.n15123 vss.n15122 1.038
R20081 vss.n10866 vss.n10865 1.035
R20082 vss.n16315 vss.n16308 1.024
R20083 vss.n16420 vss.n16413 1.024
R20084 vss.n16551 vss.n16544 1.024
R20085 vss.n16656 vss.n16649 1.024
R20086 vss.n16725 vss.n16716 1.024
R20087 vss.n16738 vss.n16737 1.024
R20088 vss.n16839 vss.n16838 1.024
R20089 vss.n16848 vss.n16841 1.024
R20090 vss.n16955 vss.n16946 1.024
R20091 vss.n16968 vss.n16967 1.024
R20092 vss.n17075 vss.n17074 1.024
R20093 vss.n17084 vss.n17083 1.024
R20094 vss.n17191 vss.n17182 1.024
R20095 vss.n17204 vss.n17203 1.024
R20096 vss.n17284 vss.n17277 1.024
R20097 vss.n15893 vss.n15883 1.024
R20098 vss.n15892 vss.n15885 1.024
R20099 vss.n16000 vss.n15993 1.024
R20100 vss.n16016 vss.n16015 1.024
R20101 vss.n16129 vss.n16119 1.024
R20102 vss.n16128 vss.n16121 1.024
R20103 vss.n16236 vss.n16229 1.024
R20104 vss.n15272 vss.n15265 1.024
R20105 vss.n15368 vss.n15361 1.024
R20106 vss.n15473 vss.n15466 1.024
R20107 vss.n15604 vss.n15597 1.024
R20108 vss.n15709 vss.n15702 1.024
R20109 vss.n15832 vss.n15825 1.024
R20110 vss.t172 vss.n12441 1.015
R20111 vss.n13450 vss.n13440 1.013
R20112 vss.n13027 vss.n13026 1.013
R20113 vss.n10582 vss.n10572 1.013
R20114 vss.n10741 vss.n10740 1.013
R20115 vss.n13637 vss.n13627 1.013
R20116 vss.n13691 vss.n13690 1.013
R20117 vss.n11386 vss.n11376 1.013
R20118 vss.n11374 vss.n11373 1.013
R20119 vss.n22631 vss.n22630 0.995
R20120 vss.n22630 vss.n22623 0.995
R20121 vss.n22555 vss.n22548 0.995
R20122 vss.n22557 vss.n22555 0.995
R20123 vss.n22423 vss.n22422 0.995
R20124 vss.n22422 vss.n22415 0.995
R20125 vss.n22347 vss.n22340 0.995
R20126 vss.n22349 vss.n22347 0.995
R20127 vss.n22215 vss.n22214 0.995
R20128 vss.n22214 vss.n22207 0.995
R20129 vss.n22139 vss.n22132 0.995
R20130 vss.n22141 vss.n22139 0.995
R20131 vss.n21559 vss.n21558 0.995
R20132 vss.n21558 vss.n21551 0.995
R20133 vss.n21483 vss.n21476 0.995
R20134 vss.n21485 vss.n21483 0.995
R20135 vss.n21351 vss.n21350 0.995
R20136 vss.n21350 vss.n21343 0.995
R20137 vss.n21275 vss.n21268 0.995
R20138 vss.n21277 vss.n21275 0.995
R20139 vss.n21143 vss.n21142 0.995
R20140 vss.n21142 vss.n21135 0.995
R20141 vss.n21067 vss.n21060 0.995
R20142 vss.n21069 vss.n21067 0.995
R20143 vss.n20935 vss.n20934 0.995
R20144 vss.n20934 vss.n20927 0.995
R20145 vss.n8794 vss.n8793 0.995
R20146 vss.n8793 vss.n8786 0.995
R20147 vss.n8718 vss.n8711 0.995
R20148 vss.n8720 vss.n8718 0.995
R20149 vss.n8586 vss.n8585 0.995
R20150 vss.n8585 vss.n8578 0.995
R20151 vss.n8510 vss.n8503 0.995
R20152 vss.n8512 vss.n8510 0.995
R20153 vss.n8378 vss.n8377 0.995
R20154 vss.n8377 vss.n8370 0.995
R20155 vss.n8302 vss.n8295 0.995
R20156 vss.n8304 vss.n8302 0.995
R20157 vss.n8170 vss.n8169 0.995
R20158 vss.n8169 vss.n8162 0.995
R20159 vss.n8094 vss.n8087 0.995
R20160 vss.n8096 vss.n8094 0.995
R20161 vss.n7962 vss.n7961 0.995
R20162 vss.n7961 vss.n7954 0.995
R20163 vss.n7886 vss.n7879 0.995
R20164 vss.n7888 vss.n7886 0.995
R20165 vss.n7753 vss.n7752 0.995
R20166 vss.n7752 vss.n7745 0.995
R20167 vss.n7677 vss.n7670 0.995
R20168 vss.n7679 vss.n7677 0.995
R20169 vss.n7545 vss.n7544 0.995
R20170 vss.n7544 vss.n7537 0.995
R20171 vss.n17285 vss.n17284 0.993
R20172 vss.n20352 vss.n20351 0.984
R20173 vss.n20351 vss.n20350 0.984
R20174 vss.n6962 vss.n6961 0.984
R20175 vss.n6961 vss.n6960 0.984
R20176 vss.n18995 vss.n18994 0.977
R20177 vss.n17658 vss.n17647 0.977
R20178 vss.n18912 vss.n18911 0.977
R20179 vss.n18904 vss.n17716 0.977
R20180 vss.n18871 vss.n17753 0.977
R20181 vss.n18866 vss.n17754 0.977
R20182 vss.n18790 vss.n17823 0.977
R20183 vss.n18785 vss.n17825 0.977
R20184 vss.n18752 vss.n17858 0.977
R20185 vss.n18745 vss.n17862 0.977
R20186 vss.n18671 vss.n18670 0.977
R20187 vss.n18663 vss.n17929 0.977
R20188 vss.n18630 vss.n17966 0.977
R20189 vss.n18625 vss.n17967 0.977
R20190 vss.n18549 vss.n18036 0.977
R20191 vss.n18544 vss.n18038 0.977
R20192 vss.n18511 vss.n18071 0.977
R20193 vss.n18504 vss.n18075 0.977
R20194 vss.n18430 vss.n18429 0.977
R20195 vss.n18422 vss.n18142 0.977
R20196 vss.n18389 vss.n18179 0.977
R20197 vss.n18384 vss.n18180 0.977
R20198 vss.n18308 vss.n18249 0.977
R20199 vss.n18303 vss.n18251 0.977
R20200 vss.n20264 vss.n19052 0.977
R20201 vss.n20259 vss.n19053 0.977
R20202 vss.n20183 vss.n19123 0.977
R20203 vss.n20178 vss.n19125 0.977
R20204 vss.n20141 vss.n20140 0.977
R20205 vss.n19165 vss.n19154 0.977
R20206 vss.n20058 vss.n20057 0.977
R20207 vss.n20050 vss.n19223 0.977
R20208 vss.n20017 vss.n19260 0.977
R20209 vss.n20012 vss.n19261 0.977
R20210 vss.n19936 vss.n19330 0.977
R20211 vss.n19931 vss.n19332 0.977
R20212 vss.n19894 vss.n19893 0.977
R20213 vss.n19372 vss.n19361 0.977
R20214 vss.n19811 vss.n19810 0.977
R20215 vss.n19803 vss.n19430 0.977
R20216 vss.n19770 vss.n19467 0.977
R20217 vss.n19765 vss.n19468 0.977
R20218 vss.n19689 vss.n19537 0.977
R20219 vss.n19684 vss.n19539 0.977
R20220 vss.n19647 vss.n19646 0.977
R20221 vss.n19579 vss.n19568 0.977
R20222 vss.n5605 vss.n5604 0.977
R20223 vss.n4268 vss.n4257 0.977
R20224 vss.n5522 vss.n5521 0.977
R20225 vss.n5514 vss.n4326 0.977
R20226 vss.n5481 vss.n4363 0.977
R20227 vss.n5476 vss.n4364 0.977
R20228 vss.n5400 vss.n4433 0.977
R20229 vss.n5395 vss.n4435 0.977
R20230 vss.n5362 vss.n4468 0.977
R20231 vss.n5355 vss.n4472 0.977
R20232 vss.n5281 vss.n5280 0.977
R20233 vss.n5273 vss.n4539 0.977
R20234 vss.n5240 vss.n4576 0.977
R20235 vss.n5235 vss.n4577 0.977
R20236 vss.n5159 vss.n4646 0.977
R20237 vss.n5154 vss.n4648 0.977
R20238 vss.n5121 vss.n4681 0.977
R20239 vss.n5114 vss.n4685 0.977
R20240 vss.n5040 vss.n5039 0.977
R20241 vss.n5032 vss.n4752 0.977
R20242 vss.n4999 vss.n4789 0.977
R20243 vss.n4994 vss.n4790 0.977
R20244 vss.n4918 vss.n4859 0.977
R20245 vss.n4913 vss.n4861 0.977
R20246 vss.n6874 vss.n5662 0.977
R20247 vss.n6869 vss.n5663 0.977
R20248 vss.n6793 vss.n5733 0.977
R20249 vss.n6788 vss.n5735 0.977
R20250 vss.n6751 vss.n6750 0.977
R20251 vss.n5775 vss.n5764 0.977
R20252 vss.n6668 vss.n6667 0.977
R20253 vss.n6660 vss.n5833 0.977
R20254 vss.n6627 vss.n5870 0.977
R20255 vss.n6622 vss.n5871 0.977
R20256 vss.n6546 vss.n5940 0.977
R20257 vss.n6541 vss.n5942 0.977
R20258 vss.n6504 vss.n6503 0.977
R20259 vss.n5982 vss.n5971 0.977
R20260 vss.n6421 vss.n6420 0.977
R20261 vss.n6413 vss.n6040 0.977
R20262 vss.n6380 vss.n6077 0.977
R20263 vss.n6375 vss.n6078 0.977
R20264 vss.n6299 vss.n6147 0.977
R20265 vss.n6294 vss.n6149 0.977
R20266 vss.n6257 vss.n6256 0.977
R20267 vss.n6189 vss.n6178 0.977
R20268 vss.n13948 vss.n13947 0.975
R20269 vss.n11688 vss.n11685 0.975
R20270 vss.n11938 vss.n11935 0.975
R20271 vss.n12262 vss.n12259 0.975
R20272 vss.n9152 vss.n9151 0.969
R20273 vss.n9063 vss.n9062 0.969
R20274 vss.n9032 vss.n9031 0.969
R20275 vss.n9125 vss.n9124 0.968
R20276 vss.n9094 vss.n9093 0.964
R20277 vss.n9002 vss.n9001 0.961
R20278 vss.n11232 vss.t174 0.95
R20279 vss.n12956 vss.t198 0.95
R20280 vss.n14997 vss.n14996 0.95
R20281 vss.n11808 vss.n11807 0.95
R20282 vss.n12395 vss.n12394 0.95
R20283 vss.n14705 vss.n14704 0.95
R20284 vss.n13442 vss.n13441 0.95
R20285 vss.n13017 vss.n13016 0.95
R20286 vss.n10574 vss.n10573 0.95
R20287 vss.n10731 vss.n10730 0.95
R20288 vss.n12027 vss.n12026 0.95
R20289 vss.n14569 vss.n14568 0.95
R20290 vss.n13629 vss.n13628 0.95
R20291 vss.n13681 vss.n13680 0.95
R20292 vss.n11378 vss.n11377 0.95
R20293 vss.n11364 vss.n11363 0.95
R20294 vss.n11307 vss.n11306 0.95
R20295 vss.n13955 vss.n13954 0.95
R20296 vss.n14175 vss.t170 0.932
R20297 vss.n17316 vss.n17315 0.919
R20298 vss.n17578 vss.n17575 0.912
R20299 vss.n4188 vss.n4185 0.912
R20300 vss.n10344 vss.n10343 0.91
R20301 vss.n10455 vss.n9154 0.909
R20302 vss.n16427 vss.n16426 0.896
R20303 vss.n16530 vss.n16529 0.896
R20304 vss.n16725 vss.n16724 0.896
R20305 vss.n16730 vss.n16729 0.896
R20306 vss.n16827 vss.n16826 0.896
R20307 vss.n16862 vss.n16853 0.896
R20308 vss.n16955 vss.n16954 0.896
R20309 vss.n16960 vss.n16959 0.896
R20310 vss.n17069 vss.n17068 0.896
R20311 vss.n17098 vss.n17089 0.896
R20312 vss.n17191 vss.n17190 0.896
R20313 vss.n17196 vss.n17195 0.896
R20314 vss.n17325 vss.n17324 0.896
R20315 vss.n15907 vss.n15906 0.896
R20316 vss.n16002 vss.n16000 0.896
R20317 vss.n16007 vss.n16006 0.896
R20318 vss.n16107 vss.n16106 0.896
R20319 vss.n16143 vss.n16142 0.896
R20320 vss.n16238 vss.n16236 0.896
R20321 vss.n15279 vss.n15278 0.896
R20322 vss.n15346 vss.n15345 0.896
R20323 vss.n15480 vss.n15479 0.896
R20324 vss.n15583 vss.n15582 0.896
R20325 vss.n15716 vss.n15715 0.896
R20326 vss.n15807 vss.n15806 0.896
R20327 vss.n12961 vss.n12960 0.89
R20328 vss.n12930 vss.n12929 0.89
R20329 vss.n18975 vss.n17661 0.888
R20330 vss.n18975 vss.n18974 0.888
R20331 vss.n18922 vss.n17704 0.888
R20332 vss.n18922 vss.n18921 0.888
R20333 vss.n18854 vss.n17765 0.888
R20334 vss.n18854 vss.n17766 0.888
R20335 vss.n18802 vss.n17811 0.888
R20336 vss.n18802 vss.n17812 0.888
R20337 vss.n18735 vss.n18734 0.888
R20338 vss.n18734 vss.n17873 0.888
R20339 vss.n18681 vss.n17917 0.888
R20340 vss.n18681 vss.n18680 0.888
R20341 vss.n18613 vss.n17978 0.888
R20342 vss.n18613 vss.n17979 0.888
R20343 vss.n18561 vss.n18024 0.888
R20344 vss.n18561 vss.n18025 0.888
R20345 vss.n18494 vss.n18493 0.888
R20346 vss.n18493 vss.n18086 0.888
R20347 vss.n18440 vss.n18130 0.888
R20348 vss.n18440 vss.n18439 0.888
R20349 vss.n18372 vss.n18191 0.888
R20350 vss.n18372 vss.n18192 0.888
R20351 vss.n18320 vss.n18237 0.888
R20352 vss.n18320 vss.n18238 0.888
R20353 vss.n20247 vss.n19065 0.888
R20354 vss.n20247 vss.n19066 0.888
R20355 vss.n20195 vss.n19111 0.888
R20356 vss.n20195 vss.n19112 0.888
R20357 vss.n20121 vss.n19168 0.888
R20358 vss.n20121 vss.n20120 0.888
R20359 vss.n20068 vss.n19211 0.888
R20360 vss.n20068 vss.n20067 0.888
R20361 vss.n20000 vss.n19272 0.888
R20362 vss.n20000 vss.n19273 0.888
R20363 vss.n19948 vss.n19318 0.888
R20364 vss.n19948 vss.n19319 0.888
R20365 vss.n19874 vss.n19375 0.888
R20366 vss.n19874 vss.n19873 0.888
R20367 vss.n19821 vss.n19418 0.888
R20368 vss.n19821 vss.n19820 0.888
R20369 vss.n19753 vss.n19479 0.888
R20370 vss.n19753 vss.n19480 0.888
R20371 vss.n19701 vss.n19525 0.888
R20372 vss.n19701 vss.n19526 0.888
R20373 vss.n19627 vss.n19582 0.888
R20374 vss.n19627 vss.n19626 0.888
R20375 vss.n5585 vss.n4271 0.888
R20376 vss.n5585 vss.n5584 0.888
R20377 vss.n5532 vss.n4314 0.888
R20378 vss.n5532 vss.n5531 0.888
R20379 vss.n5464 vss.n4375 0.888
R20380 vss.n5464 vss.n4376 0.888
R20381 vss.n5412 vss.n4421 0.888
R20382 vss.n5412 vss.n4422 0.888
R20383 vss.n5345 vss.n5344 0.888
R20384 vss.n5344 vss.n4483 0.888
R20385 vss.n5291 vss.n4527 0.888
R20386 vss.n5291 vss.n5290 0.888
R20387 vss.n5223 vss.n4588 0.888
R20388 vss.n5223 vss.n4589 0.888
R20389 vss.n5171 vss.n4634 0.888
R20390 vss.n5171 vss.n4635 0.888
R20391 vss.n5104 vss.n5103 0.888
R20392 vss.n5103 vss.n4696 0.888
R20393 vss.n5050 vss.n4740 0.888
R20394 vss.n5050 vss.n5049 0.888
R20395 vss.n4982 vss.n4801 0.888
R20396 vss.n4982 vss.n4802 0.888
R20397 vss.n4930 vss.n4847 0.888
R20398 vss.n4930 vss.n4848 0.888
R20399 vss.n6857 vss.n5675 0.888
R20400 vss.n6857 vss.n5676 0.888
R20401 vss.n6805 vss.n5721 0.888
R20402 vss.n6805 vss.n5722 0.888
R20403 vss.n6731 vss.n5778 0.888
R20404 vss.n6731 vss.n6730 0.888
R20405 vss.n6678 vss.n5821 0.888
R20406 vss.n6678 vss.n6677 0.888
R20407 vss.n6610 vss.n5882 0.888
R20408 vss.n6610 vss.n5883 0.888
R20409 vss.n6558 vss.n5928 0.888
R20410 vss.n6558 vss.n5929 0.888
R20411 vss.n6484 vss.n5985 0.888
R20412 vss.n6484 vss.n6483 0.888
R20413 vss.n6431 vss.n6028 0.888
R20414 vss.n6431 vss.n6430 0.888
R20415 vss.n6363 vss.n6089 0.888
R20416 vss.n6363 vss.n6090 0.888
R20417 vss.n6311 vss.n6135 0.888
R20418 vss.n6311 vss.n6136 0.888
R20419 vss.n6237 vss.n6192 0.888
R20420 vss.n6237 vss.n6236 0.888
R20421 vss.n12900 vss.n12899 0.869
R20422 vss.n12635 vss.n12634 0.869
R20423 vss.n9154 vss.n8921 0.853
R20424 vss.n22728 vss.n22727 0.853
R20425 vss.n22737 vss.n22736 0.853
R20426 vss.n22659 vss.n22649 0.853
R20427 vss.n22651 vss.n22650 0.853
R20428 vss.n22520 vss.n22519 0.853
R20429 vss.n22529 vss.n22528 0.853
R20430 vss.n22451 vss.n22441 0.853
R20431 vss.n22443 vss.n22442 0.853
R20432 vss.n22312 vss.n22311 0.853
R20433 vss.n22321 vss.n22320 0.853
R20434 vss.n22243 vss.n22233 0.853
R20435 vss.n22235 vss.n22234 0.853
R20436 vss.n22104 vss.n22103 0.853
R20437 vss.n22113 vss.n22112 0.853
R20438 vss.n17408 vss.n17398 0.853
R20439 vss.n17400 vss.n17399 0.853
R20440 vss.n21448 vss.n21447 0.853
R20441 vss.n21457 vss.n21456 0.853
R20442 vss.n21379 vss.n21369 0.853
R20443 vss.n21371 vss.n21370 0.853
R20444 vss.n21240 vss.n21239 0.853
R20445 vss.n21249 vss.n21248 0.853
R20446 vss.n21171 vss.n21161 0.853
R20447 vss.n21163 vss.n21162 0.853
R20448 vss.n21032 vss.n21031 0.853
R20449 vss.n21041 vss.n21040 0.853
R20450 vss.n20963 vss.n20953 0.853
R20451 vss.n20955 vss.n20954 0.853
R20452 vss.n8891 vss.n8890 0.853
R20453 vss.n8900 vss.n8899 0.853
R20454 vss.n8822 vss.n8812 0.853
R20455 vss.n8814 vss.n8813 0.853
R20456 vss.n8683 vss.n8682 0.853
R20457 vss.n8692 vss.n8691 0.853
R20458 vss.n8614 vss.n8604 0.853
R20459 vss.n8606 vss.n8605 0.853
R20460 vss.n8475 vss.n8474 0.853
R20461 vss.n8484 vss.n8483 0.853
R20462 vss.n8406 vss.n8396 0.853
R20463 vss.n8398 vss.n8397 0.853
R20464 vss.n8267 vss.n8266 0.853
R20465 vss.n8276 vss.n8275 0.853
R20466 vss.n8198 vss.n8188 0.853
R20467 vss.n8190 vss.n8189 0.853
R20468 vss.n8059 vss.n8058 0.853
R20469 vss.n8068 vss.n8067 0.853
R20470 vss.n7990 vss.n7980 0.853
R20471 vss.n7982 vss.n7981 0.853
R20472 vss.n7851 vss.n7850 0.853
R20473 vss.n7860 vss.n7859 0.853
R20474 vss.n7781 vss.n7771 0.853
R20475 vss.n7773 vss.n7772 0.853
R20476 vss.n7642 vss.n7641 0.853
R20477 vss.n7651 vss.n7650 0.853
R20478 vss.n7573 vss.n7563 0.853
R20479 vss.n7565 vss.n7564 0.853
R20480 vss.n17575 vss.n17558 0.835
R20481 vss.n4185 vss.n4168 0.835
R20482 vss.n17275 vss.n17274 0.835
R20483 vss.n10558 vss.n10557 0.829
R20484 vss.n12343 vss.n12342 0.829
R20485 vss.n13767 vss.n13766 0.829
R20486 vss.n11503 vss.n11502 0.829
R20487 vss.n14978 vss.n14977 0.823
R20488 vss.n13140 vss.n13139 0.823
R20489 vss.n11473 vss.n11472 0.823
R20490 vss.n11691 vss.n11690 0.823
R20491 vss.n13113 vss.n13112 0.823
R20492 vss.n13662 vss.n13661 0.823
R20493 vss.n12405 vss.n12404 0.823
R20494 vss.n10668 vss.n10667 0.823
R20495 vss.n12322 vss.n12321 0.823
R20496 vss.n11483 vss.n11482 0.823
R20497 vss.n13371 vss.n13370 0.823
R20498 vss.n10804 vss.n10803 0.823
R20499 vss.n14559 vss.n14558 0.823
R20500 vss.n10929 vss.n10928 0.823
R20501 vss.n13649 vss.n13648 0.823
R20502 vss.n14058 vss.n14057 0.823
R20503 vss.n9153 vss.n9152 0.818
R20504 vss.n12540 vss.n12538 0.81
R20505 vss.n12774 vss.n12772 0.81
R20506 vss.n9126 vss.n9125 0.807
R20507 vss.n18987 vss.n17655 0.8
R20508 vss.n18982 vss.n17656 0.8
R20509 vss.n17711 vss.n17710 0.8
R20510 vss.n17715 vss.n17712 0.8
R20511 vss.n18865 vss.n17758 0.8
R20512 vss.n18858 vss.n17762 0.8
R20513 vss.n18799 vss.n18798 0.8
R20514 vss.n18791 vss.n17816 0.8
R20515 vss.n17865 vss.n17864 0.8
R20516 vss.n17874 vss.n17866 0.8
R20517 vss.n17924 vss.n17923 0.8
R20518 vss.n17928 vss.n17925 0.8
R20519 vss.n18624 vss.n17971 0.8
R20520 vss.n18617 vss.n17975 0.8
R20521 vss.n18558 vss.n18557 0.8
R20522 vss.n18550 vss.n18029 0.8
R20523 vss.n18078 vss.n18077 0.8
R20524 vss.n18087 vss.n18079 0.8
R20525 vss.n18137 vss.n18136 0.8
R20526 vss.n18141 vss.n18138 0.8
R20527 vss.n18383 vss.n18184 0.8
R20528 vss.n18376 vss.n18188 0.8
R20529 vss.n18317 vss.n18316 0.8
R20530 vss.n18309 vss.n18242 0.8
R20531 vss.n20258 vss.n19058 0.8
R20532 vss.n20251 vss.n19062 0.8
R20533 vss.n20192 vss.n20191 0.8
R20534 vss.n20184 vss.n19116 0.8
R20535 vss.n20133 vss.n19162 0.8
R20536 vss.n20128 vss.n19163 0.8
R20537 vss.n19218 vss.n19217 0.8
R20538 vss.n19222 vss.n19219 0.8
R20539 vss.n20011 vss.n19265 0.8
R20540 vss.n20004 vss.n19269 0.8
R20541 vss.n19945 vss.n19944 0.8
R20542 vss.n19937 vss.n19323 0.8
R20543 vss.n19886 vss.n19369 0.8
R20544 vss.n19881 vss.n19370 0.8
R20545 vss.n19425 vss.n19424 0.8
R20546 vss.n19429 vss.n19426 0.8
R20547 vss.n19764 vss.n19472 0.8
R20548 vss.n19757 vss.n19476 0.8
R20549 vss.n19698 vss.n19697 0.8
R20550 vss.n19690 vss.n19530 0.8
R20551 vss.n19639 vss.n19576 0.8
R20552 vss.n19634 vss.n19577 0.8
R20553 vss.n19619 vss.n19618 0.8
R20554 vss.n5597 vss.n4265 0.8
R20555 vss.n5592 vss.n4266 0.8
R20556 vss.n4321 vss.n4320 0.8
R20557 vss.n4325 vss.n4322 0.8
R20558 vss.n5475 vss.n4368 0.8
R20559 vss.n5468 vss.n4372 0.8
R20560 vss.n5409 vss.n5408 0.8
R20561 vss.n5401 vss.n4426 0.8
R20562 vss.n4475 vss.n4474 0.8
R20563 vss.n4484 vss.n4476 0.8
R20564 vss.n4534 vss.n4533 0.8
R20565 vss.n4538 vss.n4535 0.8
R20566 vss.n5234 vss.n4581 0.8
R20567 vss.n5227 vss.n4585 0.8
R20568 vss.n5168 vss.n5167 0.8
R20569 vss.n5160 vss.n4639 0.8
R20570 vss.n4688 vss.n4687 0.8
R20571 vss.n4697 vss.n4689 0.8
R20572 vss.n4747 vss.n4746 0.8
R20573 vss.n4751 vss.n4748 0.8
R20574 vss.n4993 vss.n4794 0.8
R20575 vss.n4986 vss.n4798 0.8
R20576 vss.n4927 vss.n4926 0.8
R20577 vss.n4919 vss.n4852 0.8
R20578 vss.n6868 vss.n5668 0.8
R20579 vss.n6861 vss.n5672 0.8
R20580 vss.n6802 vss.n6801 0.8
R20581 vss.n6794 vss.n5726 0.8
R20582 vss.n6743 vss.n5772 0.8
R20583 vss.n6738 vss.n5773 0.8
R20584 vss.n5828 vss.n5827 0.8
R20585 vss.n5832 vss.n5829 0.8
R20586 vss.n6621 vss.n5875 0.8
R20587 vss.n6614 vss.n5879 0.8
R20588 vss.n6555 vss.n6554 0.8
R20589 vss.n6547 vss.n5933 0.8
R20590 vss.n6496 vss.n5979 0.8
R20591 vss.n6491 vss.n5980 0.8
R20592 vss.n6035 vss.n6034 0.8
R20593 vss.n6039 vss.n6036 0.8
R20594 vss.n6374 vss.n6082 0.8
R20595 vss.n6367 vss.n6086 0.8
R20596 vss.n6308 vss.n6307 0.8
R20597 vss.n6300 vss.n6140 0.8
R20598 vss.n6249 vss.n6186 0.8
R20599 vss.n6244 vss.n6187 0.8
R20600 vss.n6229 vss.n6228 0.8
R20601 vss.n9095 vss.n9094 0.796
R20602 vss.n12587 vss.n12586 0.793
R20603 vss.n12429 vss.n12428 0.793
R20604 vss.n13302 vss.n13301 0.793
R20605 vss.n14404 vss.n14401 0.792
R20606 vss.n11056 vss.n11053 0.792
R20607 vss.n9003 vss.n9002 0.785
R20608 vss.n9064 vss.n9063 0.782
R20609 vss.n9660 vss.n9659 0.78
R20610 vss.n9033 vss.n9032 0.777
R20611 vss.n21795 vss.n21794 0.768
R20612 vss.n3744 vss.n3743 0.768
R20613 vss.n16329 vss.n16322 0.768
R20614 vss.n16406 vss.n16399 0.768
R20615 vss.n16565 vss.n16558 0.768
R20616 vss.n16642 vss.n16635 0.768
R20617 vss.n16711 vss.n16702 0.768
R20618 vss.n16752 vss.n16751 0.768
R20619 vss.n16825 vss.n16824 0.768
R20620 vss.n16862 vss.n16861 0.768
R20621 vss.n16941 vss.n16932 0.768
R20622 vss.n16982 vss.n16981 0.768
R20623 vss.n17061 vss.n17060 0.768
R20624 vss.n17098 vss.n17097 0.768
R20625 vss.n17177 vss.n17168 0.768
R20626 vss.n17218 vss.n17217 0.768
R20627 vss.n17315 vss.n17314 0.768
R20628 vss.n15906 vss.n15899 0.768
R20629 vss.n15986 vss.n15979 0.768
R20630 vss.n16030 vss.n16029 0.768
R20631 vss.n16115 vss.n16105 0.768
R20632 vss.n16142 vss.n16135 0.768
R20633 vss.n16222 vss.n16215 0.768
R20634 vss.n15258 vss.n15251 0.768
R20635 vss.n15382 vss.n15375 0.768
R20636 vss.n15459 vss.n15452 0.768
R20637 vss.n15618 vss.n15611 0.768
R20638 vss.n15695 vss.n15688 0.768
R20639 vss.n15846 vss.n15839 0.768
R20640 vss.n22032 vss.n21997 0.766
R20641 vss.n3981 vss.n3946 0.766
R20642 vss.n14459 vss.n14452 0.76
R20643 vss.n14641 vss.n14634 0.76
R20644 vss.n13563 vss.n13556 0.76
R20645 vss.n14754 vss.n14747 0.76
R20646 vss.n14921 vss.n14914 0.76
R20647 vss.n14949 vss.n14942 0.76
R20648 vss.n15034 vss.n15027 0.76
R20649 vss.n10479 vss.n10472 0.76
R20650 vss.n14328 vss.n14321 0.76
R20651 vss.n13901 vss.n13894 0.76
R20652 vss.n11737 vss.n11730 0.76
R20653 vss.n14002 vss.n13995 0.76
R20654 vss.n11594 vss.n11587 0.76
R20655 vss.n12214 vss.n12207 0.76
R20656 vss.n12456 vss.n12449 0.76
R20657 vss.n12618 vss.n12611 0.76
R20658 vss.n10847 vss.n10840 0.76
R20659 vss.n10891 vss.n10884 0.76
R20660 vss.n11247 vss.n11240 0.76
R20661 vss.n11212 vss.n11205 0.76
R20662 vss.n20522 vss.n20521 0.752
R20663 vss.n20549 vss.n20548 0.752
R20664 vss.n20751 vss.n20750 0.752
R20665 vss.n20771 vss.n20770 0.752
R20666 vss.n20315 vss.n20314 0.752
R20667 vss.n20305 vss.n20304 0.752
R20668 vss.n21813 vss.n21812 0.752
R20669 vss.n21741 vss.n21740 0.752
R20670 vss.n12114 vss.n12113 0.752
R20671 vss.n12124 vss.n12123 0.752
R20672 vss.n10874 vss.n10873 0.752
R20673 vss.n11942 vss.n11941 0.752
R20674 vss.n14413 vss.n14412 0.752
R20675 vss.n14367 vss.n14366 0.752
R20676 vss.n11631 vss.n11630 0.752
R20677 vss.n11658 vss.n11657 0.752
R20678 vss.n13268 vss.n13267 0.752
R20679 vss.n13252 vss.n13251 0.752
R20680 vss.n13537 vss.n13536 0.752
R20681 vss.n14589 vss.n14588 0.752
R20682 vss.n14829 vss.n14828 0.752
R20683 vss.n14839 vss.n14838 0.752
R20684 vss.n14854 vss.n14853 0.752
R20685 vss.n14857 vss.n14856 0.752
R20686 vss.n10482 vss.n10481 0.752
R20687 vss.n10512 vss.n10511 0.752
R20688 vss.n3762 vss.n3761 0.752
R20689 vss.n3690 vss.n3689 0.752
R20690 vss.n7132 vss.n7131 0.752
R20691 vss.n7159 vss.n7158 0.752
R20692 vss.n7361 vss.n7360 0.752
R20693 vss.n7381 vss.n7380 0.752
R20694 vss.n6925 vss.n6924 0.752
R20695 vss.n6915 vss.n6914 0.752
R20696 vss.n1748 vss.n1747 0.752
R20697 vss.n1768 vss.n1767 0.752
R20698 vss.n1977 vss.n1976 0.752
R20699 vss.n2006 vss.n2005 0.752
R20700 vss.n2222 vss.n2221 0.752
R20701 vss.n2250 vss.n2249 0.752
R20702 vss.n2466 vss.n2465 0.752
R20703 vss.n2494 vss.n2493 0.752
R20704 vss.n2711 vss.n2710 0.752
R20705 vss.n2739 vss.n2738 0.752
R20706 vss.n2949 vss.n2948 0.752
R20707 vss.n2977 vss.n2976 0.752
R20708 vss.n3193 vss.n3192 0.752
R20709 vss.n3222 vss.n3221 0.752
R20710 vss.n15197 vss.n15196 0.752
R20711 vss.n15177 vss.n15176 0.752
R20712 vss.n209 vss.n208 0.752
R20713 vss.n229 vss.n228 0.752
R20714 vss.n438 vss.n437 0.752
R20715 vss.n467 vss.n466 0.752
R20716 vss.n683 vss.n682 0.752
R20717 vss.n711 vss.n710 0.752
R20718 vss.n927 vss.n926 0.752
R20719 vss.n955 vss.n954 0.752
R20720 vss.n1172 vss.n1171 0.752
R20721 vss.n1200 vss.n1199 0.752
R20722 vss.n23295 vss.n23294 0.752
R20723 vss.n23267 vss.n23266 0.752
R20724 vss.n23051 vss.n23050 0.752
R20725 vss.n23022 vss.n23021 0.752
R20726 vss.n1390 vss.n1389 0.752
R20727 vss.n22811 vss.n22810 0.752
R20728 vss.n8972 vss.n8971 0.742
R20729 vss.n21772 vss.n21760 0.739
R20730 vss.n3721 vss.n3709 0.739
R20731 vss.n10276 vss.n10275 0.723
R20732 vss.n22617 vss.n22616 0.711
R20733 vss.n22616 vss.n22609 0.711
R20734 vss.n22569 vss.n22562 0.711
R20735 vss.n22571 vss.n22569 0.711
R20736 vss.n22409 vss.n22408 0.711
R20737 vss.n22408 vss.n22401 0.711
R20738 vss.n22361 vss.n22354 0.711
R20739 vss.n22363 vss.n22361 0.711
R20740 vss.n22201 vss.n22200 0.711
R20741 vss.n22200 vss.n22193 0.711
R20742 vss.n22153 vss.n22146 0.711
R20743 vss.n22155 vss.n22153 0.711
R20744 vss.n21545 vss.n21544 0.711
R20745 vss.n21544 vss.n21537 0.711
R20746 vss.n21497 vss.n21490 0.711
R20747 vss.n21499 vss.n21497 0.711
R20748 vss.n21337 vss.n21336 0.711
R20749 vss.n21336 vss.n21329 0.711
R20750 vss.n21289 vss.n21282 0.711
R20751 vss.n21291 vss.n21289 0.711
R20752 vss.n21129 vss.n21128 0.711
R20753 vss.n21128 vss.n21121 0.711
R20754 vss.n21081 vss.n21074 0.711
R20755 vss.n21083 vss.n21081 0.711
R20756 vss.n20921 vss.n20920 0.711
R20757 vss.n20920 vss.n20913 0.711
R20758 vss.n18987 vss.n18986 0.711
R20759 vss.n18986 vss.n17656 0.711
R20760 vss.n18915 vss.n17711 0.711
R20761 vss.n18915 vss.n17712 0.711
R20762 vss.n18859 vss.n17758 0.711
R20763 vss.n18859 vss.n18858 0.711
R20764 vss.n18798 vss.n18797 0.711
R20765 vss.n18797 vss.n17816 0.711
R20766 vss.n18741 vss.n17865 0.711
R20767 vss.n18741 vss.n17866 0.711
R20768 vss.n18674 vss.n17924 0.711
R20769 vss.n18674 vss.n17925 0.711
R20770 vss.n18618 vss.n17971 0.711
R20771 vss.n18618 vss.n18617 0.711
R20772 vss.n18557 vss.n18556 0.711
R20773 vss.n18556 vss.n18029 0.711
R20774 vss.n18500 vss.n18078 0.711
R20775 vss.n18500 vss.n18079 0.711
R20776 vss.n18433 vss.n18137 0.711
R20777 vss.n18433 vss.n18138 0.711
R20778 vss.n18377 vss.n18184 0.711
R20779 vss.n18377 vss.n18376 0.711
R20780 vss.n18316 vss.n18315 0.711
R20781 vss.n18315 vss.n18242 0.711
R20782 vss.n20252 vss.n19058 0.711
R20783 vss.n20252 vss.n20251 0.711
R20784 vss.n20191 vss.n20190 0.711
R20785 vss.n20190 vss.n19116 0.711
R20786 vss.n20133 vss.n20132 0.711
R20787 vss.n20132 vss.n19163 0.711
R20788 vss.n20061 vss.n19218 0.711
R20789 vss.n20061 vss.n19219 0.711
R20790 vss.n20005 vss.n19265 0.711
R20791 vss.n20005 vss.n20004 0.711
R20792 vss.n19944 vss.n19943 0.711
R20793 vss.n19943 vss.n19323 0.711
R20794 vss.n19886 vss.n19885 0.711
R20795 vss.n19885 vss.n19370 0.711
R20796 vss.n19814 vss.n19425 0.711
R20797 vss.n19814 vss.n19426 0.711
R20798 vss.n19758 vss.n19472 0.711
R20799 vss.n19758 vss.n19757 0.711
R20800 vss.n19697 vss.n19696 0.711
R20801 vss.n19696 vss.n19530 0.711
R20802 vss.n19639 vss.n19638 0.711
R20803 vss.n19638 vss.n19577 0.711
R20804 vss.n5597 vss.n5596 0.711
R20805 vss.n5596 vss.n4266 0.711
R20806 vss.n5525 vss.n4321 0.711
R20807 vss.n5525 vss.n4322 0.711
R20808 vss.n5469 vss.n4368 0.711
R20809 vss.n5469 vss.n5468 0.711
R20810 vss.n5408 vss.n5407 0.711
R20811 vss.n5407 vss.n4426 0.711
R20812 vss.n5351 vss.n4475 0.711
R20813 vss.n5351 vss.n4476 0.711
R20814 vss.n5284 vss.n4534 0.711
R20815 vss.n5284 vss.n4535 0.711
R20816 vss.n5228 vss.n4581 0.711
R20817 vss.n5228 vss.n5227 0.711
R20818 vss.n5167 vss.n5166 0.711
R20819 vss.n5166 vss.n4639 0.711
R20820 vss.n5110 vss.n4688 0.711
R20821 vss.n5110 vss.n4689 0.711
R20822 vss.n5043 vss.n4747 0.711
R20823 vss.n5043 vss.n4748 0.711
R20824 vss.n4987 vss.n4794 0.711
R20825 vss.n4987 vss.n4986 0.711
R20826 vss.n4926 vss.n4925 0.711
R20827 vss.n4925 vss.n4852 0.711
R20828 vss.n6862 vss.n5668 0.711
R20829 vss.n6862 vss.n6861 0.711
R20830 vss.n6801 vss.n6800 0.711
R20831 vss.n6800 vss.n5726 0.711
R20832 vss.n6743 vss.n6742 0.711
R20833 vss.n6742 vss.n5773 0.711
R20834 vss.n6671 vss.n5828 0.711
R20835 vss.n6671 vss.n5829 0.711
R20836 vss.n6615 vss.n5875 0.711
R20837 vss.n6615 vss.n6614 0.711
R20838 vss.n6554 vss.n6553 0.711
R20839 vss.n6553 vss.n5933 0.711
R20840 vss.n6496 vss.n6495 0.711
R20841 vss.n6495 vss.n5980 0.711
R20842 vss.n6424 vss.n6035 0.711
R20843 vss.n6424 vss.n6036 0.711
R20844 vss.n6368 vss.n6082 0.711
R20845 vss.n6368 vss.n6367 0.711
R20846 vss.n6307 vss.n6306 0.711
R20847 vss.n6306 vss.n6140 0.711
R20848 vss.n6249 vss.n6248 0.711
R20849 vss.n6248 vss.n6187 0.711
R20850 vss.n8780 vss.n8779 0.711
R20851 vss.n8779 vss.n8772 0.711
R20852 vss.n8732 vss.n8725 0.711
R20853 vss.n8734 vss.n8732 0.711
R20854 vss.n8572 vss.n8571 0.711
R20855 vss.n8571 vss.n8564 0.711
R20856 vss.n8524 vss.n8517 0.711
R20857 vss.n8526 vss.n8524 0.711
R20858 vss.n8364 vss.n8363 0.711
R20859 vss.n8363 vss.n8356 0.711
R20860 vss.n8316 vss.n8309 0.711
R20861 vss.n8318 vss.n8316 0.711
R20862 vss.n8156 vss.n8155 0.711
R20863 vss.n8155 vss.n8148 0.711
R20864 vss.n8108 vss.n8101 0.711
R20865 vss.n8110 vss.n8108 0.711
R20866 vss.n7948 vss.n7947 0.711
R20867 vss.n7947 vss.n7940 0.711
R20868 vss.n7900 vss.n7893 0.711
R20869 vss.n7902 vss.n7900 0.711
R20870 vss.n7739 vss.n7738 0.711
R20871 vss.n7738 vss.n7731 0.711
R20872 vss.n7691 vss.n7684 0.711
R20873 vss.n7693 vss.n7691 0.711
R20874 vss.n7531 vss.n7530 0.711
R20875 vss.n7530 vss.n7523 0.711
R20876 vss.n12569 vss.n12568 0.71
R20877 vss.n13290 vss.n13289 0.71
R20878 vss.n14392 vss.n14391 0.709
R20879 vss.n11044 vss.n11043 0.709
R20880 vss.n12468 vss.n12467 0.704
R20881 vss.n8964 vss.n8963 0.699
R20882 vss.n10320 vss.n10319 0.698
R20883 vss.n12943 vss.n12942 0.697
R20884 vss.n13163 vss.n13162 0.697
R20885 vss.n13154 vss.n13153 0.697
R20886 vss.n11545 vss.n11544 0.697
R20887 vss.n11543 vss.n11542 0.697
R20888 vss.n11514 vss.n11513 0.697
R20889 vss.n12984 vss.n12983 0.697
R20890 vss.n12974 vss.n12973 0.697
R20891 vss.n12384 vss.n12383 0.697
R20892 vss.n12357 vss.n12356 0.697
R20893 vss.n10688 vss.n10687 0.697
R20894 vss.n10698 vss.n10697 0.697
R20895 vss.n13411 vss.n13410 0.697
R20896 vss.n13490 vss.n13489 0.697
R20897 vss.n13070 vss.n13069 0.697
R20898 vss.n10623 vss.n10622 0.697
R20899 vss.n10783 vss.n10782 0.697
R20900 vss.n12291 vss.n12290 0.697
R20901 vss.n14155 vss.n14154 0.697
R20902 vss.n14112 vss.n14111 0.697
R20903 vss.n13731 vss.n13730 0.697
R20904 vss.n11428 vss.n11427 0.697
R20905 vss.n11868 vss.n11867 0.697
R20906 vss.n11904 vss.n11903 0.697
R20907 vss.n13778 vss.n13777 0.697
R20908 vss.n13789 vss.n13788 0.697
R20909 vss.n21984 vss.n21983 0.697
R20910 vss.n21613 vss.n21612 0.697
R20911 vss.n3933 vss.n3932 0.697
R20912 vss.n3562 vss.n3561 0.697
R20913 vss.n10295 vss.n10294 0.693
R20914 vss.n19032 vss.n19031 0.692
R20915 vss.n5642 vss.n5641 0.692
R20916 vss.n9196 vss.n9194 0.683
R20917 vss.n15098 vss.t350 0.671
R20918 vss.n15109 vss.t345 0.671
R20919 vss.t328 vss.n9197 0.669
R20920 vss.n21620 vss.n21619 0.649
R20921 vss.n3569 vss.n3568 0.649
R20922 vss.n16441 vss.n16440 0.64
R20923 vss.n16516 vss.n16515 0.64
R20924 vss.n16711 vss.n16710 0.64
R20925 vss.n16744 vss.n16743 0.64
R20926 vss.n16813 vss.n16812 0.64
R20927 vss.n16876 vss.n16867 0.64
R20928 vss.n16941 vss.n16940 0.64
R20929 vss.n16974 vss.n16973 0.64
R20930 vss.n17055 vss.n17054 0.64
R20931 vss.n17112 vss.n17103 0.64
R20932 vss.n17177 vss.n17176 0.64
R20933 vss.n17210 vss.n17209 0.64
R20934 vss.n17298 vss.n17297 0.64
R20935 vss.n15921 vss.n15920 0.64
R20936 vss.n15988 vss.n15986 0.64
R20937 vss.n16021 vss.n16020 0.64
R20938 vss.n16093 vss.n16092 0.64
R20939 vss.n16157 vss.n16156 0.64
R20940 vss.n16224 vss.n16222 0.64
R20941 vss.n15293 vss.n15292 0.64
R20942 vss.n15332 vss.n15331 0.64
R20943 vss.n15494 vss.n15493 0.64
R20944 vss.n15569 vss.n15568 0.64
R20945 vss.n15730 vss.n15729 0.64
R20946 vss.n15797 vss.n15796 0.64
R20947 vss.n15099 vss.n15098 0.628
R20948 vss.n15100 vss.n15099 0.628
R20949 vss.n15101 vss.n15100 0.628
R20950 vss.n15102 vss.n15101 0.628
R20951 vss.n15103 vss.n15102 0.628
R20952 vss.n15104 vss.n15103 0.628
R20953 vss.n15105 vss.n15104 0.628
R20954 vss.n15106 vss.n15105 0.628
R20955 vss.n15107 vss.n15106 0.628
R20956 vss.n15108 vss.n15107 0.628
R20957 vss.n15110 vss.n15109 0.628
R20958 vss.n15111 vss.n15110 0.628
R20959 vss.n15112 vss.n15111 0.628
R20960 vss.n15113 vss.n15112 0.628
R20961 vss.n15114 vss.n15113 0.628
R20962 vss.n15115 vss.n15114 0.628
R20963 vss.n15116 vss.n15115 0.628
R20964 vss.n15117 vss.n15116 0.628
R20965 vss.n15118 vss.n15117 0.628
R20966 vss.n15119 vss.n15118 0.628
R20967 vss.n18981 vss.n17661 0.622
R20968 vss.n18974 vss.n17665 0.622
R20969 vss.n18926 vss.n17704 0.622
R20970 vss.n18921 vss.n17706 0.622
R20971 vss.n17765 vss.n17764 0.622
R20972 vss.n17774 vss.n17766 0.622
R20973 vss.n17811 vss.n17810 0.622
R20974 vss.n17815 vss.n17812 0.622
R20975 vss.n18735 vss.n17872 0.622
R20976 vss.n18730 vss.n17873 0.622
R20977 vss.n18685 vss.n17917 0.622
R20978 vss.n18680 vss.n17919 0.622
R20979 vss.n17978 vss.n17977 0.622
R20980 vss.n17987 vss.n17979 0.622
R20981 vss.n18024 vss.n18023 0.622
R20982 vss.n18028 vss.n18025 0.622
R20983 vss.n18494 vss.n18085 0.622
R20984 vss.n18489 vss.n18086 0.622
R20985 vss.n18444 vss.n18130 0.622
R20986 vss.n18439 vss.n18132 0.622
R20987 vss.n18191 vss.n18190 0.622
R20988 vss.n18200 vss.n18192 0.622
R20989 vss.n18237 vss.n18236 0.622
R20990 vss.n18241 vss.n18238 0.622
R20991 vss.n19612 vss.n19594 0.622
R20992 vss.n19065 vss.n19064 0.622
R20993 vss.n19074 vss.n19066 0.622
R20994 vss.n19111 vss.n19110 0.622
R20995 vss.n19115 vss.n19112 0.622
R20996 vss.n20127 vss.n19168 0.622
R20997 vss.n20120 vss.n19172 0.622
R20998 vss.n20072 vss.n19211 0.622
R20999 vss.n20067 vss.n19213 0.622
R21000 vss.n19272 vss.n19271 0.622
R21001 vss.n19281 vss.n19273 0.622
R21002 vss.n19318 vss.n19317 0.622
R21003 vss.n19322 vss.n19319 0.622
R21004 vss.n19880 vss.n19375 0.622
R21005 vss.n19873 vss.n19379 0.622
R21006 vss.n19825 vss.n19418 0.622
R21007 vss.n19820 vss.n19420 0.622
R21008 vss.n19479 vss.n19478 0.622
R21009 vss.n19488 vss.n19480 0.622
R21010 vss.n19525 vss.n19524 0.622
R21011 vss.n19529 vss.n19526 0.622
R21012 vss.n19633 vss.n19582 0.622
R21013 vss.n19626 vss.n19586 0.622
R21014 vss.n5591 vss.n4271 0.622
R21015 vss.n5584 vss.n4275 0.622
R21016 vss.n5536 vss.n4314 0.622
R21017 vss.n5531 vss.n4316 0.622
R21018 vss.n4375 vss.n4374 0.622
R21019 vss.n4384 vss.n4376 0.622
R21020 vss.n4421 vss.n4420 0.622
R21021 vss.n4425 vss.n4422 0.622
R21022 vss.n5345 vss.n4482 0.622
R21023 vss.n5340 vss.n4483 0.622
R21024 vss.n5295 vss.n4527 0.622
R21025 vss.n5290 vss.n4529 0.622
R21026 vss.n4588 vss.n4587 0.622
R21027 vss.n4597 vss.n4589 0.622
R21028 vss.n4634 vss.n4633 0.622
R21029 vss.n4638 vss.n4635 0.622
R21030 vss.n5104 vss.n4695 0.622
R21031 vss.n5099 vss.n4696 0.622
R21032 vss.n5054 vss.n4740 0.622
R21033 vss.n5049 vss.n4742 0.622
R21034 vss.n4801 vss.n4800 0.622
R21035 vss.n4810 vss.n4802 0.622
R21036 vss.n4847 vss.n4846 0.622
R21037 vss.n4851 vss.n4848 0.622
R21038 vss.n6222 vss.n6204 0.622
R21039 vss.n5675 vss.n5674 0.622
R21040 vss.n5684 vss.n5676 0.622
R21041 vss.n5721 vss.n5720 0.622
R21042 vss.n5725 vss.n5722 0.622
R21043 vss.n6737 vss.n5778 0.622
R21044 vss.n6730 vss.n5782 0.622
R21045 vss.n6682 vss.n5821 0.622
R21046 vss.n6677 vss.n5823 0.622
R21047 vss.n5882 vss.n5881 0.622
R21048 vss.n5891 vss.n5883 0.622
R21049 vss.n5928 vss.n5927 0.622
R21050 vss.n5932 vss.n5929 0.622
R21051 vss.n6490 vss.n5985 0.622
R21052 vss.n6483 vss.n5989 0.622
R21053 vss.n6435 vss.n6028 0.622
R21054 vss.n6430 vss.n6030 0.622
R21055 vss.n6089 vss.n6088 0.622
R21056 vss.n6098 vss.n6090 0.622
R21057 vss.n6135 vss.n6134 0.622
R21058 vss.n6139 vss.n6136 0.622
R21059 vss.n6243 vss.n6192 0.622
R21060 vss.n6236 vss.n6196 0.622
R21061 vss.n9193 vss.n9192 0.615
R21062 vss.n9060 vss.n9059 0.604
R21063 vss.n14820 vss.n13250 0.595
R21064 vss.n12147 vss.n12136 0.595
R21065 vss.t1 vss.n9202 0.58
R21066 vss.n22714 vss.n22713 0.568
R21067 vss.n22723 vss.n22722 0.568
R21068 vss.n22673 vss.n22663 0.568
R21069 vss.n22665 vss.n22664 0.568
R21070 vss.n22506 vss.n22505 0.568
R21071 vss.n22515 vss.n22514 0.568
R21072 vss.n22465 vss.n22455 0.568
R21073 vss.n22457 vss.n22456 0.568
R21074 vss.n22298 vss.n22297 0.568
R21075 vss.n22307 vss.n22306 0.568
R21076 vss.n22257 vss.n22247 0.568
R21077 vss.n22249 vss.n22248 0.568
R21078 vss.n22090 vss.n22089 0.568
R21079 vss.n22099 vss.n22098 0.568
R21080 vss.n21581 vss.n21580 0.568
R21081 vss.n21434 vss.n21433 0.568
R21082 vss.n21443 vss.n21442 0.568
R21083 vss.n21393 vss.n21383 0.568
R21084 vss.n21385 vss.n21384 0.568
R21085 vss.n21226 vss.n21225 0.568
R21086 vss.n21235 vss.n21234 0.568
R21087 vss.n21185 vss.n21175 0.568
R21088 vss.n21177 vss.n21176 0.568
R21089 vss.n21018 vss.n21017 0.568
R21090 vss.n21027 vss.n21026 0.568
R21091 vss.n20977 vss.n20967 0.568
R21092 vss.n20969 vss.n20968 0.568
R21093 vss.n8877 vss.n8876 0.568
R21094 vss.n8886 vss.n8885 0.568
R21095 vss.n8836 vss.n8826 0.568
R21096 vss.n8828 vss.n8827 0.568
R21097 vss.n8669 vss.n8668 0.568
R21098 vss.n8678 vss.n8677 0.568
R21099 vss.n8628 vss.n8618 0.568
R21100 vss.n8620 vss.n8619 0.568
R21101 vss.n8461 vss.n8460 0.568
R21102 vss.n8470 vss.n8469 0.568
R21103 vss.n8420 vss.n8410 0.568
R21104 vss.n8412 vss.n8411 0.568
R21105 vss.n8253 vss.n8252 0.568
R21106 vss.n8262 vss.n8261 0.568
R21107 vss.n8212 vss.n8202 0.568
R21108 vss.n8204 vss.n8203 0.568
R21109 vss.n8045 vss.n8044 0.568
R21110 vss.n8054 vss.n8053 0.568
R21111 vss.n8004 vss.n7994 0.568
R21112 vss.n7996 vss.n7995 0.568
R21113 vss.n7836 vss.n7835 0.568
R21114 vss.n7845 vss.n7844 0.568
R21115 vss.n7795 vss.n7785 0.568
R21116 vss.n7787 vss.n7786 0.568
R21117 vss.n7628 vss.n7627 0.568
R21118 vss.n7637 vss.n7636 0.568
R21119 vss.n7587 vss.n7577 0.568
R21120 vss.n7579 vss.n7578 0.568
R21121 vss.n9195 vss.t220 0.567
R21122 vss.n9194 vss.t221 0.567
R21123 vss.n8929 vss.n8927 0.565
R21124 vss.n18994 vss.n18993 0.533
R21125 vss.n18993 vss.n17647 0.533
R21126 vss.n18911 vss.n18910 0.533
R21127 vss.n18910 vss.n17716 0.533
R21128 vss.n18871 vss.n18870 0.533
R21129 vss.n18870 vss.n17754 0.533
R21130 vss.n18786 vss.n17823 0.533
R21131 vss.n18786 vss.n18785 0.533
R21132 vss.n18746 vss.n17858 0.533
R21133 vss.n18746 vss.n18745 0.533
R21134 vss.n18670 vss.n18669 0.533
R21135 vss.n18669 vss.n17929 0.533
R21136 vss.n18630 vss.n18629 0.533
R21137 vss.n18629 vss.n17967 0.533
R21138 vss.n18545 vss.n18036 0.533
R21139 vss.n18545 vss.n18544 0.533
R21140 vss.n18505 vss.n18071 0.533
R21141 vss.n18505 vss.n18504 0.533
R21142 vss.n18429 vss.n18428 0.533
R21143 vss.n18428 vss.n18142 0.533
R21144 vss.n18389 vss.n18388 0.533
R21145 vss.n18388 vss.n18180 0.533
R21146 vss.n18304 vss.n18249 0.533
R21147 vss.n18304 vss.n18303 0.533
R21148 vss.n19604 vss.n19594 0.533
R21149 vss.n20264 vss.n20263 0.533
R21150 vss.n20263 vss.n19053 0.533
R21151 vss.n20179 vss.n19123 0.533
R21152 vss.n20179 vss.n20178 0.533
R21153 vss.n20140 vss.n20139 0.533
R21154 vss.n20139 vss.n19154 0.533
R21155 vss.n20057 vss.n20056 0.533
R21156 vss.n20056 vss.n19223 0.533
R21157 vss.n20017 vss.n20016 0.533
R21158 vss.n20016 vss.n19261 0.533
R21159 vss.n19932 vss.n19330 0.533
R21160 vss.n19932 vss.n19931 0.533
R21161 vss.n19893 vss.n19892 0.533
R21162 vss.n19892 vss.n19361 0.533
R21163 vss.n19810 vss.n19809 0.533
R21164 vss.n19809 vss.n19430 0.533
R21165 vss.n19770 vss.n19769 0.533
R21166 vss.n19769 vss.n19468 0.533
R21167 vss.n19685 vss.n19537 0.533
R21168 vss.n19685 vss.n19684 0.533
R21169 vss.n19646 vss.n19645 0.533
R21170 vss.n19645 vss.n19568 0.533
R21171 vss.n11395 vss.n11389 0.533
R21172 vss.n13925 vss.n13920 0.533
R21173 vss.n13613 vss.n13607 0.533
R21174 vss.n11775 vss.n11774 0.533
R21175 vss.n11024 vss.n11019 0.533
R21176 vss.n11271 vss.n11266 0.533
R21177 vss.n10836 vss.n10832 0.533
R21178 vss.n12237 vss.n12232 0.533
R21179 vss.n12519 vss.n12513 0.533
R21180 vss.n10497 vss.n10492 0.533
R21181 vss.n13198 vss.n13193 0.533
R21182 vss.n13623 vss.n13617 0.533
R21183 vss.n13427 vss.n13422 0.533
R21184 vss.n13436 vss.n13431 0.533
R21185 vss.n10916 vss.n10912 0.533
R21186 vss.n10590 vss.n10585 0.533
R21187 vss.n11403 vss.n11399 0.533
R21188 vss.n10598 vss.n10594 0.533
R21189 vss.n14038 vss.n14037 0.533
R21190 vss.n11651 vss.n11646 0.533
R21191 vss.n5604 vss.n5603 0.533
R21192 vss.n5603 vss.n4257 0.533
R21193 vss.n5521 vss.n5520 0.533
R21194 vss.n5520 vss.n4326 0.533
R21195 vss.n5481 vss.n5480 0.533
R21196 vss.n5480 vss.n4364 0.533
R21197 vss.n5396 vss.n4433 0.533
R21198 vss.n5396 vss.n5395 0.533
R21199 vss.n5356 vss.n4468 0.533
R21200 vss.n5356 vss.n5355 0.533
R21201 vss.n5280 vss.n5279 0.533
R21202 vss.n5279 vss.n4539 0.533
R21203 vss.n5240 vss.n5239 0.533
R21204 vss.n5239 vss.n4577 0.533
R21205 vss.n5155 vss.n4646 0.533
R21206 vss.n5155 vss.n5154 0.533
R21207 vss.n5115 vss.n4681 0.533
R21208 vss.n5115 vss.n5114 0.533
R21209 vss.n5039 vss.n5038 0.533
R21210 vss.n5038 vss.n4752 0.533
R21211 vss.n4999 vss.n4998 0.533
R21212 vss.n4998 vss.n4790 0.533
R21213 vss.n4914 vss.n4859 0.533
R21214 vss.n4914 vss.n4913 0.533
R21215 vss.n6214 vss.n6204 0.533
R21216 vss.n6874 vss.n6873 0.533
R21217 vss.n6873 vss.n5663 0.533
R21218 vss.n6789 vss.n5733 0.533
R21219 vss.n6789 vss.n6788 0.533
R21220 vss.n6750 vss.n6749 0.533
R21221 vss.n6749 vss.n5764 0.533
R21222 vss.n6667 vss.n6666 0.533
R21223 vss.n6666 vss.n5833 0.533
R21224 vss.n6627 vss.n6626 0.533
R21225 vss.n6626 vss.n5871 0.533
R21226 vss.n6542 vss.n5940 0.533
R21227 vss.n6542 vss.n6541 0.533
R21228 vss.n6503 vss.n6502 0.533
R21229 vss.n6502 vss.n5971 0.533
R21230 vss.n6420 vss.n6419 0.533
R21231 vss.n6419 vss.n6040 0.533
R21232 vss.n6380 vss.n6379 0.533
R21233 vss.n6379 vss.n6078 0.533
R21234 vss.n6295 vss.n6147 0.533
R21235 vss.n6295 vss.n6294 0.533
R21236 vss.n6256 vss.n6255 0.533
R21237 vss.n6255 vss.n6178 0.533
R21238 vss.n12073 vss.n12072 0.533
R21239 vss.n10802 vss.n10801 0.533
R21240 vss.n10965 vss.n10964 0.533
R21241 vss.n11005 vss.n11004 0.533
R21242 vss.n11722 vss.n11721 0.533
R21243 vss.n14076 vss.n14075 0.533
R21244 vss.n13855 vss.n13854 0.533
R21245 vss.n13353 vss.n13352 0.533
R21246 vss.n14698 vss.n14697 0.533
R21247 vss.n14191 vss.n14190 0.533
R21248 vss.n9196 vss.n9195 0.517
R21249 vss.n16301 vss.n16296 0.512
R21250 vss.n16343 vss.n16336 0.512
R21251 vss.n16392 vss.n16385 0.512
R21252 vss.n16579 vss.n16572 0.512
R21253 vss.n16628 vss.n16621 0.512
R21254 vss.n16697 vss.n16688 0.512
R21255 vss.n16811 vss.n16810 0.512
R21256 vss.n16876 vss.n16875 0.512
R21257 vss.n16927 vss.n16918 0.512
R21258 vss.n16996 vss.n16995 0.512
R21259 vss.n17047 vss.n17046 0.512
R21260 vss.n17112 vss.n17111 0.512
R21261 vss.n17163 vss.n17154 0.512
R21262 vss.n17232 vss.n17231 0.512
R21263 vss.n15880 vss.n15875 0.512
R21264 vss.n15920 vss.n15913 0.512
R21265 vss.n15972 vss.n15965 0.512
R21266 vss.n16044 vss.n16043 0.512
R21267 vss.n16101 vss.n16091 0.512
R21268 vss.n16156 vss.n16149 0.512
R21269 vss.n16208 vss.n16201 0.512
R21270 vss.n16281 vss.n16274 0.512
R21271 vss.n15396 vss.n15389 0.512
R21272 vss.n15445 vss.n15438 0.512
R21273 vss.n15632 vss.n15625 0.512
R21274 vss.n15681 vss.n15674 0.512
R21275 vss.n15860 vss.n15853 0.512
R21276 vss.n10355 vss.n10354 0.509
R21277 vss.n10251 vss.n10250 0.508
R21278 vss.n10390 vss.n10389 0.507
R21279 vss.n14494 vss.n14487 0.506
R21280 vss.n14401 vss.n14394 0.506
R21281 vss.n14664 vss.n14657 0.506
R21282 vss.n13583 vss.n13576 0.506
R21283 vss.n13301 vss.n13294 0.506
R21284 vss.n13342 vss.n13335 0.506
R21285 vss.n13243 vss.n13236 0.506
R21286 vss.n14964 vss.n14957 0.506
R21287 vss.n15018 vss.n15011 0.506
R21288 vss.n10509 vss.n10502 0.506
R21289 vss.n14360 vss.n14353 0.506
R21290 vss.n13866 vss.n13859 0.506
R21291 vss.n11763 vss.n11756 0.506
R21292 vss.n11053 vss.n11046 0.506
R21293 vss.n11168 vss.n11163 0.506
R21294 vss.n13981 vss.n13974 0.506
R21295 vss.n11576 vss.n11569 0.506
R21296 vss.n12574 vss.n12573 0.506
R21297 vss.n12586 vss.n12579 0.506
R21298 vss.n12082 vss.n12075 0.506
R21299 vss.n12428 vss.n12421 0.506
R21300 vss.n12601 vss.n12594 0.506
R21301 vss.n10827 vss.n10820 0.506
R21302 vss.n10901 vss.n10894 0.506
R21303 vss.n10954 vss.n10947 0.506
R21304 vss.n11014 vss.n11007 0.506
R21305 vss.n17274 vss.n17273 0.506
R21306 vss.n10455 vss.n10454 0.505
R21307 vss.n15212 vss.n15211 0.504
R21308 vss.n10454 vss.n10453 0.495
R21309 vss.n15120 vss.n15108 0.494
R21310 vss.n9153 vss.n9126 0.473
R21311 vss.n10420 vss.n10390 0.472
R21312 vss.n9064 vss.n9033 0.471
R21313 vss.n9095 vss.n9064 0.471
R21314 vss.n9007 vss.n9005 0.471
R21315 vss.n10390 vss.n10355 0.469
R21316 vss.n15818 vss.n15817 0.468
R21317 vss.n10355 vss.n10320 0.466
R21318 vss.n9029 vss.n9028 0.464
R21319 vss.n10320 vss.n10295 0.463
R21320 vss.n9111 vss.n9110 0.461
R21321 vss.n22006 vss.n22005 0.461
R21322 vss.n21956 vss.n21955 0.461
R21323 vss.n21782 vss.n21693 0.461
R21324 vss.n22062 vss.n22061 0.461
R21325 vss.n3955 vss.n3954 0.461
R21326 vss.n3905 vss.n3904 0.461
R21327 vss.n3731 vss.n3642 0.461
R21328 vss.n4011 vss.n4010 0.461
R21329 vss.n21929 vss.n21928 0.46
R21330 vss.n3878 vss.n3877 0.46
R21331 vss.n9672 vss.n9669 0.457
R21332 vss.n10454 vss.n10420 0.457
R21333 vss.n9033 vss.n9003 0.457
R21334 vss.n10295 vss.n10276 0.454
R21335 vss.n11836 vss.n11835 0.452
R21336 vss.n13639 vss.n13638 0.452
R21337 vss.n13098 vss.n13097 0.452
R21338 vss.n13015 vss.n13014 0.452
R21339 vss.n10729 vss.n10728 0.452
R21340 vss.n10529 vss.n10528 0.452
R21341 vss.n11834 vss.n11833 0.452
R21342 vss.n10727 vss.n10726 0.452
R21343 vss.n12252 vss.n12251 0.452
R21344 vss.n11928 vss.n11927 0.452
R21345 vss.n14089 vss.n14088 0.452
R21346 vss.n11556 vss.n11555 0.452
R21347 vss.n13939 vss.n13938 0.452
R21348 vss.n14531 vss.n14530 0.452
R21349 vss.n13501 vss.n13500 0.452
R21350 vss.n14972 vss.n14971 0.452
R21351 vss.n9003 vss.n8972 0.452
R21352 vss.n10276 vss.n10251 0.449
R21353 vss.n10420 vss.n10419 0.449
R21354 vss.n17668 vss.n17667 0.444
R21355 vss.n17677 vss.n17669 0.444
R21356 vss.n18935 vss.n18934 0.444
R21357 vss.n18927 vss.n17694 0.444
R21358 vss.n18848 vss.n17772 0.444
R21359 vss.n18843 vss.n17773 0.444
R21360 vss.n18813 vss.n17804 0.444
R21361 vss.n18808 vss.n17806 0.444
R21362 vss.n18729 vss.n17877 0.444
R21363 vss.n18722 vss.n17881 0.444
R21364 vss.n18694 vss.n18693 0.444
R21365 vss.n18686 vss.n17907 0.444
R21366 vss.n18607 vss.n17985 0.444
R21367 vss.n18602 vss.n17986 0.444
R21368 vss.n18572 vss.n18017 0.444
R21369 vss.n18567 vss.n18019 0.444
R21370 vss.n18488 vss.n18090 0.444
R21371 vss.n18481 vss.n18094 0.444
R21372 vss.n18453 vss.n18452 0.444
R21373 vss.n18445 vss.n18120 0.444
R21374 vss.n18366 vss.n18198 0.444
R21375 vss.n18361 vss.n18199 0.444
R21376 vss.n18331 vss.n18230 0.444
R21377 vss.n18326 vss.n18232 0.444
R21378 vss.n20358 vss.n17591 0.444
R21379 vss.n17590 vss.n17588 0.444
R21380 vss.n20241 vss.n19072 0.444
R21381 vss.n20236 vss.n19073 0.444
R21382 vss.n20206 vss.n19104 0.444
R21383 vss.n20201 vss.n19106 0.444
R21384 vss.n19175 vss.n19174 0.444
R21385 vss.n19184 vss.n19176 0.444
R21386 vss.n20081 vss.n20080 0.444
R21387 vss.n20073 vss.n19201 0.444
R21388 vss.n19994 vss.n19279 0.444
R21389 vss.n19989 vss.n19280 0.444
R21390 vss.n19959 vss.n19311 0.444
R21391 vss.n19954 vss.n19313 0.444
R21392 vss.n19382 vss.n19381 0.444
R21393 vss.n19391 vss.n19383 0.444
R21394 vss.n19834 vss.n19833 0.444
R21395 vss.n19826 vss.n19408 0.444
R21396 vss.n19747 vss.n19486 0.444
R21397 vss.n19742 vss.n19487 0.444
R21398 vss.n19712 vss.n19518 0.444
R21399 vss.n19707 vss.n19520 0.444
R21400 vss.n19598 vss.n19597 0.444
R21401 vss.n4278 vss.n4277 0.444
R21402 vss.n4287 vss.n4279 0.444
R21403 vss.n5545 vss.n5544 0.444
R21404 vss.n5537 vss.n4304 0.444
R21405 vss.n5458 vss.n4382 0.444
R21406 vss.n5453 vss.n4383 0.444
R21407 vss.n5423 vss.n4414 0.444
R21408 vss.n5418 vss.n4416 0.444
R21409 vss.n5339 vss.n4487 0.444
R21410 vss.n5332 vss.n4491 0.444
R21411 vss.n5304 vss.n5303 0.444
R21412 vss.n5296 vss.n4517 0.444
R21413 vss.n5217 vss.n4595 0.444
R21414 vss.n5212 vss.n4596 0.444
R21415 vss.n5182 vss.n4627 0.444
R21416 vss.n5177 vss.n4629 0.444
R21417 vss.n5098 vss.n4700 0.444
R21418 vss.n5091 vss.n4704 0.444
R21419 vss.n5063 vss.n5062 0.444
R21420 vss.n5055 vss.n4730 0.444
R21421 vss.n4976 vss.n4808 0.444
R21422 vss.n4971 vss.n4809 0.444
R21423 vss.n4941 vss.n4840 0.444
R21424 vss.n4936 vss.n4842 0.444
R21425 vss.n6968 vss.n4201 0.444
R21426 vss.n4200 vss.n4198 0.444
R21427 vss.n6851 vss.n5682 0.444
R21428 vss.n6846 vss.n5683 0.444
R21429 vss.n6816 vss.n5714 0.444
R21430 vss.n6811 vss.n5716 0.444
R21431 vss.n5785 vss.n5784 0.444
R21432 vss.n5794 vss.n5786 0.444
R21433 vss.n6691 vss.n6690 0.444
R21434 vss.n6683 vss.n5811 0.444
R21435 vss.n6604 vss.n5889 0.444
R21436 vss.n6599 vss.n5890 0.444
R21437 vss.n6569 vss.n5921 0.444
R21438 vss.n6564 vss.n5923 0.444
R21439 vss.n5992 vss.n5991 0.444
R21440 vss.n6001 vss.n5993 0.444
R21441 vss.n6444 vss.n6443 0.444
R21442 vss.n6436 vss.n6018 0.444
R21443 vss.n6357 vss.n6096 0.444
R21444 vss.n6352 vss.n6097 0.444
R21445 vss.n6322 vss.n6128 0.444
R21446 vss.n6317 vss.n6130 0.444
R21447 vss.n6208 vss.n6207 0.444
R21448 vss.n9126 vss.n9095 0.443
R21449 vss.n10185 bandgapmd_0.bg_resm_0.vss 0.44
R21450 vss.n20318 vss.n17575 0.433
R21451 vss.n6928 vss.n4185 0.433
R21452 vss.n21936 vss.n21935 0.43
R21453 vss.n22013 vss.n22012 0.43
R21454 vss.n21963 vss.n21962 0.43
R21455 vss.n21778 vss.n21695 0.43
R21456 vss.n22055 vss.n22054 0.43
R21457 vss.n3885 vss.n3884 0.43
R21458 vss.n3962 vss.n3961 0.43
R21459 vss.n3912 vss.n3911 0.43
R21460 vss.n3727 vss.n3644 0.43
R21461 vss.n4004 vss.n4003 0.43
R21462 vss.n22603 vss.n22602 0.426
R21463 vss.n22602 vss.n22595 0.426
R21464 vss.n22583 vss.n22576 0.426
R21465 vss.n22585 vss.n22583 0.426
R21466 vss.n22395 vss.n22394 0.426
R21467 vss.n22394 vss.n22387 0.426
R21468 vss.n22375 vss.n22368 0.426
R21469 vss.n22377 vss.n22375 0.426
R21470 vss.n22187 vss.n22186 0.426
R21471 vss.n22186 vss.n22179 0.426
R21472 vss.n22167 vss.n22160 0.426
R21473 vss.n22169 vss.n22167 0.426
R21474 vss.n21531 vss.n21530 0.426
R21475 vss.n21530 vss.n21523 0.426
R21476 vss.n21511 vss.n21504 0.426
R21477 vss.n21513 vss.n21511 0.426
R21478 vss.n21323 vss.n21322 0.426
R21479 vss.n21322 vss.n21315 0.426
R21480 vss.n21303 vss.n21296 0.426
R21481 vss.n21305 vss.n21303 0.426
R21482 vss.n21115 vss.n21114 0.426
R21483 vss.n21114 vss.n21107 0.426
R21484 vss.n21095 vss.n21088 0.426
R21485 vss.n21097 vss.n21095 0.426
R21486 vss.n20907 vss.n20906 0.426
R21487 vss.n20906 vss.n20899 0.426
R21488 vss.n8766 vss.n8765 0.426
R21489 vss.n8765 vss.n8758 0.426
R21490 vss.n8746 vss.n8739 0.426
R21491 vss.n8748 vss.n8746 0.426
R21492 vss.n8558 vss.n8557 0.426
R21493 vss.n8557 vss.n8550 0.426
R21494 vss.n8538 vss.n8531 0.426
R21495 vss.n8540 vss.n8538 0.426
R21496 vss.n8350 vss.n8349 0.426
R21497 vss.n8349 vss.n8342 0.426
R21498 vss.n8330 vss.n8323 0.426
R21499 vss.n8332 vss.n8330 0.426
R21500 vss.n8142 vss.n8141 0.426
R21501 vss.n8141 vss.n8134 0.426
R21502 vss.n8122 vss.n8115 0.426
R21503 vss.n8124 vss.n8122 0.426
R21504 vss.n7934 vss.n7933 0.426
R21505 vss.n7933 vss.n7926 0.426
R21506 vss.n7914 vss.n7907 0.426
R21507 vss.n7916 vss.n7914 0.426
R21508 vss.n7725 vss.n7724 0.426
R21509 vss.n7724 vss.n7717 0.426
R21510 vss.n7705 vss.n7698 0.426
R21511 vss.n7707 vss.n7705 0.426
R21512 vss.n7517 vss.n7516 0.426
R21513 vss.n7516 vss.n7509 0.426
R21514 vss.n10220 vss.n10219 0.426
R21515 vss.n9038 vss.n9036 0.421
R21516 vss.n17330 vss.t316 0.407
R21517 vss.n9197 vss.n9196 0.4
R21518 vss.n21791 vss.n21790 0.398
R21519 vss.n3740 vss.n3739 0.398
R21520 vss.n11838 vss.n11837 0.395
R21521 vss.n13100 vss.n13099 0.395
R21522 vss.n14080 vss.n14079 0.395
R21523 vss.n13102 vss.n13101 0.395
R21524 vss.n12320 vss.n12319 0.395
R21525 vss.n10540 vss.n10539 0.395
R21526 vss.n10678 vss.n10677 0.395
R21527 vss.n11840 vss.n11839 0.395
R21528 vss.n12250 vss.n12249 0.395
R21529 vss.n11926 vss.n11925 0.395
R21530 vss.n14091 vss.n14090 0.395
R21531 vss.n13937 vss.n13936 0.395
R21532 vss.n11558 vss.n11557 0.395
R21533 vss.n14166 vss.n14165 0.395
R21534 vss.n14688 vss.n14687 0.395
R21535 vss.n14970 vss.n14969 0.395
R21536 vss.n16455 vss.n16454 0.384
R21537 vss.n16502 vss.n16501 0.384
R21538 vss.n16697 vss.n16696 0.384
R21539 vss.n16758 vss.n16757 0.384
R21540 vss.n16799 vss.n16798 0.384
R21541 vss.n16890 vss.n16881 0.384
R21542 vss.n16927 vss.n16926 0.384
R21543 vss.n16988 vss.n16987 0.384
R21544 vss.n17041 vss.n17040 0.384
R21545 vss.n17126 vss.n17117 0.384
R21546 vss.n17163 vss.n17162 0.384
R21547 vss.n17224 vss.n17223 0.384
R21548 vss.n17288 vss.n17287 0.384
R21549 vss.n15935 vss.n15934 0.384
R21550 vss.n15974 vss.n15972 0.384
R21551 vss.n16035 vss.n16034 0.384
R21552 vss.n16079 vss.n16078 0.384
R21553 vss.n16171 vss.n16170 0.384
R21554 vss.n16210 vss.n16208 0.384
R21555 vss.n15241 vss.n15240 0.384
R21556 vss.n15219 vss.n15218 0.384
R21557 vss.n15508 vss.n15507 0.384
R21558 vss.n15555 vss.n15554 0.384
R21559 vss.n15744 vss.n15743 0.384
R21560 vss.n15785 vss.n15784 0.384
R21561 vss.n15872 vss.n15866 0.384
R21562 vss.n15122 vss.n15121 0.382
R21563 vss.n14586 vss.n14578 0.38
R21564 vss.n14409 vss.n14405 0.38
R21565 vss.n14722 vss.n14714 0.38
R21566 vss.n14586 vss.n14579 0.38
R21567 vss.n13307 vss.n13303 0.38
R21568 vss.n14722 vss.n14715 0.38
R21569 vss.n14995 vss.n14987 0.38
R21570 vss.n12950 vss.n12943 0.38
R21571 vss.n13161 vss.n13154 0.38
R21572 vss.n14995 vss.n14994 0.38
R21573 vss.n10538 vss.n10530 0.38
R21574 vss.n13942 vss.n13940 0.38
R21575 vss.n11680 vss.n11678 0.38
R21576 vss.n13942 vss.n13941 0.38
R21577 vss.n11680 vss.n11679 0.38
R21578 vss.n11552 vss.n11545 0.38
R21579 vss.n11521 vss.n11514 0.38
R21580 vss.n12255 vss.n12253 0.38
R21581 vss.n10538 vss.n10531 0.38
R21582 vss.n12991 vss.n12984 0.38
R21583 vss.n12981 vss.n12974 0.38
R21584 vss.n12391 vss.n12384 0.38
R21585 vss.n12364 vss.n12357 0.38
R21586 vss.n10695 vss.n10688 0.38
R21587 vss.n10705 vss.n10698 0.38
R21588 vss.n13418 vss.n13411 0.38
R21589 vss.n13497 vss.n13490 0.38
R21590 vss.n13077 vss.n13070 0.38
R21591 vss.n10630 vss.n10623 0.38
R21592 vss.n10790 vss.n10783 0.38
R21593 vss.n12298 vss.n12291 0.38
R21594 vss.n12255 vss.n12254 0.38
R21595 vss.n11931 vss.n11929 0.38
R21596 vss.n11931 vss.n11930 0.38
R21597 vss.n14162 vss.n14155 0.38
R21598 vss.n14119 vss.n14112 0.38
R21599 vss.n13738 vss.n13731 0.38
R21600 vss.n11435 vss.n11428 0.38
R21601 vss.n11875 vss.n11868 0.38
R21602 vss.n11911 vss.n11904 0.38
R21603 vss.n13785 vss.n13778 0.38
R21604 vss.n13796 vss.n13789 0.38
R21605 vss.n16264 vss.n16256 0.38
R21606 vss.n17527 vss.n17518 0.376
R21607 vss.n17514 vss.n17506 0.376
R21608 vss.n21891 vss.n21890 0.376
R21609 vss.n21900 vss.n21899 0.376
R21610 vss.n21834 vss.n21830 0.376
R21611 vss.n21841 vss.n21837 0.376
R21612 vss.n21725 vss.n21720 0.376
R21613 vss.n21725 vss.n21718 0.376
R21614 vss.n21735 vss.n21716 0.376
R21615 vss.n21736 vss.n21735 0.376
R21616 vss.n21765 vss.n21764 0.376
R21617 vss.n21767 vss.n21761 0.376
R21618 vss.n21682 vss.n21681 0.376
R21619 vss.n21678 vss.n21677 0.376
R21620 vss.n21667 vss.n21659 0.376
R21621 vss.n12055 vss.n12048 0.376
R21622 vss.n12045 vss.n12038 0.376
R21623 vss.n10974 vss.n10967 0.376
R21624 vss.n10984 vss.n10977 0.376
R21625 vss.n13837 vss.n13830 0.376
R21626 vss.n13827 vss.n13820 0.376
R21627 vss.n11129 vss.n11122 0.376
R21628 vss.n11119 vss.n11112 0.376
R21629 vss.n13368 vss.n13361 0.376
R21630 vss.n13388 vss.n13381 0.376
R21631 vss.n14200 vss.n14193 0.376
R21632 vss.n14210 vss.n14203 0.376
R21633 vss.n12894 vss.n12893 0.376
R21634 vss.n12893 vss.n12880 0.376
R21635 vss.n12484 vss.n12471 0.376
R21636 vss.n3840 vss.n3839 0.376
R21637 vss.n3849 vss.n3848 0.376
R21638 vss.n3783 vss.n3779 0.376
R21639 vss.n3790 vss.n3786 0.376
R21640 vss.n3674 vss.n3669 0.376
R21641 vss.n3674 vss.n3667 0.376
R21642 vss.n3684 vss.n3665 0.376
R21643 vss.n3685 vss.n3684 0.376
R21644 vss.n3714 vss.n3713 0.376
R21645 vss.n3716 vss.n3710 0.376
R21646 vss.n3631 vss.n3630 0.376
R21647 vss.n3627 vss.n3626 0.376
R21648 vss.n3616 vss.n3608 0.376
R21649 vss.n4137 vss.n4128 0.376
R21650 vss.n4124 vss.n4116 0.376
R21651 vss.n1649 vss.n1640 0.376
R21652 vss.n1637 vss.n1628 0.376
R21653 vss.n1622 vss.n1613 0.376
R21654 vss.n1610 vss.n1601 0.376
R21655 vss.n1597 vss.n1588 0.376
R21656 vss.n1585 vss.n1576 0.376
R21657 vss.n1572 vss.n1563 0.376
R21658 vss.n1559 vss.n1550 0.376
R21659 vss.n1542 vss.n1530 0.376
R21660 vss.n1527 vss.n1518 0.376
R21661 vss.n1514 vss.n1505 0.376
R21662 vss.n1502 vss.n1493 0.376
R21663 vss.n1487 vss.n1478 0.376
R21664 vss.n1475 vss.n1466 0.376
R21665 vss.n110 vss.n101 0.376
R21666 vss.n98 vss.n89 0.376
R21667 vss.n83 vss.n74 0.376
R21668 vss.n71 vss.n62 0.376
R21669 vss.n58 vss.n49 0.376
R21670 vss.n46 vss.n37 0.376
R21671 vss.n33 vss.n24 0.376
R21672 vss.n20 vss.n11 0.376
R21673 vss.n1322 vss.n1313 0.376
R21674 vss.n1334 vss.n1325 0.376
R21675 vss.n1348 vss.n1339 0.376
R21676 vss.n1360 vss.n1351 0.376
R21677 vss.n1375 vss.n1366 0.376
R21678 vss.n1387 vss.n1378 0.376
R21679 vss.n14003 vss.n14002 0.366
R21680 vss.n11595 vss.n11594 0.366
R21681 vss.n10480 vss.n10479 0.366
R21682 vss.n10848 vss.n10847 0.366
R21683 vss.n10892 vss.n10891 0.366
R21684 vss.n14643 vss.n14641 0.366
R21685 vss.n13564 vss.n13563 0.366
R21686 vss.n21861 vss.n21860 0.362
R21687 vss.n21817 vss.n21815 0.362
R21688 vss.n3810 vss.n3809 0.362
R21689 vss.n3766 vss.n3764 0.362
R21690 vss.n19027 vss.n17629 0.355
R21691 vss.n19001 vss.n17642 0.355
R21692 vss.n17648 vss.n17642 0.355
R21693 vss.n18899 vss.n17723 0.355
R21694 vss.n18899 vss.n18898 0.355
R21695 vss.n18877 vss.n17743 0.355
R21696 vss.n18877 vss.n17744 0.355
R21697 vss.n18779 vss.n17830 0.355
R21698 vss.n18779 vss.n17831 0.355
R21699 vss.n18758 vss.n18757 0.355
R21700 vss.n18757 vss.n17854 0.355
R21701 vss.n18658 vss.n17936 0.355
R21702 vss.n18658 vss.n18657 0.355
R21703 vss.n18636 vss.n17956 0.355
R21704 vss.n18636 vss.n17957 0.355
R21705 vss.n18538 vss.n18043 0.355
R21706 vss.n18538 vss.n18044 0.355
R21707 vss.n18517 vss.n18516 0.355
R21708 vss.n18516 vss.n18067 0.355
R21709 vss.n18417 vss.n18149 0.355
R21710 vss.n18417 vss.n18416 0.355
R21711 vss.n18395 vss.n18169 0.355
R21712 vss.n18395 vss.n18170 0.355
R21713 vss.n18297 vss.n18256 0.355
R21714 vss.n18297 vss.n18257 0.355
R21715 vss.n19030 vss.n17624 0.355
R21716 vss.n17621 vss.n17618 0.355
R21717 vss.n20271 vss.n20270 0.355
R21718 vss.n20270 vss.n19043 0.355
R21719 vss.n20172 vss.n19130 0.355
R21720 vss.n20172 vss.n19131 0.355
R21721 vss.n20147 vss.n19149 0.355
R21722 vss.n19155 vss.n19149 0.355
R21723 vss.n20045 vss.n19230 0.355
R21724 vss.n20045 vss.n20044 0.355
R21725 vss.n20023 vss.n19250 0.355
R21726 vss.n20023 vss.n19251 0.355
R21727 vss.n19925 vss.n19337 0.355
R21728 vss.n19925 vss.n19338 0.355
R21729 vss.n19900 vss.n19356 0.355
R21730 vss.n19362 vss.n19356 0.355
R21731 vss.n19798 vss.n19437 0.355
R21732 vss.n19798 vss.n19797 0.355
R21733 vss.n19776 vss.n19457 0.355
R21734 vss.n19776 vss.n19458 0.355
R21735 vss.n19678 vss.n19544 0.355
R21736 vss.n19678 vss.n19545 0.355
R21737 vss.n19653 vss.n19563 0.355
R21738 vss.n19569 vss.n19563 0.355
R21739 vss.n13699 vss.n13693 0.355
R21740 vss.n14350 vss.n14344 0.355
R21741 vss.n14483 vss.n14478 0.355
R21742 vss.n11774 vss.n11770 0.355
R21743 vss.n11351 vss.n11346 0.355
R21744 vss.n10760 vss.n10754 0.355
R21745 vss.n10748 vss.n10743 0.355
R21746 vss.n12436 vss.n12432 0.355
R21747 vss.n12797 vss.n12791 0.355
R21748 vss.n13219 vss.n13214 0.355
R21749 vss.n13572 vss.n13568 0.355
R21750 vss.n14653 vss.n14648 0.355
R21751 vss.n13330 vss.n13325 0.355
R21752 vss.n11359 vss.n11355 0.355
R21753 vss.n13046 vss.n13040 0.355
R21754 vss.n13711 vss.n13705 0.355
R21755 vss.n13034 vss.n13029 0.355
R21756 vss.n14037 vss.n14032 0.355
R21757 vss.n5637 vss.n4239 0.355
R21758 vss.n5611 vss.n4252 0.355
R21759 vss.n4258 vss.n4252 0.355
R21760 vss.n5509 vss.n4333 0.355
R21761 vss.n5509 vss.n5508 0.355
R21762 vss.n5487 vss.n4353 0.355
R21763 vss.n5487 vss.n4354 0.355
R21764 vss.n5389 vss.n4440 0.355
R21765 vss.n5389 vss.n4441 0.355
R21766 vss.n5368 vss.n5367 0.355
R21767 vss.n5367 vss.n4464 0.355
R21768 vss.n5268 vss.n4546 0.355
R21769 vss.n5268 vss.n5267 0.355
R21770 vss.n5246 vss.n4566 0.355
R21771 vss.n5246 vss.n4567 0.355
R21772 vss.n5148 vss.n4653 0.355
R21773 vss.n5148 vss.n4654 0.355
R21774 vss.n5127 vss.n5126 0.355
R21775 vss.n5126 vss.n4677 0.355
R21776 vss.n5027 vss.n4759 0.355
R21777 vss.n5027 vss.n5026 0.355
R21778 vss.n5005 vss.n4779 0.355
R21779 vss.n5005 vss.n4780 0.355
R21780 vss.n4907 vss.n4866 0.355
R21781 vss.n4907 vss.n4867 0.355
R21782 vss.n5640 vss.n4234 0.355
R21783 vss.n4231 vss.n4228 0.355
R21784 vss.n6881 vss.n6880 0.355
R21785 vss.n6880 vss.n5653 0.355
R21786 vss.n6782 vss.n5740 0.355
R21787 vss.n6782 vss.n5741 0.355
R21788 vss.n6757 vss.n5759 0.355
R21789 vss.n5765 vss.n5759 0.355
R21790 vss.n6655 vss.n5840 0.355
R21791 vss.n6655 vss.n6654 0.355
R21792 vss.n6633 vss.n5860 0.355
R21793 vss.n6633 vss.n5861 0.355
R21794 vss.n6535 vss.n5947 0.355
R21795 vss.n6535 vss.n5948 0.355
R21796 vss.n6510 vss.n5966 0.355
R21797 vss.n5972 vss.n5966 0.355
R21798 vss.n6408 vss.n6047 0.355
R21799 vss.n6408 vss.n6407 0.355
R21800 vss.n6386 vss.n6067 0.355
R21801 vss.n6386 vss.n6068 0.355
R21802 vss.n6288 vss.n6154 0.355
R21803 vss.n6288 vss.n6155 0.355
R21804 vss.n6263 vss.n6173 0.355
R21805 vss.n6179 vss.n6173 0.355
R21806 vss.n15210 vss.n15209 0.355
R21807 vss.n9682 vss.t231 0.349
R21808 vss.n9115 vss.n9114 0.349
R21809 vss.n11353 vss.n11351 0.343
R21810 vss.n12798 vss.n12797 0.343
R21811 vss.n13220 vss.n13219 0.343
R21812 vss.n11362 vss.n11359 0.343
R21813 vss.n13712 vss.n13711 0.343
R21814 vss.n10761 vss.n10760 0.343
R21815 vss.n13047 vss.n13046 0.343
R21816 vss.n10751 vss.n10748 0.343
R21817 vss.n13037 vss.n13034 0.343
R21818 vss.n13701 vss.n13699 0.343
R21819 vss.n10233 vss.n10232 0.338
R21820 vss.n13469 vss.n13468 0.336
R21821 vss.n12269 vss.n12268 0.336
R21822 vss.n13409 vss.n13408 0.336
R21823 vss.n10781 vss.n10780 0.336
R21824 vss.n9140 vss.n9139 0.335
R21825 vss.n13573 vss.n13572 0.33
R21826 vss.n13331 vss.n13330 0.33
R21827 vss.n10456 vss.n10455 0.309
R21828 vss.n9197 vss.n9193 0.306
R21829 vss.n10278 vss.n10277 0.301
R21830 vss.n14036 vss.n14035 0.295
R21831 vss.n13329 vss.n13328 0.295
R21832 vss.n13218 vss.n13217 0.295
R21833 vss.n9040 vss.n9039 0.289
R21834 vss.n14264 vss.n14263 0.287
R21835 vss.n9071 vss.n9070 0.285
R21836 vss.n22698 vss.n22697 0.284
R21837 vss.n22709 vss.n22708 0.284
R21838 vss.n22689 vss.n22677 0.284
R21839 vss.n22679 vss.n22678 0.284
R21840 vss.n22490 vss.n22489 0.284
R21841 vss.n22501 vss.n22500 0.284
R21842 vss.n22481 vss.n22469 0.284
R21843 vss.n22471 vss.n22470 0.284
R21844 vss.n22282 vss.n22281 0.284
R21845 vss.n22293 vss.n22292 0.284
R21846 vss.n22273 vss.n22261 0.284
R21847 vss.n22263 vss.n22262 0.284
R21848 vss.n22072 vss.n22071 0.284
R21849 vss.n21603 vss.n21591 0.284
R21850 vss.n21593 vss.n21592 0.284
R21851 vss.n21418 vss.n21417 0.284
R21852 vss.n21429 vss.n21428 0.284
R21853 vss.n21409 vss.n21397 0.284
R21854 vss.n21399 vss.n21398 0.284
R21855 vss.n21210 vss.n21209 0.284
R21856 vss.n21221 vss.n21220 0.284
R21857 vss.n21201 vss.n21189 0.284
R21858 vss.n21191 vss.n21190 0.284
R21859 vss.n21002 vss.n21001 0.284
R21860 vss.n21013 vss.n21012 0.284
R21861 vss.n20993 vss.n20981 0.284
R21862 vss.n20983 vss.n20982 0.284
R21863 vss.n8861 vss.n8860 0.284
R21864 vss.n8872 vss.n8871 0.284
R21865 vss.n8852 vss.n8840 0.284
R21866 vss.n8842 vss.n8841 0.284
R21867 vss.n8653 vss.n8652 0.284
R21868 vss.n8664 vss.n8663 0.284
R21869 vss.n8644 vss.n8632 0.284
R21870 vss.n8634 vss.n8633 0.284
R21871 vss.n8445 vss.n8444 0.284
R21872 vss.n8456 vss.n8455 0.284
R21873 vss.n8436 vss.n8424 0.284
R21874 vss.n8426 vss.n8425 0.284
R21875 vss.n8232 vss.n8231 0.284
R21876 vss.n8229 vss.n8217 0.284
R21877 vss.n8219 vss.n8218 0.284
R21878 vss.n8029 vss.n8028 0.284
R21879 vss.n8040 vss.n8039 0.284
R21880 vss.n8020 vss.n8008 0.284
R21881 vss.n8010 vss.n8009 0.284
R21882 vss.n7820 vss.n7819 0.284
R21883 vss.n7831 vss.n7830 0.284
R21884 vss.n7811 vss.n7799 0.284
R21885 vss.n7801 vss.n7800 0.284
R21886 vss.n7612 vss.n7611 0.284
R21887 vss.n7623 vss.n7622 0.284
R21888 vss.n7603 vss.n7591 0.284
R21889 vss.n7593 vss.n7592 0.284
R21890 vss.n16780 vss.t309 0.283
R21891 vss.n15310 vss.t228 0.283
R21892 vss.n9682 vss.t230 0.277
R21893 vss.n21590 vss.n21589 0.276
R21894 vss.n20308 vss.n17556 0.27
R21895 vss.n6918 vss.n4166 0.27
R21896 vss.n17330 vss.n17329 0.269
R21897 vss.n9119 vss.n9118 0.266
R21898 vss.n18964 vss.n17675 0.266
R21899 vss.n18959 vss.n17676 0.266
R21900 vss.n18940 vss.n18939 0.266
R21901 vss.n17698 vss.n17693 0.266
R21902 vss.n18842 vss.n17777 0.266
R21903 vss.n18835 vss.n17781 0.266
R21904 vss.n18822 vss.n18821 0.266
R21905 vss.n18814 vss.n17797 0.266
R21906 vss.n17884 vss.n17883 0.266
R21907 vss.n17893 vss.n17885 0.266
R21908 vss.n18699 vss.n18698 0.266
R21909 vss.n17911 vss.n17906 0.266
R21910 vss.n18601 vss.n17990 0.266
R21911 vss.n18594 vss.n17994 0.266
R21912 vss.n18581 vss.n18580 0.266
R21913 vss.n18573 vss.n18010 0.266
R21914 vss.n18097 vss.n18096 0.266
R21915 vss.n18106 vss.n18098 0.266
R21916 vss.n18458 vss.n18457 0.266
R21917 vss.n18124 vss.n18119 0.266
R21918 vss.n18360 vss.n18203 0.266
R21919 vss.n18353 vss.n18207 0.266
R21920 vss.n18340 vss.n18339 0.266
R21921 vss.n18332 vss.n18223 0.266
R21922 vss.n20369 vss.n20368 0.266
R21923 vss.n20235 vss.n19077 0.266
R21924 vss.n20228 vss.n19081 0.266
R21925 vss.n20215 vss.n20214 0.266
R21926 vss.n20207 vss.n19097 0.266
R21927 vss.n20110 vss.n19182 0.266
R21928 vss.n20105 vss.n19183 0.266
R21929 vss.n20086 vss.n20085 0.266
R21930 vss.n19205 vss.n19200 0.266
R21931 vss.n19988 vss.n19284 0.266
R21932 vss.n19981 vss.n19288 0.266
R21933 vss.n19968 vss.n19967 0.266
R21934 vss.n19960 vss.n19304 0.266
R21935 vss.n19863 vss.n19389 0.266
R21936 vss.n19858 vss.n19390 0.266
R21937 vss.n19839 vss.n19838 0.266
R21938 vss.n19412 vss.n19407 0.266
R21939 vss.n19741 vss.n19491 0.266
R21940 vss.n19734 vss.n19495 0.266
R21941 vss.n19721 vss.n19720 0.266
R21942 vss.n19713 vss.n19511 0.266
R21943 vss.n19620 vss.n19590 0.266
R21944 vss.n19605 vss.n19591 0.266
R21945 vss.n5574 vss.n4285 0.266
R21946 vss.n5569 vss.n4286 0.266
R21947 vss.n5550 vss.n5549 0.266
R21948 vss.n4308 vss.n4303 0.266
R21949 vss.n5452 vss.n4387 0.266
R21950 vss.n5445 vss.n4391 0.266
R21951 vss.n5432 vss.n5431 0.266
R21952 vss.n5424 vss.n4407 0.266
R21953 vss.n4494 vss.n4493 0.266
R21954 vss.n4503 vss.n4495 0.266
R21955 vss.n5309 vss.n5308 0.266
R21956 vss.n4521 vss.n4516 0.266
R21957 vss.n5211 vss.n4600 0.266
R21958 vss.n5204 vss.n4604 0.266
R21959 vss.n5191 vss.n5190 0.266
R21960 vss.n5183 vss.n4620 0.266
R21961 vss.n4707 vss.n4706 0.266
R21962 vss.n4716 vss.n4708 0.266
R21963 vss.n5068 vss.n5067 0.266
R21964 vss.n4734 vss.n4729 0.266
R21965 vss.n4970 vss.n4813 0.266
R21966 vss.n4963 vss.n4817 0.266
R21967 vss.n4950 vss.n4949 0.266
R21968 vss.n4942 vss.n4833 0.266
R21969 vss.n6979 vss.n6978 0.266
R21970 vss.n6845 vss.n5687 0.266
R21971 vss.n6838 vss.n5691 0.266
R21972 vss.n6825 vss.n6824 0.266
R21973 vss.n6817 vss.n5707 0.266
R21974 vss.n6720 vss.n5792 0.266
R21975 vss.n6715 vss.n5793 0.266
R21976 vss.n6696 vss.n6695 0.266
R21977 vss.n5815 vss.n5810 0.266
R21978 vss.n6598 vss.n5894 0.266
R21979 vss.n6591 vss.n5898 0.266
R21980 vss.n6578 vss.n6577 0.266
R21981 vss.n6570 vss.n5914 0.266
R21982 vss.n6473 vss.n5999 0.266
R21983 vss.n6468 vss.n6000 0.266
R21984 vss.n6449 vss.n6448 0.266
R21985 vss.n6022 vss.n6017 0.266
R21986 vss.n6351 vss.n6101 0.266
R21987 vss.n6344 vss.n6105 0.266
R21988 vss.n6331 vss.n6330 0.266
R21989 vss.n6323 vss.n6121 0.266
R21990 vss.n6230 vss.n6200 0.266
R21991 vss.n6215 vss.n6201 0.266
R21992 vss.n10346 vss.n10344 0.264
R21993 vss.n14351 vss.n14350 0.26
R21994 vss.n14485 vss.n14483 0.26
R21995 vss.n12437 vss.n12436 0.26
R21996 vss.n14655 vss.n14653 0.26
R21997 vss.n12437 vss.n12430 0.26
R21998 vss.n14351 vss.n14342 0.26
R21999 vss.n14655 vss.n14654 0.26
R22000 vss.n14485 vss.n14484 0.26
R22001 vss.n16357 vss.n16350 0.256
R22002 vss.n16378 vss.n16371 0.256
R22003 vss.n16593 vss.n16586 0.256
R22004 vss.n16614 vss.n16607 0.256
R22005 vss.n16683 vss.n16675 0.256
R22006 vss.n16890 vss.n16889 0.256
R22007 vss.n16913 vss.n16904 0.256
R22008 vss.n17010 vss.n17009 0.256
R22009 vss.n17033 vss.n17032 0.256
R22010 vss.n17126 vss.n17125 0.256
R22011 vss.n17149 vss.n17140 0.256
R22012 vss.n17246 vss.n17245 0.256
R22013 vss.n15934 vss.n15927 0.256
R22014 vss.n15958 vss.n15951 0.256
R22015 vss.n16058 vss.n16057 0.256
R22016 vss.n16087 vss.n16077 0.256
R22017 vss.n16170 vss.n16163 0.256
R22018 vss.n16194 vss.n16187 0.256
R22019 vss.n15410 vss.n15403 0.256
R22020 vss.n15431 vss.n15424 0.256
R22021 vss.n15646 vss.n15639 0.256
R22022 vss.n15667 vss.n15660 0.256
R22023 vss.n15873 vss.n15872 0.256
R22024 vss.n10259 vss.n10257 0.254
R22025 vss.n14170 vss.n14167 0.253
R22026 vss.n14391 vss.n14386 0.253
R22027 vss.n13505 vss.n13502 0.253
R22028 vss.n13596 vss.n13593 0.253
R22029 vss.n13289 vss.n13284 0.253
R22030 vss.n13357 vss.n13354 0.253
R22031 vss.n13229 vss.n13222 0.253
R22032 vss.n13188 vss.n13184 0.253
R22033 vss.n14985 vss.n14978 0.253
R22034 vss.n13147 vss.n13140 0.253
R22035 vss.n12828 vss.n12825 0.253
R22036 vss.n10526 vss.n10522 0.253
R22037 vss.n14278 vss.n14271 0.253
R22038 vss.n13843 vss.n13839 0.253
R22039 vss.n11703 vss.n11700 0.253
R22040 vss.n11043 vss.n11036 0.253
R22041 vss.n13969 vss.n13965 0.253
R22042 vss.n11564 vss.n11561 0.253
R22043 vss.n11480 vss.n11473 0.253
R22044 vss.n11698 vss.n11691 0.253
R22045 vss.n12568 vss.n12563 0.253
R22046 vss.n12061 vss.n12057 0.253
R22047 vss.n12417 vss.n12414 0.253
R22048 vss.n12529 vss.n12522 0.253
R22049 vss.n13120 vss.n13113 0.253
R22050 vss.n13669 vss.n13662 0.253
R22051 vss.n12412 vss.n12405 0.253
R22052 vss.n10675 vss.n10668 0.253
R22053 vss.n12329 vss.n12322 0.253
R22054 vss.n11490 vss.n11483 0.253
R22055 vss.n13378 vss.n13371 0.253
R22056 vss.n13461 vss.n13454 0.253
R22057 vss.n13092 vss.n13085 0.253
R22058 vss.n10645 vss.n10638 0.253
R22059 vss.n12314 vss.n12307 0.253
R22060 vss.n10811 vss.n10804 0.253
R22061 vss.n10816 vss.n10813 0.253
R22062 vss.n10923 vss.n10919 0.253
R22063 vss.n10941 vss.n10938 0.253
R22064 vss.n11032 vss.n11028 0.253
R22065 vss.n14566 vss.n14559 0.253
R22066 vss.n14103 vss.n14096 0.253
R22067 vss.n13753 vss.n13746 0.253
R22068 vss.n11450 vss.n11443 0.253
R22069 vss.n11859 vss.n11852 0.253
R22070 vss.n10936 vss.n10929 0.253
R22071 vss.n13656 vss.n13649 0.253
R22072 vss.n14065 vss.n14058 0.253
R22073 vss.n16264 vss.n16258 0.253
R22074 vss.n9176 vss.n9174 0.248
R22075 vss.n12485 vss.n12484 0.247
R22076 vss.n20413 ldomc_0.otaldom_0.nmosbn2m_0.vss 0.247
R22077 vss.n7023 bandgapmd_0.otam_1.nmosbn2m_0.vss 0.247
R22078 vss.n13982 vss.n13981 0.247
R22079 vss.n12085 vss.n12082 0.247
R22080 vss.n10510 vss.n10509 0.247
R22081 vss.n10829 vss.n10827 0.247
R22082 vss.n10903 vss.n10901 0.247
R22083 vss.n10955 vss.n10954 0.247
R22084 vss.n11017 vss.n11014 0.247
R22085 vss.n14363 vss.n14360 0.247
R22086 vss.n13867 vss.n13866 0.247
R22087 vss.n11577 vss.n11576 0.247
R22088 vss.n11766 vss.n11763 0.247
R22089 vss.n13343 vss.n13342 0.247
R22090 vss.n14666 vss.n14664 0.247
R22091 vss.n13584 vss.n13583 0.247
R22092 vss.n14497 vss.n14494 0.247
R22093 vss.n20332 vss.n20331 0.241
R22094 vss.n6942 vss.n6941 0.241
R22095 vss.n22069 vss.n21606 0.24
R22096 vss.n13615 vss.n13613 0.232
R22097 vss.n13429 vss.n13427 0.232
R22098 vss.n10499 vss.n10497 0.232
R22099 vss.n13200 vss.n13198 0.232
R22100 vss.n13926 vss.n13925 0.231
R22101 vss.n12520 vss.n12519 0.231
R22102 vss.n13625 vss.n13623 0.231
R22103 vss.n13438 vss.n13436 0.231
R22104 vss.n11404 vss.n11403 0.231
R22105 vss.n10591 vss.n10590 0.231
R22106 vss.n10599 vss.n10598 0.231
R22107 vss.n11396 vss.n11395 0.231
R22108 vss.n11652 vss.n11651 0.231
R22109 vss.n20374 vss.n20373 0.224
R22110 vss.n6984 vss.n6983 0.224
R22111 vss.n10837 vss.n10836 0.223
R22112 vss.n12239 vss.n12237 0.223
R22113 vss.n10918 vss.n10916 0.223
R22114 vss.n11273 vss.n11271 0.222
R22115 vss.n11026 vss.n11024 0.222
R22116 vss.n21976 vss.n21975 0.212
R22117 vss.n3925 vss.n3924 0.212
R22118 vss.n9177 bandgapmd_0.bg_stupm_0.vss 0.204
R22119 vss.n8921 vss.t306 0.196
R22120 vss.n22039 vss.n22037 0.19
R22121 vss.n21842 vss.n21835 0.19
R22122 vss.n22022 vss.n22020 0.19
R22123 vss.n21680 vss.n21679 0.19
R22124 vss.n21724 vss.n21717 0.19
R22125 vss.n21768 vss.n21766 0.19
R22126 vss.n13105 vss.n13103 0.19
R22127 vss.n11843 vss.n11841 0.19
R22128 vss.n13105 vss.n13104 0.19
R22129 vss.n14083 vss.n14081 0.19
R22130 vss.n10681 vss.n10679 0.19
R22131 vss.n10681 vss.n10680 0.19
R22132 vss.n11843 vss.n11842 0.19
R22133 vss.n14083 vss.n14082 0.19
R22134 vss.n3988 vss.n3986 0.19
R22135 vss.n3791 vss.n3784 0.19
R22136 vss.n3971 vss.n3969 0.19
R22137 vss.n3629 vss.n3628 0.19
R22138 vss.n3673 vss.n3666 0.19
R22139 vss.n3717 vss.n3715 0.19
R22140 vss.n15121 vss.n15097 0.189
R22141 vss.n13164 vss.n13161 0.187
R22142 vss.n12951 vss.n12950 0.187
R22143 vss.n13164 vss.n13163 0.187
R22144 vss.n11553 vss.n11543 0.187
R22145 vss.n11522 vss.n11521 0.187
R22146 vss.n12982 vss.n12981 0.187
R22147 vss.n12992 vss.n12991 0.187
R22148 vss.n12392 vss.n12391 0.187
R22149 vss.n12365 vss.n12364 0.187
R22150 vss.n10696 vss.n10695 0.187
R22151 vss.n10706 vss.n10705 0.187
R22152 vss.n13498 vss.n13497 0.187
R22153 vss.n12299 vss.n12298 0.187
R22154 vss.n13419 vss.n13418 0.187
R22155 vss.n10791 vss.n10790 0.187
R22156 vss.n13797 vss.n13796 0.187
R22157 vss.n13786 vss.n13785 0.187
R22158 vss.n11553 vss.n11552 0.187
R22159 vss.n9171 vss.n9170 0.187
R22160 vss.n13331 vss.n13323 0.185
R22161 vss.n13573 vss.n13566 0.185
R22162 vss.n17528 vss.n17527 0.185
R22163 vss.n17515 vss.n17514 0.185
R22164 vss.n10975 vss.n10974 0.185
R22165 vss.n12056 vss.n12055 0.185
R22166 vss.n12046 vss.n12045 0.185
R22167 vss.n10985 vss.n10984 0.185
R22168 vss.n13828 vss.n13827 0.185
R22169 vss.n11120 vss.n11119 0.185
R22170 vss.n11130 vss.n11129 0.185
R22171 vss.n13838 vss.n13837 0.185
R22172 vss.n14211 vss.n14210 0.185
R22173 vss.n14201 vss.n14200 0.185
R22174 vss.n13389 vss.n13388 0.185
R22175 vss.n13369 vss.n13368 0.185
R22176 vss.n4138 vss.n4137 0.185
R22177 vss.n4125 vss.n4124 0.185
R22178 vss.n1650 vss.n1649 0.185
R22179 vss.n1611 vss.n1610 0.185
R22180 vss.n1598 vss.n1597 0.185
R22181 vss.n1560 vss.n1559 0.185
R22182 vss.n1543 vss.n1542 0.185
R22183 vss.n1503 vss.n1502 0.185
R22184 vss.n1488 vss.n1487 0.185
R22185 vss.n1638 vss.n1637 0.185
R22186 vss.n1623 vss.n1622 0.185
R22187 vss.n1586 vss.n1585 0.185
R22188 vss.n1573 vss.n1572 0.185
R22189 vss.n1528 vss.n1527 0.185
R22190 vss.n1515 vss.n1514 0.185
R22191 vss.n1476 vss.n1475 0.185
R22192 vss.n111 vss.n110 0.185
R22193 vss.n72 vss.n71 0.185
R22194 vss.n59 vss.n58 0.185
R22195 vss.n21 vss.n20 0.185
R22196 vss.n1323 vss.n1322 0.185
R22197 vss.n1361 vss.n1360 0.185
R22198 vss.n1376 vss.n1375 0.185
R22199 vss.n99 vss.n98 0.185
R22200 vss.n84 vss.n83 0.185
R22201 vss.n47 vss.n46 0.185
R22202 vss.n34 vss.n33 0.185
R22203 vss.n1335 vss.n1334 0.185
R22204 vss.n1349 vss.n1348 0.185
R22205 vss.n1388 vss.n1387 0.185
R22206 vss.n21802 ldomc_0.otaldom_0.ncsm_0.vss 0.182
R22207 vss.n3751 bandgapmd_0.otam_1.ncsm_0.vss 0.182
R22208 vss.n22032 vss.n22031 0.179
R22209 vss.n21792 vss.n21688 0.179
R22210 vss.n8921 vss.t305 0.179
R22211 vss.n3981 vss.n3980 0.179
R22212 vss.n3741 vss.n3637 0.179
R22213 vss.n19021 vss.n17630 0.177
R22214 vss.n19021 vss.n17632 0.177
R22215 vss.n19007 vss.n17636 0.177
R22216 vss.n19007 vss.n17640 0.177
R22217 vss.n18892 vss.n17730 0.177
R22218 vss.n18892 vss.n17731 0.177
R22219 vss.n18883 vss.n18882 0.177
R22220 vss.n18882 vss.n18881 0.177
R22221 vss.n18775 vss.n18774 0.177
R22222 vss.n18774 vss.n17835 0.177
R22223 vss.n18764 vss.n17844 0.177
R22224 vss.n18764 vss.n17845 0.177
R22225 vss.n18651 vss.n17943 0.177
R22226 vss.n18651 vss.n17944 0.177
R22227 vss.n18642 vss.n18641 0.177
R22228 vss.n18641 vss.n18640 0.177
R22229 vss.n18534 vss.n18533 0.177
R22230 vss.n18533 vss.n18048 0.177
R22231 vss.n18523 vss.n18057 0.177
R22232 vss.n18523 vss.n18058 0.177
R22233 vss.n18410 vss.n18156 0.177
R22234 vss.n18410 vss.n18157 0.177
R22235 vss.n18401 vss.n18400 0.177
R22236 vss.n18400 vss.n18399 0.177
R22237 vss.n18293 vss.n18292 0.177
R22238 vss.n18292 vss.n18261 0.177
R22239 vss.n18282 vss.n18270 0.177
R22240 vss.n18282 vss.n18271 0.177
R22241 vss.n20287 vss.n17622 0.177
R22242 vss.n20287 vss.n20286 0.177
R22243 vss.n20278 vss.n19038 0.177
R22244 vss.n19045 vss.n19038 0.177
R22245 vss.n20168 vss.n20167 0.177
R22246 vss.n20167 vss.n19135 0.177
R22247 vss.n20153 vss.n19143 0.177
R22248 vss.n20153 vss.n19147 0.177
R22249 vss.n20038 vss.n19237 0.177
R22250 vss.n20038 vss.n19238 0.177
R22251 vss.n20029 vss.n20028 0.177
R22252 vss.n20028 vss.n20027 0.177
R22253 vss.n19921 vss.n19920 0.177
R22254 vss.n19920 vss.n19342 0.177
R22255 vss.n19906 vss.n19350 0.177
R22256 vss.n19906 vss.n19354 0.177
R22257 vss.n19791 vss.n19444 0.177
R22258 vss.n19791 vss.n19445 0.177
R22259 vss.n19782 vss.n19781 0.177
R22260 vss.n19781 vss.n19780 0.177
R22261 vss.n19674 vss.n19673 0.177
R22262 vss.n19673 vss.n19549 0.177
R22263 vss.n19659 vss.n19557 0.177
R22264 vss.n19659 vss.n19561 0.177
R22265 vss.n21922 vss.n21921 0.177
R22266 vss.n13806 vss.n13801 0.177
R22267 vss.n11423 vss.n11417 0.177
R22268 vss.n14438 vss.n14432 0.177
R22269 vss.n13892 vss.n13886 0.177
R22270 vss.n13766 vss.n13760 0.177
R22271 vss.n14138 vss.n14132 0.177
R22272 vss.n11538 vss.n11533 0.177
R22273 vss.n11109 vss.n11103 0.177
R22274 vss.n10994 vss.n10987 0.177
R22275 vss.n11899 vss.n11893 0.177
R22276 vss.n12378 vss.n12373 0.177
R22277 vss.n11965 vss.n11959 0.177
R22278 vss.n12287 vss.n12286 0.177
R22279 vss.n12279 vss.n12272 0.177
R22280 vss.n10767 vss.n10766 0.177
R22281 vss.n10777 vss.n10772 0.177
R22282 vss.n12094 vss.n12087 0.177
R22283 vss.n12629 vss.n12623 0.177
R22284 vss.n10469 vss.n10462 0.177
R22285 vss.n13180 vss.n13175 0.177
R22286 vss.n14937 vss.n14931 0.177
R22287 vss.n14763 vss.n14757 0.177
R22288 vss.n13553 vss.n13546 0.177
R22289 vss.n14130 vss.n14124 0.177
R22290 vss.n12970 vss.n12965 0.177
R22291 vss.n13486 vss.n13485 0.177
R22292 vss.n13478 vss.n13472 0.177
R22293 vss.n13395 vss.n13394 0.177
R22294 vss.n13405 vss.n13399 0.177
R22295 vss.n12939 vss.n12934 0.177
R22296 vss.n11891 vss.n11885 0.177
R22297 vss.n10719 vss.n10714 0.177
R22298 vss.n10610 vss.n10603 0.177
R22299 vss.n13009 vss.n13004 0.177
R22300 vss.n11415 vss.n11409 0.177
R22301 vss.n10557 vss.n10552 0.177
R22302 vss.n10618 vss.n10612 0.177
R22303 vss.n12342 vss.n12336 0.177
R22304 vss.n11603 vss.n11597 0.177
R22305 vss.n11502 vss.n11497 0.177
R22306 vss.n3871 vss.n3870 0.177
R22307 vss.n5631 vss.n4240 0.177
R22308 vss.n5631 vss.n4242 0.177
R22309 vss.n5617 vss.n4246 0.177
R22310 vss.n5617 vss.n4250 0.177
R22311 vss.n5502 vss.n4340 0.177
R22312 vss.n5502 vss.n4341 0.177
R22313 vss.n5493 vss.n5492 0.177
R22314 vss.n5492 vss.n5491 0.177
R22315 vss.n5385 vss.n5384 0.177
R22316 vss.n5384 vss.n4445 0.177
R22317 vss.n5374 vss.n4454 0.177
R22318 vss.n5374 vss.n4455 0.177
R22319 vss.n5261 vss.n4553 0.177
R22320 vss.n5261 vss.n4554 0.177
R22321 vss.n5252 vss.n5251 0.177
R22322 vss.n5251 vss.n5250 0.177
R22323 vss.n5144 vss.n5143 0.177
R22324 vss.n5143 vss.n4658 0.177
R22325 vss.n5133 vss.n4667 0.177
R22326 vss.n5133 vss.n4668 0.177
R22327 vss.n5020 vss.n4766 0.177
R22328 vss.n5020 vss.n4767 0.177
R22329 vss.n5011 vss.n5010 0.177
R22330 vss.n5010 vss.n5009 0.177
R22331 vss.n4903 vss.n4902 0.177
R22332 vss.n4902 vss.n4871 0.177
R22333 vss.n4892 vss.n4880 0.177
R22334 vss.n4892 vss.n4881 0.177
R22335 vss.n6897 vss.n4232 0.177
R22336 vss.n6897 vss.n6896 0.177
R22337 vss.n6888 vss.n5648 0.177
R22338 vss.n5655 vss.n5648 0.177
R22339 vss.n6778 vss.n6777 0.177
R22340 vss.n6777 vss.n5745 0.177
R22341 vss.n6763 vss.n5753 0.177
R22342 vss.n6763 vss.n5757 0.177
R22343 vss.n6648 vss.n5847 0.177
R22344 vss.n6648 vss.n5848 0.177
R22345 vss.n6639 vss.n6638 0.177
R22346 vss.n6638 vss.n6637 0.177
R22347 vss.n6531 vss.n6530 0.177
R22348 vss.n6530 vss.n5952 0.177
R22349 vss.n6516 vss.n5960 0.177
R22350 vss.n6516 vss.n5964 0.177
R22351 vss.n6401 vss.n6054 0.177
R22352 vss.n6401 vss.n6055 0.177
R22353 vss.n6392 vss.n6391 0.177
R22354 vss.n6391 vss.n6390 0.177
R22355 vss.n6284 vss.n6283 0.177
R22356 vss.n6283 vss.n6159 0.177
R22357 vss.n6269 vss.n6167 0.177
R22358 vss.n6269 vss.n6171 0.177
R22359 vss.n20443 ldomc_0.otaldom_0.vss 0.174
R22360 vss.n7053 bandgapmd_0.otam_1.vss 0.174
R22361 vss.n11353 vss.n11352 0.172
R22362 vss.n13701 vss.n13700 0.172
R22363 vss.n10761 vss.n10752 0.172
R22364 vss.n10751 vss.n10750 0.172
R22365 vss.n13047 vss.n13038 0.172
R22366 vss.n13712 vss.n13703 0.172
R22367 vss.n11362 vss.n11361 0.172
R22368 vss.n13037 vss.n13036 0.172
R22369 vss.n12798 vss.n12789 0.172
R22370 vss.n13220 vss.n13212 0.172
R22371 vss.n21794 vss.n21793 0.169
R22372 vss.n3743 vss.n3742 0.169
R22373 vss.n10261 vss.n10259 0.168
R22374 vss.n21876 vss.n21874 0.165
R22375 vss.n21932 vss.n21930 0.165
R22376 vss.n21959 vss.n21957 0.165
R22377 vss.n3825 vss.n3823 0.165
R22378 vss.n3881 vss.n3879 0.165
R22379 vss.n3908 vss.n3906 0.165
R22380 vss.n3455 vss.n3451 0.165
R22381 vss.n1430 vss.n1426 0.165
R22382 vss.n3444 vss.n3441 0.162
R22383 vss.n1419 vss.n1416 0.162
R22384 vss.n17572 vss.n17558 0.151
R22385 vss.n4182 vss.n4168 0.151
R22386 vss.n13891 vss.n13890 0.15
R22387 vss.n11107 vss.n11106 0.15
R22388 vss.n10776 vss.n10775 0.15
R22389 vss.n14935 vss.n14934 0.15
R22390 vss.n14129 vss.n14128 0.15
R22391 vss.n13476 vss.n13475 0.15
R22392 vss.n13404 vss.n13403 0.15
R22393 vss.n12627 vss.n12626 0.15
R22394 vss.n11897 vss.n11896 0.15
R22395 vss.n11422 vss.n11421 0.15
R22396 vss.n11602 vss.n11601 0.15
R22397 vss.n21939 vss.n21923 0.15
R22398 vss.n9174 vss.n9163 0.15
R22399 vss.n3888 vss.n3872 0.15
R22400 vss.n8230 vss.n4018 0.15
R22401 vss.n10293 vss.n10292 0.147
R22402 vss.n9688 vss.n9687 0.146
R22403 vss.n9689 vss.n9688 0.146
R22404 vss.n9693 vss.n9692 0.146
R22405 vss.n9694 vss.n9693 0.146
R22406 vss.n9695 vss.n9694 0.146
R22407 vss.n9696 vss.n9695 0.146
R22408 vss.n9681 vss.n9680 0.146
R22409 vss.n9680 vss.n9679 0.146
R22410 vss.n9679 vss.n9678 0.146
R22411 vss.n9678 vss.n9677 0.146
R22412 vss.n22789 vss.n22759 0.145
R22413 vss.n21854 vss.n21846 0.144
R22414 vss.n9690 vss.n9689 0.144
R22415 vss.n9714 vss.n9681 0.144
R22416 vss.n3803 vss.n3795 0.144
R22417 vss.n17340 vss.n17333 0.142
R22418 vss.n17351 vss.n17344 0.142
R22419 vss.n17362 vss.n17355 0.142
R22420 vss.n17373 vss.n17366 0.142
R22421 vss.n17384 vss.n17377 0.142
R22422 vss.n17395 vss.n17388 0.142
R22423 vss.n17417 vss.n17410 0.142
R22424 vss.n17428 vss.n17421 0.142
R22425 vss.n17439 vss.n17432 0.142
R22426 vss.n17450 vss.n17443 0.142
R22427 vss.n17461 vss.n17454 0.142
R22428 vss.n17472 vss.n17465 0.142
R22429 vss.n17483 vss.n17476 0.142
R22430 vss.n8988 vss.n8986 0.142
R22431 vss.n3498 vss.n3491 0.142
R22432 vss.n3509 vss.n3502 0.142
R22433 vss.n3520 vss.n3513 0.142
R22434 vss.n3531 vss.n3524 0.142
R22435 vss.n3542 vss.n3535 0.142
R22436 vss.n3553 vss.n3546 0.142
R22437 vss.n4027 vss.n4020 0.142
R22438 vss.n4038 vss.n4031 0.142
R22439 vss.n4049 vss.n4042 0.142
R22440 vss.n4060 vss.n4053 0.142
R22441 vss.n4071 vss.n4064 0.142
R22442 vss.n4082 vss.n4075 0.142
R22443 vss.n4093 vss.n4086 0.142
R22444 vss.n8243 vss.n8242 0.14
R22445 vss.n9687 vss.n9686 0.14
R22446 vss.n21701 vss.n21644 0.139
R22447 vss.n3650 vss.n3593 0.139
R22448 vss.n21809 vss.n21808 0.138
R22449 vss.n3758 vss.n3757 0.138
R22450 vss.n17331 vss.n17330 0.138
R22451 vss.n22046 vss.n22043 0.135
R22452 vss.n21675 vss.n21674 0.135
R22453 vss.n3995 vss.n3992 0.135
R22454 vss.n3624 vss.n3623 0.135
R22455 vss.n21760 vss.n21702 0.133
R22456 vss.n3709 vss.n3651 0.133
R22457 vss.n9080 vss.n9078 0.133
R22458 vss.n9129 vss.n9128 0.133
R22459 vss.n17533 vss.n17531 0.132
R22460 vss.n4143 vss.n4141 0.132
R22461 vss.n17488 vss.n17486 0.131
R22462 vss.n9685 vss.n9684 0.131
R22463 vss.n4098 vss.n4096 0.131
R22464 vss.n21739 vss.n21738 0.13
R22465 vss.n22086 vss.n22069 0.13
R22466 vss.n3688 vss.n3687 0.13
R22467 vss.n20505 vss.n17545 0.129
R22468 vss.n7115 vss.n4155 0.129
R22469 vss.n15819 vss.n15818 0.129
R22470 vss.n8927 vss.n8925 0.129
R22471 vss.n17573 vss.n17558 0.129
R22472 vss.n4183 vss.n4168 0.129
R22473 vss.n20799 vss.n17500 0.128
R22474 vss.n7409 vss.n4110 0.128
R22475 vss.n16469 vss.n16468 0.128
R22476 vss.n16484 vss.n16483 0.128
R22477 vss.n16665 vss.n16664 0.128
R22478 vss.n16673 vss.n16665 0.128
R22479 vss.n16683 vss.n16677 0.128
R22480 vss.n16770 vss.n16769 0.128
R22481 vss.n16786 vss.n16785 0.128
R22482 vss.n16901 vss.n16895 0.128
R22483 vss.n16913 vss.n16912 0.128
R22484 vss.n17002 vss.n17001 0.128
R22485 vss.n17027 vss.n17026 0.128
R22486 vss.n17137 vss.n17131 0.128
R22487 vss.n17149 vss.n17148 0.128
R22488 vss.n17238 vss.n17237 0.128
R22489 vss.n17255 vss.n17254 0.128
R22490 vss.n15946 vss.n15945 0.128
R22491 vss.n15960 vss.n15958 0.128
R22492 vss.n16049 vss.n16048 0.128
R22493 vss.n16063 vss.n16062 0.128
R22494 vss.n16182 vss.n16181 0.128
R22495 vss.n16196 vss.n16194 0.128
R22496 vss.n15229 vss.n15228 0.128
R22497 vss.n15314 vss.n15313 0.128
R22498 vss.n15522 vss.n15521 0.128
R22499 vss.n15537 vss.n15536 0.128
R22500 vss.n15758 vss.n15757 0.128
R22501 vss.n15794 vss.n15793 0.128
R22502 vss.n15004 vss.n14997 0.126
R22503 vss.n13128 vss.n13122 0.126
R22504 vss.n11470 vss.n11464 0.126
R22505 vss.n11815 vss.n11808 0.126
R22506 vss.n13137 vss.n13130 0.126
R22507 vss.n13678 vss.n13671 0.126
R22508 vss.n12402 vss.n12395 0.126
R22509 vss.n10665 vss.n10659 0.126
R22510 vss.n10657 vss.n10650 0.126
R22511 vss.n11462 vss.n11455 0.126
R22512 vss.n14712 vss.n14705 0.126
R22513 vss.n13449 vss.n13442 0.126
R22514 vss.n13024 vss.n13017 0.126
R22515 vss.n10581 vss.n10574 0.126
R22516 vss.n10738 vss.n10731 0.126
R22517 vss.n12034 vss.n12027 0.126
R22518 vss.n14576 vss.n14569 0.126
R22519 vss.n13636 vss.n13629 0.126
R22520 vss.n13688 vss.n13681 0.126
R22521 vss.n11385 vss.n11378 0.126
R22522 vss.n11371 vss.n11364 0.126
R22523 vss.n11314 vss.n11307 0.126
R22524 vss.n13646 vss.n13640 0.126
R22525 vss.n13962 vss.n13955 0.126
R22526 vss.n16251 vss.n16242 0.126
R22527 vss.n12239 vss.n12238 0.126
R22528 vss.n10918 vss.n10917 0.126
R22529 vss.n10837 vss.n10830 0.126
R22530 vss.n13597 vss.n13596 0.125
R22531 vss.n13148 vss.n13147 0.125
R22532 vss.n10527 vss.n10526 0.125
R22533 vss.n11565 vss.n11564 0.125
R22534 vss.n12532 vss.n12529 0.125
R22535 vss.n12063 vss.n12061 0.125
R22536 vss.n11481 vss.n11480 0.125
R22537 vss.n13670 vss.n13669 0.125
R22538 vss.n13121 vss.n13120 0.125
R22539 vss.n12419 vss.n12417 0.125
R22540 vss.n12413 vss.n12412 0.125
R22541 vss.n10676 vss.n10675 0.125
R22542 vss.n11491 vss.n11490 0.125
R22543 vss.n12330 vss.n12329 0.125
R22544 vss.n10812 vss.n10811 0.125
R22545 vss.n10818 vss.n10816 0.125
R22546 vss.n10925 vss.n10923 0.125
R22547 vss.n10943 vss.n10941 0.125
R22548 vss.n11034 vss.n11032 0.125
R22549 vss.n10937 vss.n10936 0.125
R22550 vss.n13657 vss.n13656 0.125
R22551 vss.n14066 vss.n14065 0.125
R22552 vss.n11699 vss.n11698 0.125
R22553 vss.n14280 vss.n14278 0.125
R22554 vss.n13845 vss.n13843 0.125
R22555 vss.n13971 vss.n13969 0.125
R22556 vss.n11705 vss.n11703 0.125
R22557 vss.n13359 vss.n13357 0.125
R22558 vss.n13379 vss.n13378 0.125
R22559 vss.n13507 vss.n13505 0.125
R22560 vss.n14567 vss.n14566 0.125
R22561 vss.n14172 vss.n14170 0.125
R22562 vss.n13232 vss.n13229 0.125
R22563 vss.n13191 vss.n13188 0.125
R22564 vss.n12831 vss.n12828 0.125
R22565 vss.n14986 vss.n14985 0.125
R22566 vss.n11026 vss.n11025 0.125
R22567 vss.n11273 vss.n11272 0.125
R22568 vss.n21770 vss.n21760 0.125
R22569 vss.n21911 vss.n21910 0.125
R22570 vss.n9099 vss.n9098 0.125
R22571 vss.n3719 vss.n3709 0.125
R22572 vss.n3860 vss.n3859 0.125
R22573 vss.n21654 vss.n21649 0.125
R22574 vss.n3603 vss.n3598 0.125
R22575 vss.n21949 vss.n21948 0.124
R22576 vss.n3898 vss.n3897 0.124
R22577 vss.n10376 vss.n10375 0.122
R22578 vss.n21757 vss.n21753 0.122
R22579 vss.n3706 vss.n3702 0.122
R22580 vss.n10380 vss.n10378 0.121
R22581 vss.n22000 vss.n21998 0.121
R22582 vss.n3949 vss.n3947 0.121
R22583 vss.n12572 vss.n12571 0.119
R22584 vss.n11167 vss.n11166 0.119
R22585 vss.n21752 vss.n21706 0.118
R22586 vss.n21760 vss.n21699 0.118
R22587 vss.n9690 vss.n9682 0.118
R22588 vss.n3701 vss.n3655 0.118
R22589 vss.n3709 vss.n3648 0.118
R22590 vss.n11337 vss.n11335 0.118
R22591 vss.n12447 vss.n12445 0.118
R22592 vss.n11712 vss.n11710 0.118
R22593 vss.n14289 vss.n14287 0.118
R22594 vss.n12788 vss.n12786 0.118
R22595 vss.n13211 vss.n13209 0.118
R22596 vss.n13605 vss.n13604 0.117
R22597 vss.n14150 vss.n14148 0.117
R22598 vss.n11344 vss.n11342 0.117
R22599 vss.n13724 vss.n13723 0.117
R22600 vss.n13063 vss.n13062 0.117
R22601 vss.n13053 vss.n13051 0.117
R22602 vss.n13718 vss.n13716 0.117
R22603 vss.n14024 vss.n14023 0.117
R22604 vss.n9049 vss.n9047 0.117
R22605 vss.n13615 vss.n13614 0.116
R22606 vss.n13429 vss.n13428 0.116
R22607 vss.n10499 vss.n10498 0.116
R22608 vss.n13200 vss.n13199 0.116
R22609 vss.n11396 vss.n11387 0.116
R22610 vss.n12520 vss.n12511 0.116
R22611 vss.n10591 vss.n10583 0.116
R22612 vss.n11404 vss.n11397 0.116
R22613 vss.n13625 vss.n13624 0.116
R22614 vss.n13438 vss.n13437 0.116
R22615 vss.n10599 vss.n10592 0.116
R22616 vss.n13926 vss.n13918 0.116
R22617 vss.n11652 vss.n11644 0.116
R22618 vss.n20373 vss.n17579 0.115
R22619 vss.n6983 vss.n4189 0.115
R22620 bandgapmd_0.bg_stupm_0.vss vss.n9176 0.112
R22621 vss.n9018 vss.n9016 0.111
R22622 vss.n9067 vss.n9066 0.11
R22623 vss.n20373 vss.n20372 0.11
R22624 vss.n6983 vss.n6982 0.11
R22625 vss.n3431 vss.n3429 0.109
R22626 vss.n1406 vss.n1404 0.109
R22627 vss.n9147 vss.n9146 0.107
R22628 vss.n20397 vss.n17553 0.106
R22629 vss.n21760 vss.n21697 0.106
R22630 vss.n3709 vss.n3646 0.106
R22631 vss.n7007 vss.n4163 0.106
R22632 bandgapmd_0.bg_trimmup_0.vss vss.n9691 0.103
R22633 vss.n15125 vss.n15124 0.103
R22634 vss.n10352 vss.n10338 0.101
R22635 vss.n21774 vss.n21773 0.098
R22636 vss.n3723 vss.n3722 0.098
R22637 vss.n9192 vss.n9163 0.098
R22638 vss.n10338 vss.n10336 0.096
R22639 vss.n17561 vss.n17558 0.096
R22640 vss.n20315 vss.n17608 0.096
R22641 vss.n20315 vss.n17609 0.096
R22642 vss.n10249 vss.n10248 0.096
R22643 vss.n4171 vss.n4168 0.096
R22644 vss.n6925 vss.n4218 0.096
R22645 vss.n6925 vss.n4219 0.096
R22646 vss.n10412 vss.n10411 0.096
R22647 vss.n10408 vss.n10407 0.095
R22648 vss.n17419 vss.n17417 0.095
R22649 vss.n17430 vss.n17428 0.095
R22650 vss.n17441 vss.n17439 0.095
R22651 vss.n17452 vss.n17450 0.095
R22652 vss.n17463 vss.n17461 0.095
R22653 vss.n17474 vss.n17472 0.095
R22654 vss.n17485 vss.n17483 0.095
R22655 vss.n3500 vss.n3498 0.095
R22656 vss.n3511 vss.n3509 0.095
R22657 vss.n3522 vss.n3520 0.095
R22658 vss.n3533 vss.n3531 0.095
R22659 vss.n3544 vss.n3542 0.095
R22660 vss.n3555 vss.n3553 0.095
R22661 vss.n4029 vss.n4027 0.095
R22662 vss.n4040 vss.n4038 0.095
R22663 vss.n4051 vss.n4049 0.095
R22664 vss.n4062 vss.n4060 0.095
R22665 vss.n4073 vss.n4071 0.095
R22666 vss.n4084 vss.n4082 0.095
R22667 vss.n4095 vss.n4093 0.095
R22668 vss.n17342 vss.n17340 0.095
R22669 vss.n17353 vss.n17351 0.095
R22670 vss.n17364 vss.n17362 0.095
R22671 vss.n17375 vss.n17373 0.095
R22672 vss.n17386 vss.n17384 0.095
R22673 vss.n17397 vss.n17395 0.095
R22674 vss.n21820 vss.n21819 0.094
R22675 vss.n3769 vss.n3768 0.094
R22676 vss.n21965 vss.n21964 0.092
R22677 vss.n3914 vss.n3913 0.092
R22678 vss.n16674 vss.n16661 0.091
R22679 vss.n9673 vss.n9672 0.09
R22680 vss.n14408 vss.n14407 0.09
R22681 vss.n13306 vss.n13305 0.09
R22682 vss.n21938 vss.n21937 0.089
R22683 vss.n3887 vss.n3886 0.089
R22684 vss.n20376 vss.n20374 0.089
R22685 vss.n6986 vss.n6984 0.089
R22686 vss.n18958 vss.n17680 0.088
R22687 vss.n18941 vss.n17687 0.088
R22688 vss.n17784 vss.n17783 0.088
R22689 vss.n17796 vss.n17793 0.088
R22690 vss.n18712 vss.n17891 0.088
R22691 vss.n18700 vss.n17897 0.088
R22692 vss.n17997 vss.n17996 0.088
R22693 vss.n18009 vss.n18006 0.088
R22694 vss.n18471 vss.n18104 0.088
R22695 vss.n18459 vss.n18110 0.088
R22696 vss.n18210 vss.n18209 0.088
R22697 vss.n18222 vss.n18219 0.088
R22698 vss.n19611 vss.n17587 0.088
R22699 vss.n19084 vss.n19083 0.088
R22700 vss.n19096 vss.n19093 0.088
R22701 vss.n20104 vss.n19187 0.088
R22702 vss.n20087 vss.n19194 0.088
R22703 vss.n19291 vss.n19290 0.088
R22704 vss.n19303 vss.n19300 0.088
R22705 vss.n19857 vss.n19394 0.088
R22706 vss.n19840 vss.n19400 0.088
R22707 vss.n19498 vss.n19497 0.088
R22708 vss.n19510 vss.n19507 0.088
R22709 vss.n5568 vss.n4290 0.088
R22710 vss.n5551 vss.n4297 0.088
R22711 vss.n4394 vss.n4393 0.088
R22712 vss.n4406 vss.n4403 0.088
R22713 vss.n5322 vss.n4501 0.088
R22714 vss.n5310 vss.n4507 0.088
R22715 vss.n4607 vss.n4606 0.088
R22716 vss.n4619 vss.n4616 0.088
R22717 vss.n5081 vss.n4714 0.088
R22718 vss.n5069 vss.n4720 0.088
R22719 vss.n4820 vss.n4819 0.088
R22720 vss.n4832 vss.n4829 0.088
R22721 vss.n6221 vss.n4197 0.088
R22722 vss.n5694 vss.n5693 0.088
R22723 vss.n5706 vss.n5703 0.088
R22724 vss.n6714 vss.n5797 0.088
R22725 vss.n6697 vss.n5804 0.088
R22726 vss.n5901 vss.n5900 0.088
R22727 vss.n5913 vss.n5910 0.088
R22728 vss.n6467 vss.n6004 0.088
R22729 vss.n6450 vss.n6010 0.088
R22730 vss.n6108 vss.n6107 0.088
R22731 vss.n6120 vss.n6117 0.088
R22732 vss.n15882 vss.n15881 0.088
R22733 vss.n16304 vss.n16302 0.088
R22734 vss.n10382 vss.n10380 0.088
R22735 vss.n21749 vss.n21707 0.087
R22736 vss.n21756 vss.n21698 0.087
R22737 vss.n3698 vss.n3656 0.087
R22738 vss.n3705 vss.n3647 0.087
R22739 vss.n15432 vss.n15422 0.087
R22740 vss.n15548 vss.n15534 0.087
R22741 vss.n15668 vss.n15658 0.087
R22742 vss.n15782 vss.n15770 0.087
R22743 vss.n15949 vss.n15948 0.087
R22744 vss.n16074 vss.n16060 0.087
R22745 vss.n16185 vss.n16184 0.087
R22746 vss.n16379 vss.n16369 0.087
R22747 vss.n16495 vss.n16481 0.087
R22748 vss.n16615 vss.n16605 0.087
R22749 vss.n16914 vss.n16902 0.087
R22750 vss.n17017 vss.n17014 0.086
R22751 vss.n17150 vss.n17138 0.086
R22752 vss.n17253 vss.n17250 0.086
R22753 vss.n9671 vss.n9670 0.084
R22754 vss.n21989 vss.n21988 0.083
R22755 vss.n3938 vss.n3937 0.083
R22756 vss.n22049 vss.n21980 0.083
R22757 vss.n3998 vss.n3929 0.083
R22758 vss.n22034 vss.n22032 0.081
R22759 vss.n21826 vss.n21824 0.081
R22760 vss.n22031 vss.n22026 0.081
R22761 vss.n3983 vss.n3981 0.081
R22762 vss.n3775 vss.n3773 0.081
R22763 vss.n3980 vss.n3975 0.081
R22764 vss.n17568 vss.n17561 0.08
R22765 vss.n20395 vss.n20394 0.08
R22766 vss.n4178 vss.n4171 0.08
R22767 vss.n7005 vss.n7004 0.08
R22768 vss.n16265 vss.n16254 0.08
R22769 vss.n14437 vss.n14436 0.08
R22770 vss.n20411 vss.n17548 0.079
R22771 vss.n7021 vss.n4158 0.079
R22772 vss.n10431 vss.n10425 0.079
R22773 vss.n14762 vss.n14761 0.076
R22774 vss.n13805 vss.n13804 0.076
R22775 vss.n21886 vss.n21885 0.076
R22776 vss.n12105 vss.n12104 0.076
R22777 vss.n3835 vss.n3834 0.076
R22778 vss.n20397 vss.n17552 0.075
R22779 vss.n17540 vss.n17537 0.075
R22780 vss.n17495 vss.n17492 0.075
R22781 vss.n7007 vss.n4162 0.075
R22782 vss.n4150 vss.n4147 0.075
R22783 vss.n4105 vss.n4102 0.075
R22784 vss.n10334 vss.n10333 0.074
R22785 vss.n9683 vss.n9674 0.073
R22786 vss.n20397 vss.n17559 0.071
R22787 vss.n7007 vss.n4169 0.071
R22788 vss.n22002 vss.n22000 0.071
R22789 vss.n3951 vss.n3949 0.071
R22790 vss.n20395 vss.n17558 0.07
R22791 vss.n17564 vss.n17558 0.07
R22792 vss.n20306 vss.n20305 0.07
R22793 vss.n20405 vss.n17552 0.07
R22794 vss.n20405 vss.n17553 0.07
R22795 vss.n7005 vss.n4168 0.07
R22796 vss.n4174 vss.n4168 0.07
R22797 vss.n6916 vss.n6915 0.07
R22798 vss.n7015 vss.n4162 0.07
R22799 vss.n7015 vss.n4163 0.07
R22800 vss.n8933 vss.n8932 0.068
R22801 vss.n21990 vss.n21989 0.068
R22802 vss.n3939 vss.n3938 0.068
R22803 vss.n8981 vss.n8980 0.068
R22804 vss.n10419 vss.n10418 0.067
R22805 vss.n8970 vss.n8961 0.067
R22806 vss.n8945 vss.n8943 0.067
R22807 vss.n19022 vss.n17631 0.067
R22808 vss.n19006 vss.n17631 0.067
R22809 vss.n18950 vss.n18949 0.067
R22810 vss.n18891 vss.n18890 0.067
R22811 vss.n18890 vss.n17733 0.067
R22812 vss.n17794 vss.n17782 0.067
R22813 vss.n18766 vss.n17836 0.067
R22814 vss.n18766 vss.n18765 0.067
R22815 vss.n18709 vss.n18708 0.067
R22816 vss.n18650 vss.n18649 0.067
R22817 vss.n18649 vss.n17946 0.067
R22818 vss.n18007 vss.n17995 0.067
R22819 vss.n18525 vss.n18049 0.067
R22820 vss.n18525 vss.n18524 0.067
R22821 vss.n18468 vss.n18467 0.067
R22822 vss.n18409 vss.n18408 0.067
R22823 vss.n18408 vss.n18159 0.067
R22824 vss.n18220 vss.n18208 0.067
R22825 vss.n18284 vss.n18262 0.067
R22826 vss.n19044 vss.n19033 0.067
R22827 vss.n19094 vss.n19082 0.067
R22828 vss.n19142 vss.n19136 0.067
R22829 vss.n20152 vss.n19142 0.067
R22830 vss.n20096 vss.n20095 0.067
R22831 vss.n20037 vss.n20036 0.067
R22832 vss.n20036 vss.n19240 0.067
R22833 vss.n19301 vss.n19289 0.067
R22834 vss.n19349 vss.n19343 0.067
R22835 vss.n19905 vss.n19349 0.067
R22836 vss.n19849 vss.n19848 0.067
R22837 vss.n19790 vss.n19789 0.067
R22838 vss.n19789 vss.n19447 0.067
R22839 vss.n19508 vss.n19496 0.067
R22840 vss.n19556 vss.n19550 0.067
R22841 vss.n19658 vss.n19556 0.067
R22842 vss.n8946 vss.n8934 0.067
R22843 vss.n8971 vss.n8952 0.067
R22844 vss.n5632 vss.n4241 0.067
R22845 vss.n5616 vss.n4241 0.067
R22846 vss.n5560 vss.n5559 0.067
R22847 vss.n5501 vss.n5500 0.067
R22848 vss.n5500 vss.n4343 0.067
R22849 vss.n4404 vss.n4392 0.067
R22850 vss.n5376 vss.n4446 0.067
R22851 vss.n5376 vss.n5375 0.067
R22852 vss.n5319 vss.n5318 0.067
R22853 vss.n5260 vss.n5259 0.067
R22854 vss.n5259 vss.n4556 0.067
R22855 vss.n4617 vss.n4605 0.067
R22856 vss.n5135 vss.n4659 0.067
R22857 vss.n5135 vss.n5134 0.067
R22858 vss.n5078 vss.n5077 0.067
R22859 vss.n5019 vss.n5018 0.067
R22860 vss.n5018 vss.n4769 0.067
R22861 vss.n4830 vss.n4818 0.067
R22862 vss.n4894 vss.n4872 0.067
R22863 vss.n5654 vss.n5643 0.067
R22864 vss.n5704 vss.n5692 0.067
R22865 vss.n5752 vss.n5746 0.067
R22866 vss.n6762 vss.n5752 0.067
R22867 vss.n6706 vss.n6705 0.067
R22868 vss.n6647 vss.n6646 0.067
R22869 vss.n6646 vss.n5850 0.067
R22870 vss.n5911 vss.n5899 0.067
R22871 vss.n5959 vss.n5953 0.067
R22872 vss.n6515 vss.n5959 0.067
R22873 vss.n6459 vss.n6458 0.067
R22874 vss.n6400 vss.n6399 0.067
R22875 vss.n6399 vss.n6057 0.067
R22876 vss.n6118 vss.n6106 0.067
R22877 vss.n6166 vss.n6160 0.067
R22878 vss.n6268 vss.n6166 0.067
R22879 vss.n8980 vss.n8974 0.067
R22880 vss.n10297 vss.n10296 0.066
R22881 vss.n10357 vss.n10356 0.066
R22882 vss.n15371 vss.n15369 0.066
R22883 vss.n15385 vss.n15383 0.066
R22884 vss.n15399 vss.n15397 0.066
R22885 vss.n15413 vss.n15411 0.066
R22886 vss.n15446 vss.n15436 0.066
R22887 vss.n15460 vss.n15450 0.066
R22888 vss.n15474 vss.n15464 0.066
R22889 vss.n15488 vss.n15478 0.066
R22890 vss.n15502 vss.n15492 0.066
R22891 vss.n15516 vss.n15506 0.066
R22892 vss.n15530 vss.n15520 0.066
R22893 vss.n15551 vss.n15549 0.066
R22894 vss.n15565 vss.n15563 0.066
R22895 vss.n15579 vss.n15577 0.066
R22896 vss.n15593 vss.n15591 0.066
R22897 vss.n15607 vss.n15605 0.066
R22898 vss.n15621 vss.n15619 0.066
R22899 vss.n15635 vss.n15633 0.066
R22900 vss.n15649 vss.n15647 0.066
R22901 vss.n15682 vss.n15672 0.066
R22902 vss.n15696 vss.n15686 0.066
R22903 vss.n15710 vss.n15700 0.066
R22904 vss.n15724 vss.n15714 0.066
R22905 vss.n15738 vss.n15728 0.066
R22906 vss.n15752 vss.n15742 0.066
R22907 vss.n15766 vss.n15756 0.066
R22908 vss.n15835 vss.n15833 0.066
R22909 vss.n15849 vss.n15847 0.066
R22910 vss.n15863 vss.n15861 0.066
R22911 vss.n15896 vss.n15895 0.066
R22912 vss.n15910 vss.n15909 0.066
R22913 vss.n15924 vss.n15923 0.066
R22914 vss.n15938 vss.n15937 0.066
R22915 vss.n15963 vss.n15962 0.066
R22916 vss.n15977 vss.n15976 0.066
R22917 vss.n15991 vss.n15990 0.066
R22918 vss.n16005 vss.n16004 0.066
R22919 vss.n16019 vss.n16018 0.066
R22920 vss.n16033 vss.n16032 0.066
R22921 vss.n16047 vss.n16046 0.066
R22922 vss.n16076 vss.n16075 0.066
R22923 vss.n16090 vss.n16089 0.066
R22924 vss.n16104 vss.n16103 0.066
R22925 vss.n16118 vss.n16117 0.066
R22926 vss.n16132 vss.n16131 0.066
R22927 vss.n16146 vss.n16145 0.066
R22928 vss.n16160 vss.n16159 0.066
R22929 vss.n16174 vss.n16173 0.066
R22930 vss.n16199 vss.n16198 0.066
R22931 vss.n16213 vss.n16212 0.066
R22932 vss.n16227 vss.n16226 0.066
R22933 vss.n16284 vss.n16282 0.066
R22934 vss.n15273 vss.n15263 0.066
R22935 vss.n15287 vss.n15277 0.066
R22936 vss.n15301 vss.n15291 0.066
R22937 vss.n16318 vss.n16316 0.066
R22938 vss.n16332 vss.n16330 0.066
R22939 vss.n16346 vss.n16344 0.066
R22940 vss.n16360 vss.n16358 0.066
R22941 vss.n16393 vss.n16383 0.066
R22942 vss.n16407 vss.n16397 0.066
R22943 vss.n16421 vss.n16411 0.066
R22944 vss.n16435 vss.n16425 0.066
R22945 vss.n16449 vss.n16439 0.066
R22946 vss.n16463 vss.n16453 0.066
R22947 vss.n16477 vss.n16467 0.066
R22948 vss.n16498 vss.n16496 0.066
R22949 vss.n16512 vss.n16510 0.066
R22950 vss.n16526 vss.n16524 0.066
R22951 vss.n16540 vss.n16538 0.066
R22952 vss.n16554 vss.n16552 0.066
R22953 vss.n16568 vss.n16566 0.066
R22954 vss.n16582 vss.n16580 0.066
R22955 vss.n16596 vss.n16594 0.066
R22956 vss.n16629 vss.n16619 0.066
R22957 vss.n16643 vss.n16633 0.066
R22958 vss.n16657 vss.n16647 0.066
R22959 vss.n16698 vss.n16686 0.066
R22960 vss.n16712 vss.n16700 0.066
R22961 vss.n16726 vss.n16714 0.066
R22962 vss.n16740 vss.n16728 0.066
R22963 vss.n16754 vss.n16742 0.066
R22964 vss.n16850 vss.n16849 0.066
R22965 vss.n16864 vss.n16863 0.066
R22966 vss.n16878 vss.n16877 0.066
R22967 vss.n16892 vss.n16891 0.066
R22968 vss.n16928 vss.n16916 0.066
R22969 vss.n16942 vss.n16930 0.066
R22970 vss.n16956 vss.n16944 0.066
R22971 vss.n16970 vss.n16958 0.066
R22972 vss.n16984 vss.n16972 0.066
R22973 vss.n16998 vss.n16986 0.066
R22974 vss.n17012 vss.n17000 0.066
R22975 vss.n18284 vss.n18283 0.065
R22976 vss.n20288 vss.n19033 0.065
R22977 vss.n20542 vss.n20538 0.065
R22978 vss.n20544 vss.n20542 0.065
R22979 vss.n21748 vss.n21709 0.065
R22980 vss.n10275 vss.n10264 0.065
R22981 vss.n10570 vss.n10567 0.065
R22982 vss.n10724 vss.n10722 0.065
R22983 vss.n12994 vss.n12972 0.065
R22984 vss.n13013 vss.n13012 0.065
R22985 vss.n3697 vss.n3658 0.065
R22986 vss.n4894 vss.n4893 0.065
R22987 vss.n6898 vss.n5643 0.065
R22988 vss.n7152 vss.n7148 0.065
R22989 vss.n7154 vss.n7152 0.065
R22990 vss.n17030 vss.n17029 0.065
R22991 vss.n17044 vss.n17043 0.065
R22992 vss.n17058 vss.n17057 0.065
R22993 vss.n17072 vss.n17071 0.065
R22994 vss.n17086 vss.n17085 0.065
R22995 vss.n17100 vss.n17099 0.065
R22996 vss.n17114 vss.n17113 0.065
R22997 vss.n17128 vss.n17127 0.065
R22998 vss.n17164 vss.n17152 0.065
R22999 vss.n17178 vss.n17166 0.065
R23000 vss.n17192 vss.n17180 0.065
R23001 vss.n17206 vss.n17194 0.065
R23002 vss.n17220 vss.n17208 0.065
R23003 vss.n17234 vss.n17222 0.065
R23004 vss.n17248 vss.n17236 0.065
R23005 vss.n21752 vss.n21751 0.064
R23006 vss.n3701 vss.n3700 0.064
R23007 vss.n21819 vss.n21818 0.064
R23008 vss.n3768 vss.n3767 0.064
R23009 vss.n10319 vss.n10306 0.064
R23010 vss.n9009 vss.n9008 0.063
R23011 vss.n16251 vss.n16250 0.063
R23012 vss.n11471 vss.n11470 0.063
R23013 vss.n13679 vss.n13678 0.063
R23014 vss.n13138 vss.n13137 0.063
R23015 vss.n13129 vss.n13128 0.063
R23016 vss.n12403 vss.n12402 0.063
R23017 vss.n10666 vss.n10665 0.063
R23018 vss.n11463 vss.n11462 0.063
R23019 vss.n10658 vss.n10657 0.063
R23020 vss.n12035 vss.n12034 0.063
R23021 vss.n11315 vss.n11314 0.063
R23022 vss.n13647 vss.n13646 0.063
R23023 vss.n13963 vss.n13962 0.063
R23024 vss.n11816 vss.n11815 0.063
R23025 vss.n14713 vss.n14712 0.063
R23026 vss.n14577 vss.n14576 0.063
R23027 vss.n15005 vss.n15004 0.063
R23028 vss.n21980 vss.n21979 0.063
R23029 vss.n3929 vss.n3928 0.063
R23030 vss.n13450 vss.n13449 0.063
R23031 vss.n13027 vss.n13024 0.063
R23032 vss.n10582 vss.n10581 0.063
R23033 vss.n10741 vss.n10738 0.063
R23034 vss.n13637 vss.n13636 0.063
R23035 vss.n13691 vss.n13688 0.063
R23036 vss.n11386 vss.n11385 0.063
R23037 vss.n11374 vss.n11371 0.063
R23038 vss.n11689 vss.n11680 0.063
R23039 vss.n12263 vss.n12255 0.063
R23040 vss.n11939 vss.n11931 0.063
R23041 vss.n13949 vss.n13942 0.063
R23042 vss.n10254 vss.n10253 0.063
R23043 vss.n20385 vss.n20384 0.062
R23044 vss.n6995 vss.n6994 0.062
R23045 vss.n20397 vss.n17551 0.062
R23046 vss.n20454 vss.n20443 0.062
R23047 vss.n22009 vss.n22007 0.062
R23048 vss.n22031 vss.n22014 0.062
R23049 vss.n21622 vss.n21621 0.062
R23050 vss.n9177 vss.n9171 0.062
R23051 vss.n10294 vss.n10283 0.062
R23052 vss.n3958 vss.n3956 0.062
R23053 vss.n3980 vss.n3963 0.062
R23054 vss.n3571 vss.n3570 0.062
R23055 vss.n7007 vss.n4161 0.062
R23056 vss.n7064 vss.n7053 0.062
R23057 vss.n21895 vss.n21894 0.062
R23058 vss.n3844 vss.n3843 0.062
R23059 vss.n14390 vss.n14389 0.061
R23060 vss.n13288 vss.n13287 0.061
R23061 vss.n13842 vss.n13841 0.061
R23062 vss.n13968 vss.n13967 0.061
R23063 vss.n12567 vss.n12566 0.061
R23064 vss.n12060 vss.n12059 0.061
R23065 vss.n10525 vss.n10524 0.061
R23066 vss.n10922 vss.n10921 0.061
R23067 vss.n11031 vss.n11030 0.061
R23068 vss.n13187 vss.n13186 0.061
R23069 vss.n10342 vss.n10341 0.061
R23070 vss.n12300 vss.n12289 0.061
R23071 vss.n13499 vss.n13488 0.061
R23072 vss.n13183 vss.n13182 0.061
R23073 vss.n12393 vss.n12381 0.061
R23074 vss.n13818 vss.n13816 0.061
R23075 vss.n11554 vss.n11541 0.061
R23076 vss.n9093 vss.n9075 0.061
R23077 vss.n9001 vss.n8983 0.061
R23078 vss.n9031 vss.n9013 0.06
R23079 vss.n9151 vss.n9150 0.06
R23080 vss.n9062 vss.n9044 0.06
R23081 vss.n9124 vss.n9123 0.06
R23082 vss.n21976 vss.n21973 0.06
R23083 vss.n10222 vss.n10221 0.06
R23084 vss.n10792 vss.n10779 0.06
R23085 vss.n13420 vss.n13407 0.06
R23086 vss.n12953 vss.n12941 0.06
R23087 vss.n12355 vss.n12352 0.06
R23088 vss.n13798 vss.n13776 0.06
R23089 vss.n11524 vss.n11512 0.06
R23090 vss.n3925 vss.n3922 0.06
R23091 vss.n17317 vss.n17265 0.06
R23092 vss.n20384 vss.n20383 0.06
R23093 vss.n6994 vss.n6993 0.06
R23094 vss.n12102 vss.n12101 0.059
R23095 vss.n13283 vss.n13282 0.059
R23096 vss.n10380 vss.n10379 0.059
R23097 vss.n21754 vss.n21700 0.059
R23098 vss.n12536 vss.n12535 0.059
R23099 vss.n3703 vss.n3649 0.059
R23100 vss.n9120 vss.n9119 0.059
R23101 vss.n11237 vss.n11236 0.059
R23102 vss.n10871 vss.n10869 0.059
R23103 vss.n13524 vss.n13523 0.059
R23104 vss.n14180 vss.n14178 0.059
R23105 vss.n21616 vss.n21615 0.058
R23106 vss.n3565 vss.n3564 0.058
R23107 vss.n7504 vss.n7503 0.058
R23108 vss.n9673 vss.n9667 0.058
R23109 vss.n10241 vss.n10240 0.058
R23110 vss.n10266 vss.n10265 0.058
R23111 vss.n10285 vss.n10284 0.058
R23112 vss.n10308 vss.n10307 0.058
R23113 vss.n10326 vss.n10325 0.058
R23114 vss.n10368 vss.n10367 0.058
R23115 vss.n10400 vss.n10399 0.058
R23116 vss.n10434 vss.n10433 0.058
R23117 vss.n8941 vss.n8940 0.058
R23118 vss.n8959 vss.n8958 0.058
R23119 vss.n8990 vss.n8989 0.058
R23120 vss.n9020 vss.n9019 0.058
R23121 vss.n9051 vss.n9050 0.058
R23122 vss.n9082 vss.n9081 0.058
R23123 vss.n9101 vss.n9100 0.058
R23124 vss.n9131 vss.n9130 0.058
R23125 vss.n8923 vss.n8922 0.057
R23126 vss.n8932 vss.n8931 0.057
R23127 vss.n21785 vss.n21774 0.057
R23128 vss.n3734 vss.n3723 0.057
R23129 vss.n21759 vss.n21703 0.057
R23130 vss.n12106 vss.n12105 0.057
R23131 vss.n3708 vss.n3652 0.057
R23132 vss.n8129 vss.n8128 0.057
R23133 vss.n8027 vss.n8026 0.057
R23134 vss.n8026 vss.n8022 0.057
R23135 vss.n7921 vss.n7920 0.057
R23136 vss.n7818 vss.n7817 0.057
R23137 vss.n7817 vss.n7813 0.057
R23138 vss.n7712 vss.n7711 0.057
R23139 vss.n7610 vss.n7609 0.057
R23140 vss.n7609 vss.n7605 0.057
R23141 vss.n8948 vss.n8947 0.057
R23142 vss.n9665 vss.n9664 0.056
R23143 vss.n20391 vss.n20390 0.056
R23144 vss.n21917 vss.n21916 0.056
R23145 vss.n21748 vss.n21706 0.056
R23146 vss.n3866 vss.n3865 0.056
R23147 vss.n3697 vss.n3655 0.056
R23148 vss.n7001 vss.n7000 0.056
R23149 vss.n8920 vss.n8918 0.056
R23150 vss.n22757 vss.n22755 0.056
R23151 vss.n20894 vss.n20893 0.055
R23152 vss.n10387 vss.n10386 0.055
R23153 vss.n21671 vss.n21661 0.054
R23154 vss.n3620 vss.n3610 0.054
R23155 vss.n21518 vss.n21517 0.054
R23156 vss.n21416 vss.n21415 0.054
R23157 vss.n21415 vss.n21411 0.054
R23158 vss.n21310 vss.n21309 0.054
R23159 vss.n21208 vss.n21207 0.054
R23160 vss.n21207 vss.n21203 0.054
R23161 vss.n21102 vss.n21101 0.054
R23162 vss.n21000 vss.n20999 0.054
R23163 vss.n20999 vss.n20995 0.054
R23164 vss.n21794 vss.n21684 0.054
R23165 vss.n21722 vss.n21688 0.054
R23166 vss.n21792 vss.n21687 0.054
R23167 vss.n3743 vss.n3633 0.054
R23168 vss.n3671 vss.n3637 0.054
R23169 vss.n3741 vss.n3636 0.054
R23170 vss.n8859 vss.n8858 0.054
R23171 vss.n8858 vss.n8854 0.054
R23172 vss.n8753 vss.n8752 0.054
R23173 vss.n8651 vss.n8650 0.054
R23174 vss.n8650 vss.n8646 0.054
R23175 vss.n8545 vss.n8544 0.054
R23176 vss.n8443 vss.n8442 0.054
R23177 vss.n8442 vss.n8438 0.054
R23178 vss.n8337 vss.n8336 0.054
R23179 vss.n22696 vss.n22695 0.054
R23180 vss.n22695 vss.n22691 0.054
R23181 vss.n22590 vss.n22589 0.054
R23182 vss.n22488 vss.n22487 0.054
R23183 vss.n22487 vss.n22483 0.054
R23184 vss.n22382 vss.n22381 0.054
R23185 vss.n22280 vss.n22279 0.054
R23186 vss.n22279 vss.n22275 0.054
R23187 vss.n22174 vss.n22173 0.054
R23188 vss.n20375 vss.n17573 0.054
R23189 vss.n6985 vss.n4183 0.054
R23190 vss.n10318 vss.n10315 0.053
R23191 vss.n20391 vss.n17558 0.053
R23192 vss.n20392 vss.n17562 0.053
R23193 vss.n21635 vss.n21634 0.053
R23194 vss.n10446 vss.n10445 0.053
R23195 vss.n7001 vss.n4168 0.053
R23196 vss.n7002 vss.n4172 0.053
R23197 vss.n3584 vss.n3583 0.053
R23198 vss.n15209 vss.n3426 0.053
R23199 vss.n22842 vss.n22841 0.053
R23200 vss.n21652 vss.n21645 0.053
R23201 vss.n3601 vss.n3594 0.053
R23202 vss.n20390 vss.n20389 0.053
R23203 vss.n7000 vss.n6999 0.053
R23204 vss.n8969 vss.n8968 0.052
R23205 vss.n19031 vss.n17623 0.052
R23206 vss.n20290 vss.n19032 0.052
R23207 vss.n5641 vss.n4233 0.052
R23208 vss.n6900 vss.n5642 0.052
R23209 vss.n13309 bandgapmd_0.pnp_groupm_0.vss 0.052
R23210 vss.n14929 vss.n14927 0.052
R23211 vss.n21747 vss.n21710 0.051
R23212 vss.n3696 vss.n3659 0.051
R23213 vss.n20397 vss.n20396 0.051
R23214 vss.n10230 vss.n10229 0.051
R23215 vss.n7007 vss.n7006 0.051
R23216 vss.n10274 vss.n10272 0.051
R23217 vss.n22068 vss.n22067 0.05
R23218 vss.n19004 vss.n17641 0.05
R23219 vss.n17651 vss.n17650 0.05
R23220 vss.n18985 vss.n17659 0.05
R23221 vss.n18983 vss.n17660 0.05
R23222 vss.n18972 vss.n18971 0.05
R23223 vss.n18962 vss.n17678 0.05
R23224 vss.n18960 vss.n17679 0.05
R23225 vss.n18948 vss.n17686 0.05
R23226 vss.n18937 vss.n18936 0.05
R23227 vss.n18925 vss.n17695 0.05
R23228 vss.n18923 vss.n17705 0.05
R23229 vss.n18914 vss.n18913 0.05
R23230 vss.n18902 vss.n17717 0.05
R23231 vss.n18900 vss.n17724 0.05
R23232 vss.n18879 vss.n18878 0.05
R23233 vss.n18869 vss.n17756 0.05
R23234 vss.n18867 vss.n17757 0.05
R23235 vss.n18856 vss.n18855 0.05
R23236 vss.n18846 vss.n17775 0.05
R23237 vss.n18844 vss.n17776 0.05
R23238 vss.n18833 vss.n18832 0.05
R23239 vss.n18824 vss.n18823 0.05
R23240 vss.n18812 vss.n17798 0.05
R23241 vss.n18810 vss.n17805 0.05
R23242 vss.n18801 vss.n18800 0.05
R23243 vss.n18789 vss.n17817 0.05
R23244 vss.n18787 vss.n17824 0.05
R23245 vss.n18778 vss.n18777 0.05
R23246 vss.n18756 vss.n17856 0.05
R23247 vss.n18754 vss.n17857 0.05
R23248 vss.n18743 vss.n18742 0.05
R23249 vss.n18733 vss.n17875 0.05
R23250 vss.n18731 vss.n17876 0.05
R23251 vss.n18720 vss.n18719 0.05
R23252 vss.n18710 vss.n17894 0.05
R23253 vss.n18707 vss.n17896 0.05
R23254 vss.n18696 vss.n18695 0.05
R23255 vss.n18684 vss.n17908 0.05
R23256 vss.n18682 vss.n17918 0.05
R23257 vss.n18673 vss.n18672 0.05
R23258 vss.n18661 vss.n17930 0.05
R23259 vss.n18659 vss.n17937 0.05
R23260 vss.n18638 vss.n18637 0.05
R23261 vss.n18628 vss.n17969 0.05
R23262 vss.n18626 vss.n17970 0.05
R23263 vss.n18615 vss.n18614 0.05
R23264 vss.n18605 vss.n17988 0.05
R23265 vss.n18603 vss.n17989 0.05
R23266 vss.n18592 vss.n18591 0.05
R23267 vss.n18583 vss.n18582 0.05
R23268 vss.n18571 vss.n18011 0.05
R23269 vss.n18569 vss.n18018 0.05
R23270 vss.n18560 vss.n18559 0.05
R23271 vss.n18548 vss.n18030 0.05
R23272 vss.n18546 vss.n18037 0.05
R23273 vss.n18537 vss.n18536 0.05
R23274 vss.n18515 vss.n18069 0.05
R23275 vss.n18513 vss.n18070 0.05
R23276 vss.n18502 vss.n18501 0.05
R23277 vss.n18492 vss.n18088 0.05
R23278 vss.n18490 vss.n18089 0.05
R23279 vss.n18479 vss.n18478 0.05
R23280 vss.n18469 vss.n18107 0.05
R23281 vss.n18466 vss.n18109 0.05
R23282 vss.n18455 vss.n18454 0.05
R23283 vss.n18443 vss.n18121 0.05
R23284 vss.n18441 vss.n18131 0.05
R23285 vss.n18432 vss.n18431 0.05
R23286 vss.n18420 vss.n18143 0.05
R23287 vss.n18418 vss.n18150 0.05
R23288 vss.n18397 vss.n18396 0.05
R23289 vss.n18387 vss.n18182 0.05
R23290 vss.n18385 vss.n18183 0.05
R23291 vss.n18374 vss.n18373 0.05
R23292 vss.n18364 vss.n18201 0.05
R23293 vss.n18362 vss.n18202 0.05
R23294 vss.n18351 vss.n18350 0.05
R23295 vss.n18342 vss.n18341 0.05
R23296 vss.n18330 vss.n18224 0.05
R23297 vss.n18328 vss.n18231 0.05
R23298 vss.n18319 vss.n18318 0.05
R23299 vss.n18307 vss.n18243 0.05
R23300 vss.n18305 vss.n18250 0.05
R23301 vss.n18296 vss.n18295 0.05
R23302 vss.n19048 vss.n19047 0.05
R23303 vss.n20262 vss.n19056 0.05
R23304 vss.n20260 vss.n19057 0.05
R23305 vss.n20249 vss.n20248 0.05
R23306 vss.n20239 vss.n19075 0.05
R23307 vss.n20237 vss.n19076 0.05
R23308 vss.n20226 vss.n20225 0.05
R23309 vss.n20217 vss.n20216 0.05
R23310 vss.n20205 vss.n19098 0.05
R23311 vss.n20203 vss.n19105 0.05
R23312 vss.n20194 vss.n20193 0.05
R23313 vss.n20182 vss.n19117 0.05
R23314 vss.n20180 vss.n19124 0.05
R23315 vss.n20171 vss.n20170 0.05
R23316 vss.n20150 vss.n19148 0.05
R23317 vss.n19158 vss.n19157 0.05
R23318 vss.n20131 vss.n19166 0.05
R23319 vss.n20129 vss.n19167 0.05
R23320 vss.n20118 vss.n20117 0.05
R23321 vss.n20108 vss.n19185 0.05
R23322 vss.n20106 vss.n19186 0.05
R23323 vss.n20094 vss.n19193 0.05
R23324 vss.n20083 vss.n20082 0.05
R23325 vss.n20071 vss.n19202 0.05
R23326 vss.n20069 vss.n19212 0.05
R23327 vss.n20060 vss.n20059 0.05
R23328 vss.n20048 vss.n19224 0.05
R23329 vss.n20046 vss.n19231 0.05
R23330 vss.n20025 vss.n20024 0.05
R23331 vss.n20015 vss.n19263 0.05
R23332 vss.n20013 vss.n19264 0.05
R23333 vss.n20002 vss.n20001 0.05
R23334 vss.n19992 vss.n19282 0.05
R23335 vss.n19990 vss.n19283 0.05
R23336 vss.n19979 vss.n19978 0.05
R23337 vss.n19970 vss.n19969 0.05
R23338 vss.n19958 vss.n19305 0.05
R23339 vss.n19956 vss.n19312 0.05
R23340 vss.n19947 vss.n19946 0.05
R23341 vss.n19935 vss.n19324 0.05
R23342 vss.n19933 vss.n19331 0.05
R23343 vss.n19924 vss.n19923 0.05
R23344 vss.n19903 vss.n19355 0.05
R23345 vss.n19365 vss.n19364 0.05
R23346 vss.n19884 vss.n19373 0.05
R23347 vss.n19882 vss.n19374 0.05
R23348 vss.n19871 vss.n19870 0.05
R23349 vss.n19861 vss.n19392 0.05
R23350 vss.n19859 vss.n19393 0.05
R23351 vss.n19847 vss.n19399 0.05
R23352 vss.n19836 vss.n19835 0.05
R23353 vss.n19824 vss.n19409 0.05
R23354 vss.n19822 vss.n19419 0.05
R23355 vss.n19813 vss.n19812 0.05
R23356 vss.n19801 vss.n19431 0.05
R23357 vss.n19799 vss.n19438 0.05
R23358 vss.n19778 vss.n19777 0.05
R23359 vss.n19768 vss.n19470 0.05
R23360 vss.n19766 vss.n19471 0.05
R23361 vss.n19755 vss.n19754 0.05
R23362 vss.n19745 vss.n19489 0.05
R23363 vss.n19743 vss.n19490 0.05
R23364 vss.n19732 vss.n19731 0.05
R23365 vss.n19723 vss.n19722 0.05
R23366 vss.n19711 vss.n19512 0.05
R23367 vss.n19709 vss.n19519 0.05
R23368 vss.n19700 vss.n19699 0.05
R23369 vss.n19688 vss.n19531 0.05
R23370 vss.n19686 vss.n19538 0.05
R23371 vss.n19677 vss.n19676 0.05
R23372 vss.n19656 vss.n19562 0.05
R23373 vss.n19572 vss.n19571 0.05
R23374 vss.n19637 vss.n19580 0.05
R23375 vss.n19635 vss.n19581 0.05
R23376 vss.n21783 vss.n21781 0.05
R23377 vss.n21777 vss.n21685 0.05
R23378 vss.n10238 vss.n10237 0.05
R23379 vss.n14143 vss.n14141 0.05
R23380 vss.n11883 vss.n11881 0.05
R23381 vss.n3732 vss.n3730 0.05
R23382 vss.n3726 vss.n3634 0.05
R23383 vss.n5614 vss.n4251 0.05
R23384 vss.n4261 vss.n4260 0.05
R23385 vss.n5595 vss.n4269 0.05
R23386 vss.n5593 vss.n4270 0.05
R23387 vss.n5582 vss.n5581 0.05
R23388 vss.n5572 vss.n4288 0.05
R23389 vss.n5570 vss.n4289 0.05
R23390 vss.n5558 vss.n4296 0.05
R23391 vss.n5547 vss.n5546 0.05
R23392 vss.n5535 vss.n4305 0.05
R23393 vss.n5533 vss.n4315 0.05
R23394 vss.n5524 vss.n5523 0.05
R23395 vss.n5512 vss.n4327 0.05
R23396 vss.n5510 vss.n4334 0.05
R23397 vss.n5489 vss.n5488 0.05
R23398 vss.n5479 vss.n4366 0.05
R23399 vss.n5477 vss.n4367 0.05
R23400 vss.n5466 vss.n5465 0.05
R23401 vss.n5456 vss.n4385 0.05
R23402 vss.n5454 vss.n4386 0.05
R23403 vss.n5443 vss.n5442 0.05
R23404 vss.n5434 vss.n5433 0.05
R23405 vss.n5422 vss.n4408 0.05
R23406 vss.n5420 vss.n4415 0.05
R23407 vss.n5411 vss.n5410 0.05
R23408 vss.n5399 vss.n4427 0.05
R23409 vss.n5397 vss.n4434 0.05
R23410 vss.n5388 vss.n5387 0.05
R23411 vss.n5366 vss.n4466 0.05
R23412 vss.n5364 vss.n4467 0.05
R23413 vss.n5353 vss.n5352 0.05
R23414 vss.n5343 vss.n4485 0.05
R23415 vss.n5341 vss.n4486 0.05
R23416 vss.n5330 vss.n5329 0.05
R23417 vss.n5320 vss.n4504 0.05
R23418 vss.n5317 vss.n4506 0.05
R23419 vss.n5306 vss.n5305 0.05
R23420 vss.n5294 vss.n4518 0.05
R23421 vss.n5292 vss.n4528 0.05
R23422 vss.n5283 vss.n5282 0.05
R23423 vss.n5271 vss.n4540 0.05
R23424 vss.n5269 vss.n4547 0.05
R23425 vss.n5248 vss.n5247 0.05
R23426 vss.n5238 vss.n4579 0.05
R23427 vss.n5236 vss.n4580 0.05
R23428 vss.n5225 vss.n5224 0.05
R23429 vss.n5215 vss.n4598 0.05
R23430 vss.n5213 vss.n4599 0.05
R23431 vss.n5202 vss.n5201 0.05
R23432 vss.n5193 vss.n5192 0.05
R23433 vss.n5181 vss.n4621 0.05
R23434 vss.n5179 vss.n4628 0.05
R23435 vss.n5170 vss.n5169 0.05
R23436 vss.n5158 vss.n4640 0.05
R23437 vss.n5156 vss.n4647 0.05
R23438 vss.n5147 vss.n5146 0.05
R23439 vss.n5125 vss.n4679 0.05
R23440 vss.n5123 vss.n4680 0.05
R23441 vss.n5112 vss.n5111 0.05
R23442 vss.n5102 vss.n4698 0.05
R23443 vss.n5100 vss.n4699 0.05
R23444 vss.n5089 vss.n5088 0.05
R23445 vss.n5079 vss.n4717 0.05
R23446 vss.n5076 vss.n4719 0.05
R23447 vss.n5065 vss.n5064 0.05
R23448 vss.n5053 vss.n4731 0.05
R23449 vss.n5051 vss.n4741 0.05
R23450 vss.n5042 vss.n5041 0.05
R23451 vss.n5030 vss.n4753 0.05
R23452 vss.n5028 vss.n4760 0.05
R23453 vss.n5007 vss.n5006 0.05
R23454 vss.n4997 vss.n4792 0.05
R23455 vss.n4995 vss.n4793 0.05
R23456 vss.n4984 vss.n4983 0.05
R23457 vss.n4974 vss.n4811 0.05
R23458 vss.n4972 vss.n4812 0.05
R23459 vss.n4961 vss.n4960 0.05
R23460 vss.n4952 vss.n4951 0.05
R23461 vss.n4940 vss.n4834 0.05
R23462 vss.n4938 vss.n4841 0.05
R23463 vss.n4929 vss.n4928 0.05
R23464 vss.n4917 vss.n4853 0.05
R23465 vss.n4915 vss.n4860 0.05
R23466 vss.n4906 vss.n4905 0.05
R23467 vss.n5658 vss.n5657 0.05
R23468 vss.n6872 vss.n5666 0.05
R23469 vss.n6870 vss.n5667 0.05
R23470 vss.n6859 vss.n6858 0.05
R23471 vss.n6849 vss.n5685 0.05
R23472 vss.n6847 vss.n5686 0.05
R23473 vss.n6836 vss.n6835 0.05
R23474 vss.n6827 vss.n6826 0.05
R23475 vss.n6815 vss.n5708 0.05
R23476 vss.n6813 vss.n5715 0.05
R23477 vss.n6804 vss.n6803 0.05
R23478 vss.n6792 vss.n5727 0.05
R23479 vss.n6790 vss.n5734 0.05
R23480 vss.n6781 vss.n6780 0.05
R23481 vss.n6760 vss.n5758 0.05
R23482 vss.n5768 vss.n5767 0.05
R23483 vss.n6741 vss.n5776 0.05
R23484 vss.n6739 vss.n5777 0.05
R23485 vss.n6728 vss.n6727 0.05
R23486 vss.n6718 vss.n5795 0.05
R23487 vss.n6716 vss.n5796 0.05
R23488 vss.n6704 vss.n5803 0.05
R23489 vss.n6693 vss.n6692 0.05
R23490 vss.n6681 vss.n5812 0.05
R23491 vss.n6679 vss.n5822 0.05
R23492 vss.n6670 vss.n6669 0.05
R23493 vss.n6658 vss.n5834 0.05
R23494 vss.n6656 vss.n5841 0.05
R23495 vss.n6635 vss.n6634 0.05
R23496 vss.n6625 vss.n5873 0.05
R23497 vss.n6623 vss.n5874 0.05
R23498 vss.n6612 vss.n6611 0.05
R23499 vss.n6602 vss.n5892 0.05
R23500 vss.n6600 vss.n5893 0.05
R23501 vss.n6589 vss.n6588 0.05
R23502 vss.n6580 vss.n6579 0.05
R23503 vss.n6568 vss.n5915 0.05
R23504 vss.n6566 vss.n5922 0.05
R23505 vss.n6557 vss.n6556 0.05
R23506 vss.n6545 vss.n5934 0.05
R23507 vss.n6543 vss.n5941 0.05
R23508 vss.n6534 vss.n6533 0.05
R23509 vss.n6513 vss.n5965 0.05
R23510 vss.n5975 vss.n5974 0.05
R23511 vss.n6494 vss.n5983 0.05
R23512 vss.n6492 vss.n5984 0.05
R23513 vss.n6481 vss.n6480 0.05
R23514 vss.n6471 vss.n6002 0.05
R23515 vss.n6469 vss.n6003 0.05
R23516 vss.n6457 vss.n6009 0.05
R23517 vss.n6446 vss.n6445 0.05
R23518 vss.n6434 vss.n6019 0.05
R23519 vss.n6432 vss.n6029 0.05
R23520 vss.n6423 vss.n6422 0.05
R23521 vss.n6411 vss.n6041 0.05
R23522 vss.n6409 vss.n6048 0.05
R23523 vss.n6388 vss.n6387 0.05
R23524 vss.n6378 vss.n6080 0.05
R23525 vss.n6376 vss.n6081 0.05
R23526 vss.n6365 vss.n6364 0.05
R23527 vss.n6355 vss.n6099 0.05
R23528 vss.n6353 vss.n6100 0.05
R23529 vss.n6342 vss.n6341 0.05
R23530 vss.n6333 vss.n6332 0.05
R23531 vss.n6321 vss.n6122 0.05
R23532 vss.n6319 vss.n6129 0.05
R23533 vss.n6310 vss.n6309 0.05
R23534 vss.n6298 vss.n6141 0.05
R23535 vss.n6296 vss.n6148 0.05
R23536 vss.n6287 vss.n6286 0.05
R23537 vss.n6266 vss.n6172 0.05
R23538 vss.n6182 vss.n6181 0.05
R23539 vss.n6247 vss.n6190 0.05
R23540 vss.n6245 vss.n6191 0.05
R23541 vss.n20386 vss.n17567 0.05
R23542 vss.n6996 vss.n4177 0.05
R23543 vss.n17563 vss.n17557 0.049
R23544 vss.n20470 vss.n20459 0.049
R23545 vss.n20485 vss.n20474 0.049
R23546 vss.n20500 vss.n20489 0.049
R23547 vss.n20534 vss.n20520 0.049
R23548 vss.n20563 vss.n20561 0.049
R23549 vss.n20578 vss.n20576 0.049
R23550 vss.n9674 vss.n9156 0.049
R23551 vss.n10451 vss.n10448 0.049
R23552 vss.n4173 vss.n4167 0.049
R23553 vss.n7080 vss.n7069 0.049
R23554 vss.n7095 vss.n7084 0.049
R23555 vss.n7110 vss.n7099 0.049
R23556 vss.n7144 vss.n7130 0.049
R23557 vss.n7173 vss.n7171 0.049
R23558 vss.n7188 vss.n7186 0.049
R23559 vss.n8918 vss.n8916 0.049
R23560 vss.n22755 vss.n22753 0.049
R23561 vss.n17570 vss.n17566 0.048
R23562 vss.n4180 vss.n4176 0.048
R23563 vss.n21754 vss.n21697 0.048
R23564 vss.n14823 vss.n14821 0.048
R23565 vss.n12761 vss.n12760 0.048
R23566 vss.n12764 vss.n12763 0.048
R23567 vss.n15074 vss.n15073 0.048
R23568 vss.n15071 vss.n15070 0.048
R23569 vss.n3703 vss.n3646 0.048
R23570 vss.n15819 vss.n15783 0.048
R23571 vss.n8981 vss.n8973 0.047
R23572 vss.n20388 vss.n17565 0.047
R23573 vss.n6998 vss.n4175 0.047
R23574 vss.n9674 vss.n9662 0.046
R23575 vss.n20390 vss.n17564 0.046
R23576 vss.n21889 vss.n21888 0.046
R23577 vss.n10322 vss.n10321 0.046
R23578 vss.n3838 vss.n3837 0.046
R23579 vss.n7000 vss.n4174 0.046
R23580 vss.n3455 vss.n3435 0.046
R23581 vss.n1430 vss.n1410 0.046
R23582 vss.n10537 vss.n10536 0.046
R23583 vss.n14993 vss.n14992 0.046
R23584 vss.n17578 vss.n17576 0.045
R23585 vss.n4188 vss.n4186 0.045
R23586 vss.n17565 vss.n17558 0.045
R23587 bandgapmd_0.bg_resm_0.vss vss.t2 0.045
R23588 vss.n4175 vss.n4168 0.045
R23589 vss.n4018 vss.n4017 0.044
R23590 vss.n22063 vss.n22060 0.044
R23591 vss.n10237 vss.n10236 0.044
R23592 vss.n4012 vss.n4009 0.044
R23593 vss.n22036 vss.n22034 0.043
R23594 vss.n22043 vss.n22041 0.043
R23595 vss.n21828 vss.n21826 0.043
R23596 vss.n21846 vss.n21844 0.043
R23597 vss.n22026 vss.n22024 0.043
R23598 vss.n21975 vss.n21974 0.043
R23599 vss.n21684 vss.n21683 0.043
R23600 vss.n21675 vss.n21665 0.043
R23601 vss.n21723 vss.n21722 0.043
R23602 vss.n21738 vss.n21715 0.043
R23603 vss.n21749 vss.n21706 0.043
R23604 vss.n21762 vss.n21687 0.043
R23605 vss.n21770 vss.n21769 0.043
R23606 vss.n21703 vss.n21699 0.043
R23607 vss.n9692 bandgapmd_0.bg_trimmup_0.vss 0.043
R23608 vss.n3985 vss.n3983 0.043
R23609 vss.n3992 vss.n3990 0.043
R23610 vss.n3777 vss.n3775 0.043
R23611 vss.n3795 vss.n3793 0.043
R23612 vss.n3975 vss.n3973 0.043
R23613 vss.n3924 vss.n3923 0.043
R23614 vss.n3633 vss.n3632 0.043
R23615 vss.n3624 vss.n3614 0.043
R23616 vss.n3672 vss.n3671 0.043
R23617 vss.n3687 vss.n3664 0.043
R23618 vss.n3698 vss.n3655 0.043
R23619 vss.n3711 vss.n3636 0.043
R23620 vss.n3719 vss.n3718 0.043
R23621 vss.n3652 vss.n3648 0.043
R23622 vss.n8201 vss.n8200 0.043
R23623 vss.n8187 vss.n8186 0.043
R23624 vss.n8173 vss.n8172 0.043
R23625 vss.n8159 vss.n8158 0.043
R23626 vss.n8145 vss.n8144 0.043
R23627 vss.n8131 vss.n8130 0.043
R23628 vss.n8127 vss.n8126 0.043
R23629 vss.n8113 vss.n8112 0.043
R23630 vss.n8099 vss.n8098 0.043
R23631 vss.n8085 vss.n8084 0.043
R23632 vss.n8071 vss.n8070 0.043
R23633 vss.n8057 vss.n8056 0.043
R23634 vss.n8043 vss.n8042 0.043
R23635 vss.n8007 vss.n8006 0.043
R23636 vss.n7993 vss.n7992 0.043
R23637 vss.n7979 vss.n7978 0.043
R23638 vss.n7965 vss.n7964 0.043
R23639 vss.n7951 vss.n7950 0.043
R23640 vss.n7937 vss.n7936 0.043
R23641 vss.n7923 vss.n7922 0.043
R23642 vss.n7919 vss.n7918 0.043
R23643 vss.n7905 vss.n7904 0.043
R23644 vss.n7891 vss.n7890 0.043
R23645 vss.n7877 vss.n7876 0.043
R23646 vss.n7863 vss.n7862 0.043
R23647 vss.n7834 vss.n7833 0.043
R23648 vss.n7798 vss.n7797 0.043
R23649 vss.n7784 vss.n7783 0.043
R23650 vss.n7770 vss.n7769 0.043
R23651 vss.n7756 vss.n7755 0.043
R23652 vss.n7742 vss.n7741 0.043
R23653 vss.n7728 vss.n7727 0.043
R23654 vss.n7714 vss.n7713 0.043
R23655 vss.n7710 vss.n7709 0.043
R23656 vss.n7696 vss.n7695 0.043
R23657 vss.n7682 vss.n7681 0.043
R23658 vss.n7668 vss.n7667 0.043
R23659 vss.n7654 vss.n7653 0.043
R23660 vss.n7640 vss.n7639 0.043
R23661 vss.n7626 vss.n7625 0.043
R23662 vss.n7590 vss.n7589 0.043
R23663 vss.n7576 vss.n7575 0.043
R23664 vss.n7562 vss.n7561 0.043
R23665 vss.n7548 vss.n7547 0.043
R23666 vss.n7534 vss.n7533 0.043
R23667 vss.n7520 vss.n7519 0.043
R23668 vss.n7506 vss.n7505 0.043
R23669 vss.n15108 vss.t354 0.043
R23670 vss.n15107 vss.t332 0.043
R23671 vss.n15106 vss.t336 0.043
R23672 vss.n15105 vss.t339 0.043
R23673 vss.n15104 vss.t352 0.043
R23674 vss.n15103 vss.t344 0.043
R23675 vss.n15102 vss.t349 0.043
R23676 vss.n15101 vss.t338 0.043
R23677 vss.n15100 vss.t342 0.043
R23678 vss.n15099 vss.t333 0.043
R23679 vss.n15098 vss.t348 0.043
R23680 vss.n15119 vss.t347 0.043
R23681 vss.n15118 vss.t351 0.043
R23682 vss.n15117 vss.t331 0.043
R23683 vss.n15116 vss.t335 0.043
R23684 vss.n15115 vss.t346 0.043
R23685 vss.n15114 vss.t340 0.043
R23686 vss.n15113 vss.t343 0.043
R23687 vss.n15112 vss.t334 0.043
R23688 vss.n15111 vss.t337 0.043
R23689 vss.n15110 vss.t353 0.043
R23690 vss.n15109 vss.t341 0.043
R23691 vss.n9151 vss.n9141 0.042
R23692 vss.n9031 vss.n9030 0.042
R23693 vss.n9062 vss.n9061 0.042
R23694 vss.n9124 vss.n9112 0.042
R23695 vss.n9093 vss.n9092 0.042
R23696 vss.n17572 vss.n17571 0.042
R23697 vss.n21635 vss.n21632 0.042
R23698 vss.n21606 vss.n21605 0.042
R23699 vss.n10432 vss.n10431 0.042
R23700 vss.n4182 vss.n4181 0.042
R23701 vss.n3584 vss.n3581 0.042
R23702 vss.n15155 vss.n15125 0.042
R23703 vss.n9001 vss.n9000 0.042
R23704 vss.n19615 vss.n19614 0.041
R23705 vss.n21579 vss.n21578 0.041
R23706 vss.n21576 vss.n21575 0.041
R23707 vss.n21562 vss.n21561 0.041
R23708 vss.n21548 vss.n21547 0.041
R23709 vss.n21534 vss.n21533 0.041
R23710 vss.n21520 vss.n21519 0.041
R23711 vss.n21516 vss.n21515 0.041
R23712 vss.n21502 vss.n21501 0.041
R23713 vss.n21488 vss.n21487 0.041
R23714 vss.n21474 vss.n21473 0.041
R23715 vss.n21460 vss.n21459 0.041
R23716 vss.n21446 vss.n21445 0.041
R23717 vss.n21432 vss.n21431 0.041
R23718 vss.n21396 vss.n21395 0.041
R23719 vss.n21382 vss.n21381 0.041
R23720 vss.n21368 vss.n21367 0.041
R23721 vss.n21354 vss.n21353 0.041
R23722 vss.n21340 vss.n21339 0.041
R23723 vss.n21326 vss.n21325 0.041
R23724 vss.n21312 vss.n21311 0.041
R23725 vss.n21308 vss.n21307 0.041
R23726 vss.n21294 vss.n21293 0.041
R23727 vss.n21280 vss.n21279 0.041
R23728 vss.n21266 vss.n21265 0.041
R23729 vss.n21252 vss.n21251 0.041
R23730 vss.n21238 vss.n21237 0.041
R23731 vss.n21224 vss.n21223 0.041
R23732 vss.n21188 vss.n21187 0.041
R23733 vss.n21174 vss.n21173 0.041
R23734 vss.n21160 vss.n21159 0.041
R23735 vss.n21146 vss.n21145 0.041
R23736 vss.n21132 vss.n21131 0.041
R23737 vss.n21118 vss.n21117 0.041
R23738 vss.n21104 vss.n21103 0.041
R23739 vss.n21100 vss.n21099 0.041
R23740 vss.n21086 vss.n21085 0.041
R23741 vss.n21072 vss.n21071 0.041
R23742 vss.n21058 vss.n21057 0.041
R23743 vss.n21044 vss.n21043 0.041
R23744 vss.n21030 vss.n21029 0.041
R23745 vss.n21016 vss.n21015 0.041
R23746 vss.n20980 vss.n20979 0.041
R23747 vss.n20966 vss.n20965 0.041
R23748 vss.n20952 vss.n20951 0.041
R23749 vss.n20938 vss.n20937 0.041
R23750 vss.n20924 vss.n20923 0.041
R23751 vss.n20910 vss.n20909 0.041
R23752 vss.n20896 vss.n20895 0.041
R23753 vss.n6225 vss.n6224 0.041
R23754 vss.n8903 vss.n8902 0.041
R23755 vss.n8889 vss.n8888 0.041
R23756 vss.n8875 vss.n8874 0.041
R23757 vss.n8839 vss.n8838 0.041
R23758 vss.n8825 vss.n8824 0.041
R23759 vss.n8811 vss.n8810 0.041
R23760 vss.n8797 vss.n8796 0.041
R23761 vss.n8783 vss.n8782 0.041
R23762 vss.n8769 vss.n8768 0.041
R23763 vss.n8755 vss.n8754 0.041
R23764 vss.n8751 vss.n8750 0.041
R23765 vss.n8737 vss.n8736 0.041
R23766 vss.n8723 vss.n8722 0.041
R23767 vss.n8709 vss.n8708 0.041
R23768 vss.n8695 vss.n8694 0.041
R23769 vss.n8681 vss.n8680 0.041
R23770 vss.n8667 vss.n8666 0.041
R23771 vss.n8631 vss.n8630 0.041
R23772 vss.n8617 vss.n8616 0.041
R23773 vss.n8603 vss.n8602 0.041
R23774 vss.n8589 vss.n8588 0.041
R23775 vss.n8575 vss.n8574 0.041
R23776 vss.n8561 vss.n8560 0.041
R23777 vss.n8547 vss.n8546 0.041
R23778 vss.n8543 vss.n8542 0.041
R23779 vss.n8529 vss.n8528 0.041
R23780 vss.n8515 vss.n8514 0.041
R23781 vss.n8501 vss.n8500 0.041
R23782 vss.n8487 vss.n8486 0.041
R23783 vss.n8473 vss.n8472 0.041
R23784 vss.n8459 vss.n8458 0.041
R23785 vss.n8423 vss.n8422 0.041
R23786 vss.n8409 vss.n8408 0.041
R23787 vss.n8395 vss.n8394 0.041
R23788 vss.n8381 vss.n8380 0.041
R23789 vss.n8367 vss.n8366 0.041
R23790 vss.n8353 vss.n8352 0.041
R23791 vss.n8339 vss.n8338 0.041
R23792 vss.n8335 vss.n8334 0.041
R23793 vss.n8321 vss.n8320 0.041
R23794 vss.n8307 vss.n8306 0.041
R23795 vss.n8293 vss.n8292 0.041
R23796 vss.n8279 vss.n8278 0.041
R23797 vss.n8265 vss.n8264 0.041
R23798 vss.n8251 vss.n8250 0.041
R23799 vss.n15175 vss.n3455 0.041
R23800 vss.n15217 vss.n15212 0.041
R23801 vss.n15881 vss.n15865 0.041
R23802 vss.n16302 vss.n16293 0.041
R23803 vss.n16684 vss.n16674 0.041
R23804 vss.n22740 vss.n22739 0.041
R23805 vss.n22726 vss.n22725 0.041
R23806 vss.n22712 vss.n22711 0.041
R23807 vss.n22676 vss.n22675 0.041
R23808 vss.n22662 vss.n22661 0.041
R23809 vss.n22648 vss.n22647 0.041
R23810 vss.n22634 vss.n22633 0.041
R23811 vss.n22620 vss.n22619 0.041
R23812 vss.n22606 vss.n22605 0.041
R23813 vss.n22592 vss.n22591 0.041
R23814 vss.n22588 vss.n22587 0.041
R23815 vss.n22574 vss.n22573 0.041
R23816 vss.n22560 vss.n22559 0.041
R23817 vss.n22546 vss.n22545 0.041
R23818 vss.n22532 vss.n22531 0.041
R23819 vss.n22518 vss.n22517 0.041
R23820 vss.n22504 vss.n22503 0.041
R23821 vss.n22468 vss.n22467 0.041
R23822 vss.n22454 vss.n22453 0.041
R23823 vss.n22440 vss.n22439 0.041
R23824 vss.n22426 vss.n22425 0.041
R23825 vss.n22412 vss.n22411 0.041
R23826 vss.n22398 vss.n22397 0.041
R23827 vss.n22384 vss.n22383 0.041
R23828 vss.n22380 vss.n22379 0.041
R23829 vss.n22366 vss.n22365 0.041
R23830 vss.n22352 vss.n22351 0.041
R23831 vss.n22338 vss.n22337 0.041
R23832 vss.n22324 vss.n22323 0.041
R23833 vss.n22310 vss.n22309 0.041
R23834 vss.n22296 vss.n22295 0.041
R23835 vss.n22260 vss.n22259 0.041
R23836 vss.n22246 vss.n22245 0.041
R23837 vss.n22232 vss.n22231 0.041
R23838 vss.n22218 vss.n22217 0.041
R23839 vss.n22204 vss.n22203 0.041
R23840 vss.n22190 vss.n22189 0.041
R23841 vss.n22176 vss.n22175 0.041
R23842 vss.n22172 vss.n22171 0.041
R23843 vss.n22158 vss.n22157 0.041
R23844 vss.n22144 vss.n22143 0.041
R23845 vss.n22130 vss.n22129 0.041
R23846 vss.n22116 vss.n22115 0.041
R23847 vss.n22102 vss.n22101 0.041
R23848 vss.n22088 vss.n22087 0.041
R23849 vss.n22809 vss.n1430 0.041
R23850 vss.n9183 vss.n9182 0.041
R23851 vss.n9180 vss.n9179 0.041
R23852 vss.n9181 vss.n9180 0.041
R23853 vss.n9187 vss.n9186 0.041
R23854 vss.n9188 vss.n9187 0.041
R23855 vss.n9189 vss.n9188 0.041
R23856 vss.n9190 vss.n9189 0.041
R23857 vss.n20401 vss.n17554 0.04
R23858 vss.n7011 vss.n4164 0.04
R23859 vss.n20398 vss.n17558 0.04
R23860 vss.n20388 vss.n20387 0.04
R23861 vss.n20404 vss.n20403 0.04
R23862 vss.n17549 ldomc_0.otaldom_0.nmosbn2m_0.vss 0.04
R23863 vss.n9167 vss.n9166 0.04
R23864 vss.n9165 vss.n9164 0.04
R23865 vss.n10417 vss.n10397 0.04
R23866 vss.n10417 vss.n10415 0.04
R23867 vss.n10430 vss.n10427 0.04
R23868 vss.n10430 vss.n10428 0.04
R23869 vss.n10447 vss.n10446 0.04
R23870 vss.n7008 vss.n4168 0.04
R23871 vss.n6998 vss.n6997 0.04
R23872 vss.n7014 vss.n7013 0.04
R23873 vss.n4159 bandgapmd_0.otam_1.nmosbn2m_0.vss 0.04
R23874 vss.n1876 vss.n1875 0.04
R23875 vss.n2002 vss.n2000 0.04
R23876 vss.n2121 vss.n2120 0.04
R23877 vss.n2244 vss.n2240 0.04
R23878 vss.n2246 vss.n2244 0.04
R23879 vss.n2365 vss.n2364 0.04
R23880 vss.n2488 vss.n2484 0.04
R23881 vss.n2490 vss.n2488 0.04
R23882 vss.n2733 vss.n2729 0.04
R23883 vss.n2735 vss.n2733 0.04
R23884 vss.n2848 vss.n2847 0.04
R23885 vss.n2971 vss.n2967 0.04
R23886 vss.n2973 vss.n2971 0.04
R23887 vss.n3092 vss.n3091 0.04
R23888 vss.n3215 vss.n3211 0.04
R23889 vss.n3337 vss.n3336 0.04
R23890 vss.n15216 ldomc_0.vdm_0.vss 0.04
R23891 vss.n337 vss.n336 0.04
R23892 vss.n463 vss.n461 0.04
R23893 vss.n582 vss.n581 0.04
R23894 vss.n705 vss.n701 0.04
R23895 vss.n707 vss.n705 0.04
R23896 vss.n826 vss.n825 0.04
R23897 vss.n949 vss.n945 0.04
R23898 vss.n951 vss.n949 0.04
R23899 vss.n1194 vss.n1190 0.04
R23900 vss.n1196 vss.n1194 0.04
R23901 vss.n23409 vss.n23408 0.04
R23902 vss.n23291 vss.n23289 0.04
R23903 vss.n23289 vss.n23285 0.04
R23904 vss.n23166 vss.n23165 0.04
R23905 vss.n23047 vss.n23045 0.04
R23906 vss.n22921 vss.n22920 0.04
R23907 vss.n21901 vss.n21896 0.04
R23908 vss.n3850 vss.n3845 0.04
R23909 vss.n21978 vss.n21977 0.04
R23910 vss.n3927 vss.n3926 0.04
R23911 vss.n8945 vss.n8944 0.04
R23912 vss.n9666 vss.n9665 0.04
R23913 vss.n8951 vss.n8950 0.039
R23914 vss.n10415 vss.n10413 0.039
R23915 vss.n20362 vss.n20361 0.039
R23916 vss.n20371 vss.n17580 0.039
R23917 vss.n20381 vss.n20380 0.039
R23918 vss.n14824 vss.n14823 0.039
R23919 vss.n14826 vss.n14824 0.039
R23920 vss.n14827 vss.n14826 0.039
R23921 vss.n14850 vss.n14842 0.039
R23922 vss.n14851 vss.n14850 0.039
R23923 vss.n6972 vss.n6971 0.039
R23924 vss.n6981 vss.n4190 0.039
R23925 vss.n6991 vss.n6990 0.039
R23926 vss.n9667 vss.n9666 0.039
R23927 vss.n11097 vss.n11086 0.039
R23928 vss.n20387 vss.n17558 0.038
R23929 vss.n12897 vss.n12896 0.038
R23930 vss.n6997 vss.n4168 0.038
R23931 vss.n3451 vss.n3450 0.038
R23932 vss.n1426 vss.n1425 0.038
R23933 vss.n10318 vss.n10317 0.037
R23934 vss.n10385 vss.n10364 0.037
R23935 vss.n10385 vss.n10384 0.037
R23936 vss.n9073 vss.n9072 0.037
R23937 vss.n9075 vss.n9073 0.037
R23938 vss.n9148 vss.n9147 0.037
R23939 vss.n9150 vss.n9148 0.037
R23940 vss.n15064 vss.n15063 0.037
R23941 vss.n20394 vss.n20393 0.037
R23942 vss.n14842 vss.n14841 0.037
R23943 vss.n14852 vss.n14851 0.037
R23944 vss.n7004 vss.n7003 0.037
R23945 vss.n10338 vss.n10337 0.037
R23946 vss.n9121 vss.n9120 0.037
R23947 vss.n9123 vss.n9121 0.037
R23948 vss.n9042 vss.n9041 0.036
R23949 vss.n9044 vss.n9042 0.036
R23950 vss.n12903 vss.n12902 0.036
R23951 vss.n12876 vss.n12875 0.036
R23952 vss.n7848 vss.n7847 0.036
R23953 vss.n10274 vss.n10273 0.035
R23954 vss.n9013 vss.n9011 0.035
R23955 vss.n10349 vss.n10348 0.035
R23956 vss.n10350 vss.n10349 0.035
R23957 vss.n14867 vss.n14866 0.035
R23958 vss.n10262 vss.n10255 0.035
R23959 vss.n19624 vss.n19623 0.034
R23960 vss.n6234 vss.n6233 0.034
R23961 vss.n20385 vss.n17558 0.034
R23962 vss.n6995 vss.n4168 0.034
R23963 vss.n17564 vss.n17559 0.034
R23964 vss.n21874 vss.n21867 0.034
R23965 vss.n21930 vss.n21927 0.034
R23966 vss.n21957 vss.n21954 0.034
R23967 vss.n21626 vss.n21623 0.034
R23968 vss.n12861 vss.n12860 0.034
R23969 vss.n3823 vss.n3816 0.034
R23970 vss.n3879 vss.n3876 0.034
R23971 vss.n3906 vss.n3903 0.034
R23972 vss.n4174 vss.n4169 0.034
R23973 vss.n3575 vss.n3572 0.034
R23974 vss.n21896 vss.n21895 0.034
R23975 vss.n3845 vss.n3844 0.034
R23976 vss.n22056 vss.n22053 0.034
R23977 vss.n4005 vss.n4002 0.034
R23978 vss.n20305 vss.n20303 0.033
R23979 vss.n6915 vss.n6913 0.033
R23980 vss.n20393 vss.n17561 0.033
R23981 vss.n20505 vss.n20504 0.033
R23982 vss.n20768 vss.n20764 0.033
R23983 vss.n20769 vss.n20768 0.033
R23984 vss.n21756 vss.n21697 0.033
R23985 vss.n14898 vss.n14897 0.033
R23986 vss.n3705 vss.n3646 0.033
R23987 vss.n7003 vss.n4171 0.033
R23988 vss.n7115 vss.n7114 0.033
R23989 vss.n7378 vss.n7374 0.033
R23990 vss.n7379 vss.n7378 0.033
R23991 vss.n15125 bandgapmd_0.vss 0.033
R23992 vss.n20383 vss.n17558 0.033
R23993 vss.n6993 vss.n4168 0.033
R23994 vss.n10413 vss.n10412 0.033
R23995 vss.n9011 vss.n9010 0.033
R23996 vss.n10347 vss.n10342 0.032
R23997 vss.n20892 vss.n20860 0.032
R23998 vss.n12824 vss.n12823 0.032
R23999 vss.n12534 vss.n12533 0.032
R24000 vss.n12149 vss.n12148 0.032
R24001 vss.n12846 vss.n12845 0.032
R24002 vss.n7502 vss.n7470 0.032
R24003 vss.n13645 vss.n13644 0.031
R24004 vss.n10656 vss.n10655 0.031
R24005 vss.n11469 vss.n11468 0.031
R24006 vss.n13677 vss.n13676 0.031
R24007 vss.n13136 vss.n13135 0.031
R24008 vss.n13127 vss.n13126 0.031
R24009 vss.n10664 vss.n10663 0.031
R24010 vss.n11461 vss.n11460 0.031
R24011 vss.n21711 vss.n21710 0.03
R24012 vss.n3660 vss.n3659 0.03
R24013 vss.n10228 vss.n10226 0.03
R24014 vss.n21967 vss.n21966 0.03
R24015 vss.n10282 vss.n10281 0.03
R24016 vss.n10382 vss.n10381 0.03
R24017 vss.n12777 vss.n12776 0.03
R24018 vss.n14883 vss.n14882 0.03
R24019 vss.n3916 vss.n3915 0.03
R24020 vss.n1814 vss.n1812 0.03
R24021 vss.n1829 vss.n1827 0.03
R24022 vss.n1844 vss.n1842 0.03
R24023 vss.n1859 vss.n1857 0.03
R24024 vss.n1874 vss.n1872 0.03
R24025 vss.n1907 vss.n1895 0.03
R24026 vss.n1923 vss.n1911 0.03
R24027 vss.n1939 vss.n1927 0.03
R24028 vss.n1955 vss.n1943 0.03
R24029 vss.n1971 vss.n1959 0.03
R24030 vss.n1991 vss.n1975 0.03
R24031 vss.n2022 vss.n2020 0.03
R24032 vss.n2038 vss.n2036 0.03
R24033 vss.n2054 vss.n2052 0.03
R24034 vss.n2070 vss.n2068 0.03
R24035 vss.n2086 vss.n2084 0.03
R24036 vss.n2119 vss.n2117 0.03
R24037 vss.n2135 vss.n2123 0.03
R24038 vss.n2151 vss.n2139 0.03
R24039 vss.n2167 vss.n2155 0.03
R24040 vss.n2183 vss.n2171 0.03
R24041 vss.n2216 vss.n2204 0.03
R24042 vss.n2236 vss.n2220 0.03
R24043 vss.n2266 vss.n2264 0.03
R24044 vss.n2282 vss.n2280 0.03
R24045 vss.n2299 vss.n2296 0.03
R24046 vss.n2315 vss.n2313 0.03
R24047 vss.n2331 vss.n2329 0.03
R24048 vss.n2347 vss.n2345 0.03
R24049 vss.n2363 vss.n2361 0.03
R24050 vss.n2379 vss.n2367 0.03
R24051 vss.n2395 vss.n2383 0.03
R24052 vss.n2412 vss.n2400 0.03
R24053 vss.n2428 vss.n2416 0.03
R24054 vss.n2444 vss.n2432 0.03
R24055 vss.n2460 vss.n2448 0.03
R24056 vss.n2480 vss.n2464 0.03
R24057 vss.n2527 vss.n2525 0.03
R24058 vss.n2543 vss.n2541 0.03
R24059 vss.n2559 vss.n2557 0.03
R24060 vss.n2575 vss.n2573 0.03
R24061 vss.n2591 vss.n2589 0.03
R24062 vss.n2607 vss.n2605 0.03
R24063 vss.n2624 vss.n2612 0.03
R24064 vss.n2640 vss.n2628 0.03
R24065 vss.n2656 vss.n2644 0.03
R24066 vss.n2672 vss.n2660 0.03
R24067 vss.n2688 vss.n2676 0.03
R24068 vss.n2704 vss.n2692 0.03
R24069 vss.n2755 vss.n2753 0.03
R24070 vss.n2771 vss.n2769 0.03
R24071 vss.n2787 vss.n2785 0.03
R24072 vss.n2803 vss.n2801 0.03
R24073 vss.n2818 vss.n2816 0.03
R24074 vss.n2832 vss.n2831 0.03
R24075 vss.n2862 vss.n2850 0.03
R24076 vss.n2878 vss.n2866 0.03
R24077 vss.n2894 vss.n2882 0.03
R24078 vss.n2910 vss.n2898 0.03
R24079 vss.n2927 vss.n2915 0.03
R24080 vss.n2943 vss.n2931 0.03
R24081 vss.n2963 vss.n2947 0.03
R24082 vss.n2993 vss.n2991 0.03
R24083 vss.n3009 vss.n3007 0.03
R24084 vss.n3026 vss.n3024 0.03
R24085 vss.n3042 vss.n3040 0.03
R24086 vss.n3058 vss.n3056 0.03
R24087 vss.n3074 vss.n3072 0.03
R24088 vss.n3090 vss.n3088 0.03
R24089 vss.n3106 vss.n3094 0.03
R24090 vss.n3139 vss.n3127 0.03
R24091 vss.n3155 vss.n3143 0.03
R24092 vss.n3171 vss.n3159 0.03
R24093 vss.n3187 vss.n3175 0.03
R24094 vss.n3207 vss.n3191 0.03
R24095 vss.n3238 vss.n3236 0.03
R24096 vss.n3254 vss.n3252 0.03
R24097 vss.n3270 vss.n3268 0.03
R24098 vss.n3286 vss.n3284 0.03
R24099 vss.n3302 vss.n3300 0.03
R24100 vss.n3318 vss.n3316 0.03
R24101 vss.n3350 vss.n3339 0.03
R24102 vss.n3365 vss.n3354 0.03
R24103 vss.n3380 vss.n3369 0.03
R24104 vss.n3395 vss.n3384 0.03
R24105 vss.n3410 vss.n3399 0.03
R24106 vss.n275 vss.n273 0.03
R24107 vss.n290 vss.n288 0.03
R24108 vss.n305 vss.n303 0.03
R24109 vss.n320 vss.n318 0.03
R24110 vss.n335 vss.n333 0.03
R24111 vss.n368 vss.n356 0.03
R24112 vss.n384 vss.n372 0.03
R24113 vss.n400 vss.n388 0.03
R24114 vss.n416 vss.n404 0.03
R24115 vss.n432 vss.n420 0.03
R24116 vss.n452 vss.n436 0.03
R24117 vss.n483 vss.n481 0.03
R24118 vss.n499 vss.n497 0.03
R24119 vss.n515 vss.n513 0.03
R24120 vss.n531 vss.n529 0.03
R24121 vss.n547 vss.n545 0.03
R24122 vss.n580 vss.n578 0.03
R24123 vss.n596 vss.n584 0.03
R24124 vss.n612 vss.n600 0.03
R24125 vss.n628 vss.n616 0.03
R24126 vss.n644 vss.n632 0.03
R24127 vss.n677 vss.n665 0.03
R24128 vss.n697 vss.n681 0.03
R24129 vss.n727 vss.n725 0.03
R24130 vss.n743 vss.n741 0.03
R24131 vss.n760 vss.n757 0.03
R24132 vss.n776 vss.n774 0.03
R24133 vss.n792 vss.n790 0.03
R24134 vss.n808 vss.n806 0.03
R24135 vss.n824 vss.n822 0.03
R24136 vss.n840 vss.n828 0.03
R24137 vss.n856 vss.n844 0.03
R24138 vss.n873 vss.n861 0.03
R24139 vss.n889 vss.n877 0.03
R24140 vss.n905 vss.n893 0.03
R24141 vss.n921 vss.n909 0.03
R24142 vss.n941 vss.n925 0.03
R24143 vss.n988 vss.n986 0.03
R24144 vss.n1004 vss.n1002 0.03
R24145 vss.n1020 vss.n1018 0.03
R24146 vss.n1036 vss.n1034 0.03
R24147 vss.n1052 vss.n1050 0.03
R24148 vss.n1068 vss.n1066 0.03
R24149 vss.n1085 vss.n1073 0.03
R24150 vss.n1101 vss.n1089 0.03
R24151 vss.n1117 vss.n1105 0.03
R24152 vss.n1133 vss.n1121 0.03
R24153 vss.n1149 vss.n1137 0.03
R24154 vss.n1165 vss.n1153 0.03
R24155 vss.n1216 vss.n1214 0.03
R24156 vss.n1232 vss.n1230 0.03
R24157 vss.n1248 vss.n1246 0.03
R24158 vss.n1264 vss.n1262 0.03
R24159 vss.n1280 vss.n1278 0.03
R24160 vss.n1297 vss.n1295 0.03
R24161 vss.n23407 vss.n23405 0.03
R24162 vss.n23391 vss.n23389 0.03
R24163 vss.n23375 vss.n23373 0.03
R24164 vss.n23359 vss.n23357 0.03
R24165 vss.n23343 vss.n23341 0.03
R24166 vss.n23327 vss.n23325 0.03
R24167 vss.n23311 vss.n23309 0.03
R24168 vss.n23281 vss.n23265 0.03
R24169 vss.n23261 vss.n23249 0.03
R24170 vss.n23244 vss.n23232 0.03
R24171 vss.n23228 vss.n23216 0.03
R24172 vss.n23212 vss.n23200 0.03
R24173 vss.n23196 vss.n23184 0.03
R24174 vss.n23180 vss.n23168 0.03
R24175 vss.n23164 vss.n23162 0.03
R24176 vss.n23131 vss.n23129 0.03
R24177 vss.n23115 vss.n23113 0.03
R24178 vss.n23099 vss.n23097 0.03
R24179 vss.n23083 vss.n23081 0.03
R24180 vss.n23067 vss.n23065 0.03
R24181 vss.n23036 vss.n23020 0.03
R24182 vss.n23016 vss.n23004 0.03
R24183 vss.n23000 vss.n22988 0.03
R24184 vss.n22984 vss.n22972 0.03
R24185 vss.n22968 vss.n22956 0.03
R24186 vss.n22952 vss.n22940 0.03
R24187 vss.n22919 vss.n22917 0.03
R24188 vss.n22904 vss.n22902 0.03
R24189 vss.n22889 vss.n22887 0.03
R24190 vss.n22874 vss.n22872 0.03
R24191 vss.n22859 vss.n22857 0.03
R24192 vss.n17555 vss.n17550 0.03
R24193 vss.n4165 vss.n4160 0.03
R24194 vss.n20398 vss.n20397 0.029
R24195 vss.n20394 vss.n17560 0.029
R24196 vss.n17571 vss.n17568 0.029
R24197 vss.n21635 vss.n21629 0.029
R24198 vss.n14869 vss.n14868 0.029
R24199 vss.n12737 vss.n12736 0.029
R24200 vss.n7008 vss.n7007 0.029
R24201 vss.n7004 vss.n4170 0.029
R24202 vss.n4181 vss.n4178 0.029
R24203 vss.n3584 vss.n3578 0.029
R24204 vss.n2188 vss.n2187 0.029
R24205 vss.n16252 vss.n16240 0.029
R24206 vss.n649 vss.n648 0.029
R24207 vss.n20402 vss.n17555 0.029
R24208 vss.n7012 vss.n4165 0.029
R24209 vss.n21885 vss.n21878 0.028
R24210 vss.n21937 vss.n21934 0.028
R24211 vss.n21964 vss.n21961 0.028
R24212 vss.n9195 vss.t218 0.028
R24213 vss.n9194 vss.t219 0.028
R24214 vss.n10411 vss.n10409 0.028
R24215 vss.n12800 vss.n12799 0.028
R24216 vss.n12544 vss.n12543 0.028
R24217 vss.n3834 vss.n3827 0.028
R24218 vss.n3886 vss.n3883 0.028
R24219 vss.n3913 vss.n3910 0.028
R24220 vss.n15123 vss.n8920 0.028
R24221 vss.n15209 vss.n3414 0.028
R24222 vss.n22758 vss.n22757 0.028
R24223 vss.n22844 vss.n22842 0.028
R24224 vss.n21799 vss.n21645 0.028
R24225 vss.n3748 vss.n3594 0.028
R24226 vss.n15062 vss.n12735 0.027
R24227 vss.n21636 vss.n21635 0.027
R24228 vss.n3585 vss.n3584 0.027
R24229 vss.n10305 vss.n10304 0.027
R24230 vss.n20389 vss.n17558 0.027
R24231 vss.n6999 vss.n4168 0.027
R24232 vss.n21905 vss.n21856 0.027
R24233 vss.n21940 vss.n21939 0.027
R24234 vss.n12778 vss.n12777 0.027
R24235 vss.n10725 vss.n10724 0.027
R24236 vss.n13111 vss.n12994 0.027
R24237 vss.n14884 vss.n14883 0.027
R24238 vss.n3854 vss.n3805 0.027
R24239 vss.n3889 vss.n3888 0.027
R24240 vss.n2709 vss.n2708 0.027
R24241 vss.n1170 vss.n1169 0.027
R24242 vss.n10384 vss.n10383 0.026
R24243 vss.n15061 vss.n15060 0.026
R24244 vss.n12823 vss.n12822 0.026
R24245 vss.n12148 vss.n12147 0.026
R24246 vss.n12847 vss.n12846 0.026
R24247 vss.n8983 vss.n8981 0.026
R24248 vss.n8970 vss.n8969 0.026
R24249 vss.n17569 vss.n17568 0.025
R24250 vss.n20593 vss.n20591 0.025
R24251 vss.n20608 vss.n20606 0.025
R24252 vss.n20623 vss.n20621 0.025
R24253 vss.n20638 vss.n20636 0.025
R24254 vss.n20653 vss.n20651 0.025
R24255 vss.n20684 vss.n20673 0.025
R24256 vss.n20699 vss.n20688 0.025
R24257 vss.n20714 vss.n20703 0.025
R24258 vss.n20729 vss.n20718 0.025
R24259 vss.n20744 vss.n20733 0.025
R24260 vss.n20785 vss.n20783 0.025
R24261 vss.n20816 vss.n20814 0.025
R24262 vss.n20831 vss.n20829 0.025
R24263 vss.n21878 vss.n21876 0.025
R24264 vss.n21934 vss.n21932 0.025
R24265 vss.n21961 vss.n21959 0.025
R24266 vss.n21627 vss.n21626 0.025
R24267 vss.n10243 vss.n10242 0.025
R24268 vss.n10244 vss.n10243 0.025
R24269 vss.n10247 vss.n10246 0.025
R24270 vss.n10268 vss.n10267 0.025
R24271 vss.n10271 vss.n10270 0.025
R24272 vss.n10287 vss.n10286 0.025
R24273 vss.n10288 vss.n10287 0.025
R24274 vss.n10291 vss.n10290 0.025
R24275 vss.n10310 vss.n10309 0.025
R24276 vss.n10311 vss.n10310 0.025
R24277 vss.n10314 vss.n10313 0.025
R24278 vss.n10328 vss.n10327 0.025
R24279 vss.n10329 vss.n10328 0.025
R24280 vss.n10332 vss.n10331 0.025
R24281 vss.n10370 vss.n10369 0.025
R24282 vss.n10371 vss.n10370 0.025
R24283 vss.n10374 vss.n10373 0.025
R24284 vss.n10402 vss.n10401 0.025
R24285 vss.n10403 vss.n10402 0.025
R24286 vss.n10406 vss.n10405 0.025
R24287 vss.n10436 vss.n10435 0.025
R24288 vss.n10437 vss.n10436 0.025
R24289 vss.n10440 vss.n10439 0.025
R24290 vss.n10452 vss.n10432 0.025
R24291 vss.n8942 vss.n8939 0.025
R24292 vss.n8939 vss.n8938 0.025
R24293 vss.n8936 vss.n8935 0.025
R24294 vss.n8960 vss.n8957 0.025
R24295 vss.n8957 vss.n8956 0.025
R24296 vss.n8954 vss.n8953 0.025
R24297 vss.n8992 vss.n8991 0.025
R24298 vss.n8993 vss.n8992 0.025
R24299 vss.n8996 vss.n8995 0.025
R24300 vss.n9022 vss.n9021 0.025
R24301 vss.n9023 vss.n9022 0.025
R24302 vss.n9026 vss.n9025 0.025
R24303 vss.n9053 vss.n9052 0.025
R24304 vss.n9054 vss.n9053 0.025
R24305 vss.n9057 vss.n9056 0.025
R24306 vss.n9084 vss.n9083 0.025
R24307 vss.n9085 vss.n9084 0.025
R24308 vss.n9088 vss.n9087 0.025
R24309 vss.n9103 vss.n9102 0.025
R24310 vss.n9104 vss.n9103 0.025
R24311 vss.n9107 vss.n9106 0.025
R24312 vss.n9133 vss.n9132 0.025
R24313 vss.n9134 vss.n9133 0.025
R24314 vss.n9137 vss.n9136 0.025
R24315 vss.n11407 vss.n11405 0.025
R24316 vss.n14908 vss.n14898 0.025
R24317 vss.n3827 vss.n3825 0.025
R24318 vss.n3883 vss.n3881 0.025
R24319 vss.n3910 vss.n3908 0.025
R24320 vss.n4179 vss.n4178 0.025
R24321 vss.n7203 vss.n7201 0.025
R24322 vss.n7218 vss.n7216 0.025
R24323 vss.n7233 vss.n7231 0.025
R24324 vss.n7248 vss.n7246 0.025
R24325 vss.n7263 vss.n7261 0.025
R24326 vss.n7294 vss.n7283 0.025
R24327 vss.n7309 vss.n7298 0.025
R24328 vss.n7324 vss.n7313 0.025
R24329 vss.n7339 vss.n7328 0.025
R24330 vss.n7354 vss.n7343 0.025
R24331 vss.n7395 vss.n7393 0.025
R24332 vss.n7426 vss.n7424 0.025
R24333 vss.n7441 vss.n7439 0.025
R24334 vss.n3576 vss.n3575 0.025
R24335 vss.n3439 vss.n3437 0.025
R24336 vss.n1414 vss.n1412 0.025
R24337 vss.n19616 vss.n19592 0.024
R24338 vss.n20366 vss.n20365 0.024
R24339 vss.n20396 vss.n20395 0.024
R24340 vss.n21755 vss.n21699 0.024
R24341 vss.n21626 vss.n21625 0.024
R24342 vss.n8968 vss.n8967 0.024
R24343 vss.n12906 vss.n12904 0.024
R24344 vss.n12493 vss.n12491 0.024
R24345 vss.n12863 vss.n12861 0.024
R24346 vss.n12738 vss.n12737 0.024
R24347 vss.n12739 vss.n12738 0.024
R24348 vss.n12740 vss.n12739 0.024
R24349 vss.n12741 vss.n12740 0.024
R24350 vss.n12742 vss.n12741 0.024
R24351 vss.n12743 vss.n12742 0.024
R24352 vss.n12744 vss.n12743 0.024
R24353 vss.n12745 vss.n12744 0.024
R24354 vss.n12746 vss.n12745 0.024
R24355 vss.n12747 vss.n12746 0.024
R24356 vss.n12748 vss.n12747 0.024
R24357 vss.n12749 vss.n12748 0.024
R24358 vss.n12750 vss.n12749 0.024
R24359 vss.n12751 vss.n12750 0.024
R24360 vss.n12752 vss.n12751 0.024
R24361 vss.n12753 vss.n12752 0.024
R24362 vss.n12754 vss.n12753 0.024
R24363 vss.n12755 vss.n12754 0.024
R24364 vss.n12756 vss.n12755 0.024
R24365 vss.n12757 vss.n12756 0.024
R24366 vss.n12758 vss.n12757 0.024
R24367 vss.n12759 vss.n12758 0.024
R24368 vss.n12760 vss.n12759 0.024
R24369 vss.n12762 vss.n12761 0.024
R24370 vss.n12763 vss.n12762 0.024
R24371 vss.n12765 vss.n12764 0.024
R24372 vss.n12766 vss.n12765 0.024
R24373 vss.n12767 vss.n12766 0.024
R24374 vss.n12768 vss.n12767 0.024
R24375 vss.n12769 vss.n12768 0.024
R24376 vss.n15096 vss.n15095 0.024
R24377 vss.n15095 vss.n15094 0.024
R24378 vss.n15094 vss.n15093 0.024
R24379 vss.n15093 vss.n15092 0.024
R24380 vss.n15092 vss.n15091 0.024
R24381 vss.n15091 vss.n15090 0.024
R24382 vss.n15090 vss.n15089 0.024
R24383 vss.n15089 vss.n15088 0.024
R24384 vss.n15088 vss.n15087 0.024
R24385 vss.n15087 vss.n15086 0.024
R24386 vss.n15086 vss.n15085 0.024
R24387 vss.n15085 vss.n15084 0.024
R24388 vss.n15084 vss.n15083 0.024
R24389 vss.n15083 vss.n15082 0.024
R24390 vss.n15082 vss.n15081 0.024
R24391 vss.n15081 vss.n15080 0.024
R24392 vss.n15080 vss.n15079 0.024
R24393 vss.n15079 vss.n15078 0.024
R24394 vss.n15078 vss.n15077 0.024
R24395 vss.n15077 vss.n15076 0.024
R24396 vss.n15076 vss.n15075 0.024
R24397 vss.n15075 vss.n15074 0.024
R24398 vss.n15073 vss.n15072 0.024
R24399 vss.n15072 vss.n15071 0.024
R24400 vss.n15070 vss.n15069 0.024
R24401 vss.n15069 vss.n15068 0.024
R24402 vss.n15068 vss.n15067 0.024
R24403 vss.n15067 vss.n15066 0.024
R24404 vss.n15066 vss.n15065 0.024
R24405 vss.n15065 vss.n15064 0.024
R24406 vss.n3704 vss.n3648 0.024
R24407 vss.n6226 vss.n6202 0.024
R24408 vss.n6976 vss.n6975 0.024
R24409 vss.n7006 vss.n7005 0.024
R24410 vss.n3575 vss.n3574 0.024
R24411 vss.n1799 vss.n1797 0.024
R24412 vss.n3123 vss.n3111 0.024
R24413 vss.n3333 vss.n3332 0.024
R24414 vss.n260 vss.n258 0.024
R24415 vss.n23146 vss.n23145 0.024
R24416 vss.n22936 vss.n22924 0.024
R24417 vss.n22069 vss.n22068 0.024
R24418 vss.n9072 vss.n9071 0.023
R24419 vss.n20400 vss.n20399 0.023
R24420 vss.n20845 vss.n20844 0.023
R24421 vss.n9156 vss.n9155 0.023
R24422 vss.n12301 vss.n10792 0.023
R24423 vss.n12301 vss.n12300 0.023
R24424 vss.n14700 vss.n13420 0.023
R24425 vss.n14700 vss.n13499 0.023
R24426 vss.n14975 vss.n12953 0.023
R24427 vss.n14975 vss.n13183 0.023
R24428 vss.n12710 vss.n12355 0.023
R24429 vss.n12710 vss.n12393 0.023
R24430 vss.n14078 vss.n13798 0.023
R24431 vss.n14078 vss.n13818 0.023
R24432 vss.n11832 vss.n11524 0.023
R24433 vss.n11832 vss.n11554 0.023
R24434 vss.n14837 vss.n14827 0.023
R24435 vss.n14866 vss.n14865 0.023
R24436 vss.n7010 vss.n7009 0.023
R24437 vss.n7455 vss.n7454 0.023
R24438 vss.n8215 vss.n8214 0.023
R24439 vss.n1765 vss.n1761 0.023
R24440 vss.n1766 vss.n1765 0.023
R24441 vss.n2000 vss.n1996 0.023
R24442 vss.n2511 vss.n2509 0.023
R24443 vss.n3216 vss.n3215 0.023
R24444 vss.n16766 vss.n16756 0.023
R24445 vss.n16778 vss.n16768 0.023
R24446 vss.n16797 vss.n16796 0.023
R24447 vss.n16808 vss.n16807 0.023
R24448 vss.n16822 vss.n16821 0.023
R24449 vss.n16836 vss.n16835 0.023
R24450 vss.n226 vss.n222 0.023
R24451 vss.n227 vss.n226 0.023
R24452 vss.n461 vss.n457 0.023
R24453 vss.n972 vss.n970 0.023
R24454 vss.n23045 vss.n23041 0.023
R24455 vss.n20376 vss.n20375 0.022
R24456 vss.n21760 vss.n21698 0.022
R24457 vss.n22086 vss.n22085 0.022
R24458 vss.n12902 vss.n12901 0.022
R24459 vss.n12636 vss.n12633 0.022
R24460 vss.n10725 vss.n10570 0.022
R24461 vss.n13111 vss.n13013 0.022
R24462 vss.n12878 vss.n12876 0.022
R24463 vss.n3709 vss.n3647 0.022
R24464 vss.n6986 vss.n6985 0.022
R24465 vss.n8249 vss.n8248 0.022
R24466 vss.n2846 bandgapmd_0.otam_1.pdiffaloadm_0.vss 0.022
R24467 vss.n3449 vss.n3446 0.022
R24468 ldomc_0.otaldom_0.pdiffaloadm_0.vss vss.n23411 0.022
R24469 vss.n1424 vss.n1421 0.022
R24470 vss.n10442 vss.n10441 0.022
R24471 vss.n21635 vss.n21616 0.021
R24472 vss.n3584 vss.n3565 0.021
R24473 vss.n10351 vss.n10350 0.021
R24474 vss.n10304 vss.n10303 0.021
R24475 vss.n10363 vss.n10362 0.021
R24476 vss.n19617 vss.n19616 0.021
R24477 vss.n20403 vss.n17553 0.021
R24478 vss.n19622 vss.n19588 0.021
R24479 vss.n20402 vss.n20400 0.021
R24480 vss.n20656 vss.n20655 0.021
R24481 vss.n21800 vss.n21642 0.021
R24482 vss.n10236 vss.n10233 0.021
R24483 vss.n10353 vss.n10352 0.021
R24484 vss.n12491 vss.n12490 0.021
R24485 vss.n12543 vss.n12542 0.021
R24486 vss.n11099 vss.n11097 0.021
R24487 vss.n14266 vss.n14264 0.021
R24488 vss.n12898 vss.n12897 0.021
R24489 vss.n3749 vss.n3591 0.021
R24490 vss.n6227 vss.n6226 0.021
R24491 vss.n7013 vss.n4163 0.021
R24492 vss.n6232 vss.n6198 0.021
R24493 vss.n7012 vss.n7010 0.021
R24494 vss.n7266 vss.n7265 0.021
R24495 vss.n1891 vss.n1879 0.021
R24496 vss.n2101 vss.n2100 0.021
R24497 vss.n2609 vss.n2608 0.021
R24498 vss.n15549 vss.n15548 0.021
R24499 vss.n15783 vss.n15782 0.021
R24500 vss.n15306 vss.n15305 0.021
R24501 vss.n15308 vss.n15307 0.021
R24502 vss.n15325 vss.n15324 0.021
R24503 vss.n15328 vss.n15326 0.021
R24504 vss.n15342 vss.n15340 0.021
R24505 vss.n15356 vss.n15354 0.021
R24506 vss.n16075 vss.n16074 0.021
R24507 vss.n16496 vss.n16495 0.021
R24508 vss.n17029 vss.n17017 0.021
R24509 vss.n17265 vss.n17253 0.021
R24510 vss.n352 vss.n340 0.021
R24511 vss.n562 vss.n561 0.021
R24512 vss.n1070 vss.n1069 0.021
R24513 vss.n21656 vss.n21651 0.021
R24514 vss.n3605 vss.n3600 0.021
R24515 vss.n20378 vss.n20377 0.021
R24516 vss.n6988 vss.n6987 0.021
R24517 vss.n9036 vss.n9035 0.02
R24518 vss.n9713 vss.n9712 0.02
R24519 vss.n17560 vss.n17558 0.02
R24520 vss.n19615 vss.n19588 0.02
R24521 vss.n15061 vss.n12769 0.02
R24522 vss.n4170 vss.n4168 0.02
R24523 vss.n6225 vss.n6198 0.02
R24524 vss.n15415 vss.n15413 0.02
R24525 vss.n15436 vss.n15434 0.02
R24526 vss.n15651 vss.n15649 0.02
R24527 vss.n15672 vss.n15670 0.02
R24528 vss.n15821 vss.n15819 0.02
R24529 vss.n15947 vss.n15938 0.02
R24530 vss.n15962 vss.n15961 0.02
R24531 vss.n16183 vss.n16174 0.02
R24532 vss.n16198 vss.n16197 0.02
R24533 vss.n16286 vss.n16284 0.02
R24534 vss.n16362 vss.n16360 0.02
R24535 vss.n16383 vss.n16381 0.02
R24536 vss.n16598 vss.n16596 0.02
R24537 vss.n16619 vss.n16617 0.02
R24538 vss.n16686 vss.n16685 0.02
R24539 vss.n16893 vss.n16892 0.02
R24540 vss.n16916 vss.n16915 0.02
R24541 vss.n9712 vss.n9709 0.02
R24542 vss.n21672 vss.n21669 0.019
R24543 vss.n3621 vss.n3618 0.019
R24544 vss.n20360 vss.n20359 0.019
R24545 vss.n21755 vss.n21754 0.019
R24546 vss.n21703 vss.n21702 0.019
R24547 vss.n13309 vss.n13308 0.019
R24548 vss.n14973 vss.n14968 0.019
R24549 vss.n14821 bandgapmd_0.pnp_groupm_0.vss 0.019
R24550 vss.n3704 vss.n3703 0.019
R24551 vss.n3652 vss.n3651 0.019
R24552 vss.n6970 vss.n6969 0.019
R24553 vss.n8216 vss.n8215 0.019
R24554 vss.n17129 vss.n17128 0.019
R24555 vss.n17152 vss.n17151 0.019
R24556 vss.n16254 vss.n16253 0.019
R24557 vss.n22842 vss 0.019
R24558 vss.n9184 vss.n9183 0.019
R24559 vss.n10221 vss.n10214 0.019
R24560 vss.n10214 vss.n10210 0.018
R24561 vss.n9709 vss.n9705 0.018
R24562 vss.n21632 vss.n21631 0.018
R24563 vss.n3581 vss.n3580 0.018
R24564 vss.n19613 vss.n17585 0.018
R24565 vss.n20749 vss.n20748 0.018
R24566 vss.n21867 vss.n21865 0.018
R24567 vss.n21927 vss.n21926 0.018
R24568 vss.n21760 vss.n21700 0.018
R24569 vss.n21615 vss.n21614 0.018
R24570 vss.n10224 vss.n10223 0.018
R24571 vss.n14093 vss.n14092 0.018
R24572 vss.n13758 vss.n13757 0.018
R24573 vss.n11495 vss.n11454 0.018
R24574 vss.n11849 vss.n11848 0.018
R24575 vss.n13451 vss.n13152 0.018
R24576 vss.n13110 vss.n13096 0.018
R24577 vss.n10686 vss.n10649 0.018
R24578 vss.n12334 vss.n12318 0.018
R24579 vss.n3816 vss.n3814 0.018
R24580 vss.n3876 vss.n3875 0.018
R24581 vss.n3709 vss.n3649 0.018
R24582 vss.n3564 vss.n3563 0.018
R24583 vss.n6223 vss.n4195 0.018
R24584 vss.n7359 vss.n7358 0.018
R24585 vss.n2610 vss.n2609 0.018
R24586 vss.n15215 vss.n15214 0.018
R24587 vss.n15532 vss.n15530 0.018
R24588 vss.n15563 vss.n15553 0.018
R24589 vss.n15768 vss.n15766 0.018
R24590 vss.n16059 vss.n16047 0.018
R24591 vss.n16089 vss.n16088 0.018
R24592 vss.n16479 vss.n16477 0.018
R24593 vss.n16510 vss.n16500 0.018
R24594 vss.n17013 vss.n17012 0.018
R24595 vss.n17043 vss.n17031 0.018
R24596 vss.n17249 vss.n17248 0.018
R24597 vss.n1071 vss.n1070 0.018
R24598 vss.n17569 vss.n17558 0.017
R24599 vss.n19614 vss.n17584 0.017
R24600 vss.n17535 vss.n17533 0.017
R24601 vss.n17545 vss.n17542 0.017
R24602 vss.n17490 vss.n17488 0.017
R24603 vss.n21941 vss.n21940 0.017
R24604 vss.n21970 vss.n21969 0.017
R24605 vss.n21760 vss.n21759 0.017
R24606 vss.n21653 vss.n21641 0.017
R24607 vss.n9176 vss.n9175 0.017
R24608 vss.n9192 vss.n9191 0.017
R24609 vss.n9178 vss.n9177 0.017
R24610 vss.n10411 vss.n10410 0.017
R24611 vss.n11219 vss.n11218 0.017
R24612 vss.n11101 vss.n11099 0.017
R24613 vss.n14268 vss.n14266 0.017
R24614 vss.n11134 vss.n11133 0.017
R24615 vss.n14443 vss.n14442 0.017
R24616 vss.n15007 vss.n15006 0.017
R24617 vss.n12895 vss.n12878 0.017
R24618 vss.n3890 vss.n3889 0.017
R24619 vss.n3919 vss.n3918 0.017
R24620 vss.n3709 vss.n3708 0.017
R24621 vss.n3602 vss.n3590 0.017
R24622 vss.n4179 vss.n4168 0.017
R24623 vss.n6224 vss.n4194 0.017
R24624 vss.n4145 vss.n4143 0.017
R24625 vss.n4155 vss.n4152 0.017
R24626 vss.n4100 vss.n4098 0.017
R24627 vss.n1708 vss.n1697 0.017
R24628 vss.n1723 vss.n1712 0.017
R24629 vss.n1738 vss.n1727 0.017
R24630 vss.n1782 vss.n1780 0.017
R24631 vss.n15401 vss.n15399 0.017
R24632 vss.n15450 vss.n15448 0.017
R24633 vss.n15637 vss.n15635 0.017
R24634 vss.n15686 vss.n15684 0.017
R24635 vss.n15864 vss.n15863 0.017
R24636 vss.n15936 vss.n15924 0.017
R24637 vss.n15976 vss.n15975 0.017
R24638 vss.n16172 vss.n16160 0.017
R24639 vss.n16212 vss.n16211 0.017
R24640 vss.n16272 vss.n16270 0.017
R24641 vss.n16348 vss.n16346 0.017
R24642 vss.n16397 vss.n16395 0.017
R24643 vss.n16584 vss.n16582 0.017
R24644 vss.n16633 vss.n16631 0.017
R24645 vss.n16700 vss.n16699 0.017
R24646 vss.n16879 vss.n16878 0.017
R24647 vss.n16930 vss.n16929 0.017
R24648 vss.n17115 vss.n17114 0.017
R24649 vss.n17166 vss.n17165 0.017
R24650 vss.n169 vss.n158 0.017
R24651 vss.n184 vss.n173 0.017
R24652 vss.n199 vss.n188 0.017
R24653 vss.n243 vss.n241 0.017
R24654 vss.n21631 vss.n21630 0.017
R24655 vss.n3580 vss.n3579 0.017
R24656 vss.n19623 vss.n19587 0.016
R24657 vss.n6233 vss.n6197 0.016
R24658 vss.n20377 vss.n20376 0.016
R24659 vss.n17500 vss.n17497 0.016
R24660 vss.n20801 vss.n20799 0.016
R24661 vss.n21903 vss.n21902 0.016
R24662 vss.n21888 vss.n21887 0.016
R24663 vss.n10389 vss.n10388 0.016
R24664 vss.n12541 vss.n12536 0.016
R24665 vss.n12148 vss.n12108 0.016
R24666 vss.n14840 vss.n14837 0.016
R24667 vss.n14865 vss.n14855 0.016
R24668 vss.n3852 vss.n3851 0.016
R24669 vss.n3837 vss.n3836 0.016
R24670 vss.n6987 vss.n6986 0.016
R24671 vss.n4110 vss.n4107 0.016
R24672 vss.n7411 vss.n7409 0.016
R24673 vss.n1996 vss.n1995 0.016
R24674 vss.n3218 vss.n3216 0.016
R24675 vss.n3433 vss.n3431 0.016
R24676 vss.n15518 vss.n15516 0.016
R24677 vss.n15577 vss.n15567 0.016
R24678 vss.n15754 vss.n15752 0.016
R24679 vss.n16045 vss.n16033 0.016
R24680 vss.n16103 vss.n16102 0.016
R24681 vss.n16465 vss.n16463 0.016
R24682 vss.n16524 vss.n16514 0.016
R24683 vss.n16999 vss.n16998 0.016
R24684 vss.n17057 vss.n17045 0.016
R24685 vss.n17235 vss.n17234 0.016
R24686 vss.n17317 vss.n15217 0.016
R24687 vss.n457 vss.n456 0.016
R24688 vss.n23041 vss.n23040 0.016
R24689 vss.n1408 vss.n1406 0.016
R24690 vss.n16781 vss.n16779 0.016
R24691 vss.n16784 vss.n16781 0.016
R24692 vss.n10245 vss.n10244 0.016
R24693 vss.n10269 vss.n10268 0.016
R24694 vss.n10289 vss.n10288 0.016
R24695 vss.n10312 vss.n10311 0.016
R24696 vss.n10330 vss.n10329 0.016
R24697 vss.n10372 vss.n10371 0.016
R24698 vss.n10404 vss.n10403 0.016
R24699 vss.n10438 vss.n10437 0.016
R24700 vss.n8938 vss.n8937 0.016
R24701 vss.n8956 vss.n8955 0.016
R24702 vss.n8994 vss.n8993 0.016
R24703 vss.n9024 vss.n9023 0.016
R24704 vss.n9055 vss.n9054 0.016
R24705 vss.n9086 vss.n9085 0.016
R24706 vss.n9105 vss.n9104 0.016
R24707 vss.n9135 vss.n9134 0.016
R24708 vss.n21916 vss.n21915 0.016
R24709 vss.n3865 vss.n3864 0.016
R24710 vss.n9647 vss.n9646 0.015
R24711 vss.n18950 vss.n17679 0.015
R24712 vss.n18949 vss.n18948 0.015
R24713 vss.n18832 vss.n17782 0.015
R24714 vss.n18824 vss.n17794 0.015
R24715 vss.n18710 vss.n18709 0.015
R24716 vss.n18708 vss.n18707 0.015
R24717 vss.n18591 vss.n17995 0.015
R24718 vss.n18583 vss.n18007 0.015
R24719 vss.n18469 vss.n18468 0.015
R24720 vss.n18467 vss.n18466 0.015
R24721 vss.n18350 vss.n18208 0.015
R24722 vss.n18342 vss.n18220 0.015
R24723 vss.n20225 vss.n19082 0.015
R24724 vss.n20217 vss.n19094 0.015
R24725 vss.n20096 vss.n19186 0.015
R24726 vss.n20095 vss.n20094 0.015
R24727 vss.n19978 vss.n19289 0.015
R24728 vss.n19970 vss.n19301 0.015
R24729 vss.n19849 vss.n19393 0.015
R24730 vss.n19848 vss.n19847 0.015
R24731 vss.n19731 vss.n19496 0.015
R24732 vss.n19723 vss.n19508 0.015
R24733 vss.n20384 vss.n17572 0.015
R24734 vss.n20401 vss.n17552 0.015
R24735 vss.n20516 vss.n20505 0.015
R24736 vss.n21865 vss.n21863 0.015
R24737 vss.n21946 vss.n21941 0.015
R24738 vss.n21954 vss.n21953 0.015
R24739 vss.n9684 vss.n9683 0.015
R24740 vss.n10239 vss.n10238 0.015
R24741 vss.n10231 vss.n10230 0.015
R24742 vss.n10378 vss.n10377 0.015
R24743 vss.n12923 vss.n12906 0.015
R24744 vss.n12510 vss.n12493 0.015
R24745 vss.n12874 vss.n12863 0.015
R24746 vss.n3814 vss.n3812 0.015
R24747 vss.n3895 vss.n3890 0.015
R24748 vss.n3903 vss.n3902 0.015
R24749 vss.n5560 vss.n4289 0.015
R24750 vss.n5559 vss.n5558 0.015
R24751 vss.n5442 vss.n4392 0.015
R24752 vss.n5434 vss.n4404 0.015
R24753 vss.n5320 vss.n5319 0.015
R24754 vss.n5318 vss.n5317 0.015
R24755 vss.n5201 vss.n4605 0.015
R24756 vss.n5193 vss.n4617 0.015
R24757 vss.n5079 vss.n5078 0.015
R24758 vss.n5077 vss.n5076 0.015
R24759 vss.n4960 vss.n4818 0.015
R24760 vss.n4952 vss.n4830 0.015
R24761 vss.n6835 vss.n5692 0.015
R24762 vss.n6827 vss.n5704 0.015
R24763 vss.n6706 vss.n5796 0.015
R24764 vss.n6705 vss.n6704 0.015
R24765 vss.n6588 vss.n5899 0.015
R24766 vss.n6580 vss.n5911 0.015
R24767 vss.n6459 vss.n6003 0.015
R24768 vss.n6458 vss.n6457 0.015
R24769 vss.n6341 vss.n6106 0.015
R24770 vss.n6333 vss.n6118 0.015
R24771 vss.n6994 vss.n4182 0.015
R24772 vss.n7011 vss.n4162 0.015
R24773 vss.n7126 vss.n7115 0.015
R24774 vss.n15387 vss.n15385 0.015
R24775 vss.n15464 vss.n15462 0.015
R24776 vss.n15623 vss.n15621 0.015
R24777 vss.n15700 vss.n15698 0.015
R24778 vss.n15851 vss.n15849 0.015
R24779 vss.n15922 vss.n15910 0.015
R24780 vss.n15990 vss.n15989 0.015
R24781 vss.n16158 vss.n16146 0.015
R24782 vss.n16226 vss.n16225 0.015
R24783 vss.n15263 vss.n15261 0.015
R24784 vss.n16334 vss.n16332 0.015
R24785 vss.n16411 vss.n16409 0.015
R24786 vss.n16570 vss.n16568 0.015
R24787 vss.n16647 vss.n16645 0.015
R24788 vss.n16714 vss.n16713 0.015
R24789 vss.n16865 vss.n16864 0.015
R24790 vss.n16944 vss.n16943 0.015
R24791 vss.n21977 vss.n21976 0.015
R24792 vss.n3926 vss.n3925 0.015
R24793 vss.n9119 vss.n9117 0.015
R24794 vss.n15311 vss.n15309 0.014
R24795 vss.n15323 vss.n15311 0.014
R24796 vss.n9646 vss.n9642 0.014
R24797 vss.n10352 vss.n10351 0.014
R24798 vss.n19024 vss.n19023 0.014
R24799 vss.n19005 vss.n19004 0.014
R24800 vss.n17732 vss.n17724 0.014
R24801 vss.n18880 vss.n18879 0.014
R24802 vss.n18777 vss.n17833 0.014
R24803 vss.n17856 vss.n17843 0.014
R24804 vss.n17945 vss.n17937 0.014
R24805 vss.n18639 vss.n18638 0.014
R24806 vss.n18536 vss.n18046 0.014
R24807 vss.n18069 vss.n18056 0.014
R24808 vss.n18158 vss.n18150 0.014
R24809 vss.n18398 vss.n18397 0.014
R24810 vss.n18295 vss.n18259 0.014
R24811 vss.n19047 vss.n19046 0.014
R24812 vss.n20170 vss.n19133 0.014
R24813 vss.n20151 vss.n20150 0.014
R24814 vss.n19239 vss.n19231 0.014
R24815 vss.n20026 vss.n20025 0.014
R24816 vss.n19923 vss.n19340 0.014
R24817 vss.n19904 vss.n19903 0.014
R24818 vss.n19446 vss.n19438 0.014
R24819 vss.n19779 vss.n19778 0.014
R24820 vss.n19676 vss.n19547 0.014
R24821 vss.n19657 vss.n19656 0.014
R24822 vss.n20364 vss.n17583 0.014
R24823 vss.n20405 vss.n20404 0.014
R24824 vss.n20363 vss.n20362 0.014
R24825 vss.n20399 vss.n17557 0.014
R24826 vss.n21758 vss.n21701 0.014
R24827 vss.n14911 vss.n14908 0.014
R24828 vss.n3707 vss.n3650 0.014
R24829 vss.n5634 vss.n5633 0.014
R24830 vss.n5615 vss.n5614 0.014
R24831 vss.n4342 vss.n4334 0.014
R24832 vss.n5490 vss.n5489 0.014
R24833 vss.n5387 vss.n4443 0.014
R24834 vss.n4466 vss.n4453 0.014
R24835 vss.n4555 vss.n4547 0.014
R24836 vss.n5249 vss.n5248 0.014
R24837 vss.n5146 vss.n4656 0.014
R24838 vss.n4679 vss.n4666 0.014
R24839 vss.n4768 vss.n4760 0.014
R24840 vss.n5008 vss.n5007 0.014
R24841 vss.n4905 vss.n4869 0.014
R24842 vss.n5657 vss.n5656 0.014
R24843 vss.n6780 vss.n5743 0.014
R24844 vss.n6761 vss.n6760 0.014
R24845 vss.n5849 vss.n5841 0.014
R24846 vss.n6636 vss.n6635 0.014
R24847 vss.n6533 vss.n5950 0.014
R24848 vss.n6514 vss.n6513 0.014
R24849 vss.n6056 vss.n6048 0.014
R24850 vss.n6389 vss.n6388 0.014
R24851 vss.n6286 vss.n6157 0.014
R24852 vss.n6267 vss.n6266 0.014
R24853 vss.n6974 vss.n4193 0.014
R24854 vss.n7015 vss.n7014 0.014
R24855 vss.n6973 vss.n6972 0.014
R24856 vss.n7009 vss.n4167 0.014
R24857 vss.n8248 vss.n8244 0.014
R24858 vss.n17101 vss.n17100 0.014
R24859 vss.n17180 vss.n17179 0.014
R24860 vss.n10225 vss.n10224 0.014
R24861 vss.n9674 vss.n9673 0.014
R24862 vss.n21605 vss.n21604 0.013
R24863 vss.n21913 vss.n21912 0.013
R24864 vss.n3862 vss.n3861 0.013
R24865 vss.n9649 vss.n9647 0.013
R24866 vss.n21629 vss.n21628 0.013
R24867 vss.n3578 vss.n3577 0.013
R24868 vss.n18962 vss.n18961 0.013
R24869 vss.n18938 vss.n18937 0.013
R24870 vss.n18834 vss.n17776 0.013
R24871 vss.n17798 vss.n17795 0.013
R24872 vss.n18719 vss.n17882 0.013
R24873 vss.n18697 vss.n18696 0.013
R24874 vss.n18593 vss.n17989 0.013
R24875 vss.n18011 vss.n18008 0.013
R24876 vss.n18478 vss.n18095 0.013
R24877 vss.n18456 vss.n18455 0.013
R24878 vss.n18352 vss.n18202 0.013
R24879 vss.n18224 vss.n18221 0.013
R24880 vss.n18269 vss.n17623 0.013
R24881 vss.n20290 vss.n20289 0.013
R24882 vss.n20227 vss.n19076 0.013
R24883 vss.n19098 vss.n19095 0.013
R24884 vss.n20108 vss.n20107 0.013
R24885 vss.n20084 vss.n20083 0.013
R24886 vss.n19980 vss.n19283 0.013
R24887 vss.n19305 vss.n19302 0.013
R24888 vss.n19861 vss.n19860 0.013
R24889 vss.n19837 vss.n19836 0.013
R24890 vss.n19733 vss.n19490 0.013
R24891 vss.n19512 vss.n19509 0.013
R24892 vss.n19621 vss.n19589 0.013
R24893 vss.n20366 vss.n17581 0.013
R24894 vss.n20380 vss.n17574 0.013
R24895 vss.n20536 vss.n20534 0.013
R24896 vss.n20669 ldomc_0.otaldom_0.nmosbn1m_0.vss 0.013
R24897 vss.n9657 vss.n9656 0.013
R24898 vss.n9649 vss.n9648 0.013
R24899 vss.n9642 vss.n9641 0.013
R24900 vss.n9746 vss.n9745 0.013
R24901 vss.n9740 vss.n9739 0.013
R24902 vss.n9734 vss.n9733 0.013
R24903 vss.n9728 vss.n9727 0.013
R24904 vss.n9722 vss.n9721 0.013
R24905 vss.n9716 vss.n9715 0.013
R24906 vss.n9705 vss.n9704 0.013
R24907 vss.n9676 vss.n9675 0.013
R24908 vss.n10192 vss.n10191 0.013
R24909 vss.n10198 vss.n10197 0.013
R24910 vss.n10204 vss.n10203 0.013
R24911 vss.n10210 vss.n10209 0.013
R24912 vss.n9661 vss.n9660 0.013
R24913 vss.n10336 vss.n10334 0.013
R24914 vss.n10336 vss.n10335 0.013
R24915 vss.n10451 vss.n10447 0.013
R24916 vss.n8980 vss.n8979 0.013
R24917 vss.n12176 vss.n12174 0.013
R24918 vss.n12190 vss.n12188 0.013
R24919 vss.n12025 vss.n12023 0.013
R24920 vss.n11980 vss.n11978 0.013
R24921 vss.n11968 vss.n11967 0.013
R24922 vss.n11950 vss.n11940 0.013
R24923 vss.n11222 vss.n11221 0.013
R24924 vss.n11148 vss.n11101 0.013
R24925 vss.n14092 vss.n14078 0.013
R24926 vss.n14078 vss.n13758 0.013
R24927 vss.n11832 vss.n11495 0.013
R24928 vss.n11848 vss.n11832 0.013
R24929 vss.n14975 vss.n13152 0.013
R24930 vss.n12710 vss.n12334 0.013
R24931 vss.n14421 vss.n14268 0.013
R24932 vss.n14314 vss.n14304 0.013
R24933 vss.n14056 vss.n14054 0.013
R24934 vss.n11628 vss.n11618 0.013
R24935 vss.n11639 vss.n11629 0.013
R24936 vss.n11667 vss.n11666 0.013
R24937 vss.n14804 vss.n14794 0.013
R24938 vss.n14790 vss.n14780 0.013
R24939 vss.n14686 vss.n14684 0.013
R24940 vss.n14619 vss.n14617 0.013
R24941 vss.n14607 vss.n14606 0.013
R24942 vss.n14597 vss.n14587 0.013
R24943 vss.n14446 vss.n14445 0.013
R24944 vss.n13235 vss.n13234 0.013
R24945 vss.n14976 vss.n14975 0.013
R24946 vss.n15010 vss.n15009 0.013
R24947 vss.n15025 vss.n15024 0.013
R24948 vss.n15041 vss.n15040 0.013
R24949 vss.n12859 vss.n12847 0.013
R24950 vss.n5572 vss.n5571 0.013
R24951 vss.n5548 vss.n5547 0.013
R24952 vss.n5444 vss.n4386 0.013
R24953 vss.n4408 vss.n4405 0.013
R24954 vss.n5329 vss.n4492 0.013
R24955 vss.n5307 vss.n5306 0.013
R24956 vss.n5203 vss.n4599 0.013
R24957 vss.n4621 vss.n4618 0.013
R24958 vss.n5088 vss.n4705 0.013
R24959 vss.n5066 vss.n5065 0.013
R24960 vss.n4962 vss.n4812 0.013
R24961 vss.n4834 vss.n4831 0.013
R24962 vss.n4879 vss.n4233 0.013
R24963 vss.n6900 vss.n6899 0.013
R24964 vss.n6837 vss.n5686 0.013
R24965 vss.n5708 vss.n5705 0.013
R24966 vss.n6718 vss.n6717 0.013
R24967 vss.n6694 vss.n6693 0.013
R24968 vss.n6590 vss.n5893 0.013
R24969 vss.n5915 vss.n5912 0.013
R24970 vss.n6471 vss.n6470 0.013
R24971 vss.n6447 vss.n6446 0.013
R24972 vss.n6343 vss.n6100 0.013
R24973 vss.n6122 vss.n6119 0.013
R24974 vss.n6231 vss.n6199 0.013
R24975 vss.n6976 vss.n4191 0.013
R24976 vss.n6990 vss.n4184 0.013
R24977 vss.n7146 vss.n7144 0.013
R24978 vss.n7279 bandgapmd_0.otam_1.nmosbn1m_0.vss 0.013
R24979 vss.n8130 vss.n8129 0.013
R24980 vss.n8128 vss.n8127 0.013
R24981 vss.n7922 vss.n7921 0.013
R24982 vss.n7920 vss.n7919 0.013
R24983 vss.n7713 vss.n7712 0.013
R24984 vss.n7711 vss.n7710 0.013
R24985 vss.n7505 vss.n7504 0.013
R24986 vss.n15504 vss.n15502 0.013
R24987 vss.n15591 vss.n15581 0.013
R24988 vss.n15740 vss.n15738 0.013
R24989 vss.n16031 vss.n16019 0.013
R24990 vss.n16117 vss.n16116 0.013
R24991 vss.n15303 vss.n15301 0.013
R24992 vss.n16451 vss.n16449 0.013
R24993 vss.n16538 vss.n16528 0.013
R24994 vss.n16755 vss.n16754 0.013
R24995 vss.n16985 vss.n16984 0.013
R24996 vss.n17071 vss.n17059 0.013
R24997 vss.n17221 vss.n17220 0.013
R24998 vss.n9071 vss.n9069 0.013
R24999 vss.n20405 vss.n17554 0.012
R25000 vss.n7015 vss.n4164 0.012
R25001 vss.n21628 vss.n21627 0.012
R25002 vss.n3577 vss.n3576 0.012
R25003 vss.n17650 vss.n17649 0.012
R25004 vss.n18902 vss.n18901 0.012
R25005 vss.n17756 vss.n17742 0.012
R25006 vss.n17832 vss.n17824 0.012
R25007 vss.n18755 vss.n18754 0.012
R25008 vss.n18661 vss.n18660 0.012
R25009 vss.n17969 vss.n17955 0.012
R25010 vss.n18045 vss.n18037 0.012
R25011 vss.n18514 vss.n18513 0.012
R25012 vss.n18420 vss.n18419 0.012
R25013 vss.n18182 vss.n18168 0.012
R25014 vss.n18258 vss.n18250 0.012
R25015 vss.n19056 vss.n19054 0.012
R25016 vss.n19132 vss.n19124 0.012
R25017 vss.n19157 vss.n19156 0.012
R25018 vss.n20048 vss.n20047 0.012
R25019 vss.n19263 vss.n19249 0.012
R25020 vss.n19339 vss.n19331 0.012
R25021 vss.n19364 vss.n19363 0.012
R25022 vss.n19801 vss.n19800 0.012
R25023 vss.n19470 vss.n19456 0.012
R25024 vss.n19546 vss.n19538 0.012
R25025 vss.n19571 vss.n19570 0.012
R25026 vss.n20518 vss.n20516 0.012
R25027 vss.n20576 vss.n20565 0.012
R25028 vss.n20655 vss.n20654 0.012
R25029 vss.n20657 ldomc_0.otaldom_0.nmosbn1m_0.vss 0.012
R25030 vss.n21519 vss.n21518 0.012
R25031 vss.n21517 vss.n21516 0.012
R25032 vss.n21311 vss.n21310 0.012
R25033 vss.n21309 vss.n21308 0.012
R25034 vss.n21103 vss.n21102 0.012
R25035 vss.n21101 vss.n21100 0.012
R25036 vss.n20895 vss.n20894 0.012
R25037 vss.n22007 vss.n22004 0.012
R25038 vss.n22049 vss.n21978 0.012
R25039 vss.n21969 vss.n21967 0.012
R25040 vss.n21751 vss.n21748 0.012
R25041 vss.n21653 vss.n21652 0.012
R25042 vss.n21656 vss.n21641 0.012
R25043 vss.n21750 vss.n21704 0.012
R25044 vss.n21753 vss.n21704 0.012
R25045 vss.n22052 vss.n21802 0.012
R25046 vss.n22050 vss.n21950 0.012
R25047 vss.n10210 vss.n10208 0.012
R25048 vss.n10208 vss.n10204 0.012
R25049 vss.n10204 vss.n10202 0.012
R25050 vss.n10202 vss.n10198 0.012
R25051 vss.n10198 vss.n10196 0.012
R25052 vss.n10196 vss.n10192 0.012
R25053 vss.n9703 vss.n9676 0.012
R25054 vss.n9705 vss.n9703 0.012
R25055 vss.n9716 vss.n9714 0.012
R25056 vss.n9720 vss.n9716 0.012
R25057 vss.n9722 vss.n9720 0.012
R25058 vss.n9726 vss.n9722 0.012
R25059 vss.n9728 vss.n9726 0.012
R25060 vss.n9732 vss.n9728 0.012
R25061 vss.n9734 vss.n9732 0.012
R25062 vss.n9738 vss.n9734 0.012
R25063 vss.n9740 vss.n9738 0.012
R25064 vss.n9744 vss.n9740 0.012
R25065 vss.n9746 vss.n9744 0.012
R25066 vss.n10183 vss.n9746 0.012
R25067 vss.n10425 vss.n10424 0.012
R25068 vss.n10430 vss.n10429 0.012
R25069 vss.n10452 vss.n10451 0.012
R25070 vss.n12590 vss.n12589 0.012
R25071 vss.n14110 vss.n14109 0.012
R25072 vss.n14095 vss.n14094 0.012
R25073 vss.n13756 vss.n13755 0.012
R25074 vss.n13742 vss.n13740 0.012
R25075 vss.n11439 vss.n11437 0.012
R25076 vss.n11453 vss.n11452 0.012
R25077 vss.n11851 vss.n11850 0.012
R25078 vss.n11866 vss.n11865 0.012
R25079 vss.n13095 vss.n13094 0.012
R25080 vss.n13081 vss.n13079 0.012
R25081 vss.n12317 vss.n12316 0.012
R25082 vss.n14411 vss.n14410 0.012
R25083 vss.n14385 vss.n14377 0.012
R25084 vss.n14953 vss.n14951 0.012
R25085 vss.n14967 vss.n14966 0.012
R25086 vss.n14896 vss.n14884 0.012
R25087 vss.n3956 vss.n3953 0.012
R25088 vss.n3998 vss.n3927 0.012
R25089 vss.n3918 vss.n3916 0.012
R25090 vss.n3700 vss.n3697 0.012
R25091 vss.n3602 vss.n3601 0.012
R25092 vss.n3605 vss.n3590 0.012
R25093 vss.n3699 vss.n3653 0.012
R25094 vss.n3702 vss.n3653 0.012
R25095 vss.n4001 vss.n3751 0.012
R25096 vss.n3999 vss.n3899 0.012
R25097 vss.n4260 vss.n4259 0.012
R25098 vss.n5512 vss.n5511 0.012
R25099 vss.n4366 vss.n4352 0.012
R25100 vss.n4442 vss.n4434 0.012
R25101 vss.n5365 vss.n5364 0.012
R25102 vss.n5271 vss.n5270 0.012
R25103 vss.n4579 vss.n4565 0.012
R25104 vss.n4655 vss.n4647 0.012
R25105 vss.n5124 vss.n5123 0.012
R25106 vss.n5030 vss.n5029 0.012
R25107 vss.n4792 vss.n4778 0.012
R25108 vss.n4868 vss.n4860 0.012
R25109 vss.n5666 vss.n5664 0.012
R25110 vss.n5742 vss.n5734 0.012
R25111 vss.n5767 vss.n5766 0.012
R25112 vss.n6658 vss.n6657 0.012
R25113 vss.n5873 vss.n5859 0.012
R25114 vss.n5949 vss.n5941 0.012
R25115 vss.n5974 vss.n5973 0.012
R25116 vss.n6411 vss.n6410 0.012
R25117 vss.n6080 vss.n6066 0.012
R25118 vss.n6156 vss.n6148 0.012
R25119 vss.n6181 vss.n6180 0.012
R25120 vss.n7128 vss.n7126 0.012
R25121 vss.n7186 vss.n7175 0.012
R25122 vss.n7265 vss.n7264 0.012
R25123 vss.n7267 bandgapmd_0.otam_1.nmosbn1m_0.vss 0.012
R25124 vss.n8230 vss.n8216 0.012
R25125 vss.n8042 vss.n8041 0.012
R25126 vss.n8021 vss.n8007 0.012
R25127 vss.n7833 vss.n7832 0.012
R25128 vss.n7812 vss.n7798 0.012
R25129 vss.n7625 vss.n7624 0.012
R25130 vss.n7604 vss.n7590 0.012
R25131 vss.n8754 vss.n8753 0.012
R25132 vss.n8752 vss.n8751 0.012
R25133 vss.n8546 vss.n8545 0.012
R25134 vss.n8544 vss.n8543 0.012
R25135 vss.n8338 vss.n8337 0.012
R25136 vss.n8336 vss.n8335 0.012
R25137 vss.n15373 vss.n15371 0.012
R25138 vss.n15478 vss.n15476 0.012
R25139 vss.n15609 vss.n15607 0.012
R25140 vss.n15714 vss.n15712 0.012
R25141 vss.n15837 vss.n15835 0.012
R25142 vss.n15908 vss.n15896 0.012
R25143 vss.n16004 vss.n16003 0.012
R25144 vss.n16144 vss.n16132 0.012
R25145 vss.n16240 vss.n16239 0.012
R25146 vss.n15277 vss.n15275 0.012
R25147 vss.n16320 vss.n16318 0.012
R25148 vss.n16425 vss.n16423 0.012
R25149 vss.n16556 vss.n16554 0.012
R25150 vss.n16661 vss.n16659 0.012
R25151 vss.n16728 vss.n16727 0.012
R25152 vss.n16851 vss.n16850 0.012
R25153 vss.n16958 vss.n16957 0.012
R25154 vss.n17087 vss.n17086 0.012
R25155 vss.n17194 vss.n17193 0.012
R25156 vss.n22591 vss.n22590 0.012
R25157 vss.n22589 vss.n22588 0.012
R25158 vss.n22383 vss.n22382 0.012
R25159 vss.n22381 vss.n22380 0.012
R25160 vss.n22175 vss.n22174 0.012
R25161 vss.n22173 vss.n22172 0.012
R25162 vss.n10431 vss.n10430 0.012
R25163 vss.n10383 vss.n10382 0.012
R25164 vss.n20406 vss.n17550 0.011
R25165 vss.n7016 vss.n4160 0.011
R25166 vss.n10304 vss.n10298 0.011
R25167 vss.n10364 vss.n10363 0.011
R25168 vss.n18971 vss.n17666 0.011
R25169 vss.n17695 vss.n17692 0.011
R25170 vss.n18846 vss.n18845 0.011
R25171 vss.n18811 vss.n18810 0.011
R25172 vss.n18721 vss.n17876 0.011
R25173 vss.n17908 vss.n17905 0.011
R25174 vss.n18605 vss.n18604 0.011
R25175 vss.n18570 vss.n18569 0.011
R25176 vss.n18480 vss.n18089 0.011
R25177 vss.n18121 vss.n18118 0.011
R25178 vss.n18364 vss.n18363 0.011
R25179 vss.n18329 vss.n18328 0.011
R25180 vss.n20239 vss.n20238 0.011
R25181 vss.n20204 vss.n20203 0.011
R25182 vss.n20117 vss.n19173 0.011
R25183 vss.n19202 vss.n19199 0.011
R25184 vss.n19992 vss.n19991 0.011
R25185 vss.n19957 vss.n19956 0.011
R25186 vss.n19870 vss.n19380 0.011
R25187 vss.n19409 vss.n19406 0.011
R25188 vss.n19745 vss.n19744 0.011
R25189 vss.n19710 vss.n19709 0.011
R25190 vss.n17589 vss.n17586 0.011
R25191 vss.n17579 vss.n17574 0.011
R25192 vss.n20547 vss.n20546 0.011
R25193 vss.n21431 vss.n21430 0.011
R25194 vss.n21410 vss.n21396 0.011
R25195 vss.n21223 vss.n21222 0.011
R25196 vss.n21202 vss.n21188 0.011
R25197 vss.n21015 vss.n21014 0.011
R25198 vss.n20994 vss.n20980 0.011
R25199 vss.n21950 vss.n21949 0.011
R25200 vss.n21918 vss.n21911 0.011
R25201 vss.n21621 vss.n21620 0.011
R25202 vss.n21626 vss.n21624 0.011
R25203 vss.n10249 vss.n10239 0.011
R25204 vss.n10250 vss.n10231 0.011
R25205 vss.n10323 vss.n10322 0.011
R25206 vss.n10354 vss.n10323 0.011
R25207 vss.n12818 vss.n12800 0.011
R25208 vss.n12562 vss.n12544 0.011
R25209 vss.n12588 vss.n12575 0.011
R25210 vss.n12301 vss.n12036 0.011
R25211 vss.n12009 vss.n12008 0.011
R25212 vss.n11996 vss.n11995 0.011
R25213 vss.n11993 vss.n11992 0.011
R25214 vss.n11956 vss.n11955 0.011
R25215 vss.n11953 vss.n11952 0.011
R25216 vss.n13453 vss.n13452 0.011
R25217 vss.n13111 vss.n13110 0.011
R25218 vss.n10634 vss.n10632 0.011
R25219 vss.n10648 vss.n10647 0.011
R25220 vss.n10725 vss.n10686 0.011
R25221 vss.n14078 vss.n14077 0.011
R25222 vss.n14041 vss.n14040 0.011
R25223 vss.n14028 vss.n14027 0.011
R25224 vss.n11643 vss.n11642 0.011
R25225 vss.n11655 vss.n11654 0.011
R25226 vss.n14700 vss.n14699 0.011
R25227 vss.n14670 vss.n14669 0.011
R25228 vss.n14646 vss.n14645 0.011
R25229 vss.n14632 vss.n14631 0.011
R25230 vss.n14604 vss.n14603 0.011
R25231 vss.n14601 vss.n14600 0.011
R25232 vss.n12844 vss.n12832 0.011
R25233 vss.n3899 vss.n3898 0.011
R25234 vss.n3867 vss.n3860 0.011
R25235 vss.n3570 vss.n3569 0.011
R25236 vss.n3575 vss.n3573 0.011
R25237 vss.n5581 vss.n4276 0.011
R25238 vss.n4305 vss.n4302 0.011
R25239 vss.n5456 vss.n5455 0.011
R25240 vss.n5421 vss.n5420 0.011
R25241 vss.n5331 vss.n4486 0.011
R25242 vss.n4518 vss.n4515 0.011
R25243 vss.n5215 vss.n5214 0.011
R25244 vss.n5180 vss.n5179 0.011
R25245 vss.n5090 vss.n4699 0.011
R25246 vss.n4731 vss.n4728 0.011
R25247 vss.n4974 vss.n4973 0.011
R25248 vss.n4939 vss.n4938 0.011
R25249 vss.n6849 vss.n6848 0.011
R25250 vss.n6814 vss.n6813 0.011
R25251 vss.n6727 vss.n5783 0.011
R25252 vss.n5812 vss.n5809 0.011
R25253 vss.n6602 vss.n6601 0.011
R25254 vss.n6567 vss.n6566 0.011
R25255 vss.n6480 vss.n5990 0.011
R25256 vss.n6019 vss.n6016 0.011
R25257 vss.n6355 vss.n6354 0.011
R25258 vss.n6320 vss.n6319 0.011
R25259 vss.n4199 vss.n4196 0.011
R25260 vss.n4189 vss.n4184 0.011
R25261 vss.n7157 vss.n7156 0.011
R25262 vss.n8144 vss.n8143 0.011
R25263 vss.n8125 vss.n8113 0.011
R25264 vss.n7936 vss.n7935 0.011
R25265 vss.n7917 vss.n7905 0.011
R25266 vss.n7727 vss.n7726 0.011
R25267 vss.n7708 vss.n7696 0.011
R25268 vss.n7519 vss.n7518 0.011
R25269 vss.n8874 vss.n8873 0.011
R25270 vss.n8853 vss.n8839 0.011
R25271 vss.n8666 vss.n8665 0.011
R25272 vss.n8645 vss.n8631 0.011
R25273 vss.n8458 vss.n8457 0.011
R25274 vss.n8437 vss.n8423 0.011
R25275 vss.n15369 vss.n15359 0.011
R25276 vss.n15490 vss.n15488 0.011
R25277 vss.n15605 vss.n15595 0.011
R25278 vss.n15726 vss.n15724 0.011
R25279 vss.n15833 vss.n15823 0.011
R25280 vss.n15895 vss.n15894 0.011
R25281 vss.n16017 vss.n16005 0.011
R25282 vss.n16131 vss.n16130 0.011
R25283 vss.n15289 vss.n15287 0.011
R25284 vss.n16316 vss.n16306 0.011
R25285 vss.n16437 vss.n16435 0.011
R25286 vss.n16552 vss.n16542 0.011
R25287 vss.n16741 vss.n16740 0.011
R25288 vss.n16971 vss.n16970 0.011
R25289 vss.n17085 vss.n17073 0.011
R25290 vss.n17207 vss.n17206 0.011
R25291 vss.n22711 vss.n22710 0.011
R25292 vss.n22690 vss.n22676 0.011
R25293 vss.n22503 vss.n22502 0.011
R25294 vss.n22482 vss.n22468 0.011
R25295 vss.n22295 vss.n22294 0.011
R25296 vss.n22274 vss.n22260 0.011
R25297 vss.n20386 vss.n17566 0.01
R25298 vss.n6996 vss.n4176 0.01
R25299 vss.n10246 vss.n10245 0.01
R25300 vss.n10270 vss.n10269 0.01
R25301 vss.n10290 vss.n10289 0.01
R25302 vss.n10313 vss.n10312 0.01
R25303 vss.n10331 vss.n10330 0.01
R25304 vss.n10373 vss.n10372 0.01
R25305 vss.n10405 vss.n10404 0.01
R25306 vss.n10439 vss.n10438 0.01
R25307 vss.n8937 vss.n8936 0.01
R25308 vss.n8955 vss.n8954 0.01
R25309 vss.n8995 vss.n8994 0.01
R25310 vss.n9025 vss.n9024 0.01
R25311 vss.n9056 vss.n9055 0.01
R25312 vss.n9087 vss.n9086 0.01
R25313 vss.n9106 vss.n9105 0.01
R25314 vss.n9136 vss.n9135 0.01
R25315 vss.n17659 vss.n17657 0.01
R25316 vss.n18913 vss.n17714 0.01
R25317 vss.n18868 vss.n18867 0.01
R25318 vss.n18789 vss.n18788 0.01
R25319 vss.n18744 vss.n18743 0.01
R25320 vss.n18672 vss.n17927 0.01
R25321 vss.n18627 vss.n18626 0.01
R25322 vss.n18548 vss.n18547 0.01
R25323 vss.n18503 vss.n18502 0.01
R25324 vss.n18431 vss.n18140 0.01
R25325 vss.n18386 vss.n18385 0.01
R25326 vss.n18307 vss.n18306 0.01
R25327 vss.n20261 vss.n20260 0.01
R25328 vss.n20182 vss.n20181 0.01
R25329 vss.n19166 vss.n19164 0.01
R25330 vss.n20059 vss.n19221 0.01
R25331 vss.n20014 vss.n20013 0.01
R25332 vss.n19935 vss.n19934 0.01
R25333 vss.n19373 vss.n19371 0.01
R25334 vss.n19812 vss.n19428 0.01
R25335 vss.n19767 vss.n19766 0.01
R25336 vss.n19688 vss.n19687 0.01
R25337 vss.n19580 vss.n19578 0.01
R25338 vss.n20365 vss.n20364 0.01
R25339 vss.n20370 vss.n17577 0.01
R25340 vss.n20363 vss.n17580 0.01
R25341 vss.n20372 vss.n20371 0.01
R25342 vss.n20392 vss.n17563 0.01
R25343 vss.n20502 vss.n20500 0.01
R25344 vss.n21533 vss.n21532 0.01
R25345 vss.n21514 vss.n21502 0.01
R25346 vss.n21445 vss.n21444 0.01
R25347 vss.n21394 vss.n21382 0.01
R25348 vss.n21325 vss.n21324 0.01
R25349 vss.n21306 vss.n21294 0.01
R25350 vss.n21237 vss.n21236 0.01
R25351 vss.n21186 vss.n21174 0.01
R25352 vss.n21117 vss.n21116 0.01
R25353 vss.n21098 vss.n21086 0.01
R25354 vss.n21029 vss.n21028 0.01
R25355 vss.n20978 vss.n20966 0.01
R25356 vss.n20909 vss.n20908 0.01
R25357 vss.n21905 vss.n21903 0.01
R25358 vss.n22014 vss.n22011 0.01
R25359 vss.n21806 vss.n21803 0.01
R25360 vss.n21922 vss.n21920 0.01
R25361 vss.n21784 vss.n21783 0.01
R25362 vss.n21669 vss.n21668 0.01
R25363 vss.n22052 vss.n22051 0.01
R25364 vss.n21634 vss.n21633 0.01
R25365 vss.n9642 vss.n9640 0.01
R25366 vss.n9655 vss.n9649 0.01
R25367 vss.n9657 vss.n9655 0.01
R25368 vss.n10184 vss.n10183 0.01
R25369 vss.n10388 vss.n10387 0.01
R25370 vss.n12609 vss.n12608 0.01
R25371 vss.n12264 vss.n12248 0.01
R25372 vss.n11184 vss.n11183 0.01
R25373 vss.n11169 vss.n11162 0.01
R25374 vss.n13950 vss.n13935 0.01
R25375 vss.n14724 vss.n14723 0.01
R25376 vss.n14912 vss.n14911 0.01
R25377 vss.n3854 vss.n3852 0.01
R25378 vss.n3963 vss.n3960 0.01
R25379 vss.n3755 vss.n3752 0.01
R25380 vss.n3871 vss.n3869 0.01
R25381 vss.n3733 vss.n3732 0.01
R25382 vss.n3618 vss.n3617 0.01
R25383 vss.n4001 vss.n4000 0.01
R25384 vss.n4269 vss.n4267 0.01
R25385 vss.n5523 vss.n4324 0.01
R25386 vss.n5478 vss.n5477 0.01
R25387 vss.n5399 vss.n5398 0.01
R25388 vss.n5354 vss.n5353 0.01
R25389 vss.n5282 vss.n4537 0.01
R25390 vss.n5237 vss.n5236 0.01
R25391 vss.n5158 vss.n5157 0.01
R25392 vss.n5113 vss.n5112 0.01
R25393 vss.n5041 vss.n4750 0.01
R25394 vss.n4996 vss.n4995 0.01
R25395 vss.n4917 vss.n4916 0.01
R25396 vss.n6871 vss.n6870 0.01
R25397 vss.n6792 vss.n6791 0.01
R25398 vss.n5776 vss.n5774 0.01
R25399 vss.n6669 vss.n5831 0.01
R25400 vss.n6624 vss.n6623 0.01
R25401 vss.n6545 vss.n6544 0.01
R25402 vss.n5983 vss.n5981 0.01
R25403 vss.n6422 vss.n6038 0.01
R25404 vss.n6377 vss.n6376 0.01
R25405 vss.n6298 vss.n6297 0.01
R25406 vss.n6190 vss.n6188 0.01
R25407 vss.n6975 vss.n6974 0.01
R25408 vss.n6980 vss.n4187 0.01
R25409 vss.n6973 vss.n4190 0.01
R25410 vss.n6982 vss.n6981 0.01
R25411 vss.n7002 vss.n4173 0.01
R25412 vss.n7112 vss.n7110 0.01
R25413 vss.n8213 vss.n8201 0.01
R25414 vss.n8056 vss.n8055 0.01
R25415 vss.n8005 vss.n7993 0.01
R25416 vss.n7847 vss.n7846 0.01
R25417 vss.n7796 vss.n7784 0.01
R25418 vss.n7639 vss.n7638 0.01
R25419 vss.n7588 vss.n7576 0.01
R25420 vss.n3583 vss.n3582 0.01
R25421 vss.n8888 vss.n8887 0.01
R25422 vss.n8837 vss.n8825 0.01
R25423 vss.n8768 vss.n8767 0.01
R25424 vss.n8749 vss.n8737 0.01
R25425 vss.n8680 vss.n8679 0.01
R25426 vss.n8629 vss.n8617 0.01
R25427 vss.n8560 vss.n8559 0.01
R25428 vss.n8541 vss.n8529 0.01
R25429 vss.n8472 vss.n8471 0.01
R25430 vss.n8421 vss.n8409 0.01
R25431 vss.n8352 vss.n8351 0.01
R25432 vss.n8333 vss.n8321 0.01
R25433 vss.n8264 vss.n8263 0.01
R25434 vss.n1743 vss.n1742 0.01
R25435 vss.n15492 vss.n15490 0.01
R25436 vss.n15595 vss.n15593 0.01
R25437 vss.n15728 vss.n15726 0.01
R25438 vss.n15823 vss.n15821 0.01
R25439 vss.n15894 vss.n15882 0.01
R25440 vss.n16018 vss.n16017 0.01
R25441 vss.n16130 vss.n16118 0.01
R25442 vss.n15291 vss.n15289 0.01
R25443 vss.n16306 vss.n16304 0.01
R25444 vss.n16439 vss.n16437 0.01
R25445 vss.n16542 vss.n16540 0.01
R25446 vss.n16742 vss.n16741 0.01
R25447 vss.n16972 vss.n16971 0.01
R25448 vss.n22725 vss.n22724 0.01
R25449 vss.n22674 vss.n22662 0.01
R25450 vss.n22605 vss.n22604 0.01
R25451 vss.n22586 vss.n22574 0.01
R25452 vss.n22517 vss.n22516 0.01
R25453 vss.n22466 vss.n22454 0.01
R25454 vss.n22397 vss.n22396 0.01
R25455 vss.n22378 vss.n22366 0.01
R25456 vss.n22309 vss.n22308 0.01
R25457 vss.n22258 vss.n22246 0.01
R25458 vss.n22189 vss.n22188 0.01
R25459 vss.n22170 vss.n22158 0.01
R25460 vss.n22101 vss.n22100 0.01
R25461 vss.n204 vss.n203 0.01
R25462 vss.n22053 vss.n21639 0.01
R25463 vss.n4002 vss.n3588 0.01
R25464 vss.n20389 vss.n20388 0.01
R25465 vss.n6999 vss.n6998 0.01
R25466 vss.n20382 vss.n17567 0.009
R25467 vss.n6992 vss.n4177 0.009
R25468 vss.n18973 vss.n17660 0.009
R25469 vss.n18924 vss.n18923 0.009
R25470 vss.n18855 vss.n17763 0.009
R25471 vss.n18801 vss.n17813 0.009
R25472 vss.n18733 vss.n18732 0.009
R25473 vss.n18683 vss.n18682 0.009
R25474 vss.n18614 vss.n17976 0.009
R25475 vss.n18560 vss.n18026 0.009
R25476 vss.n18492 vss.n18491 0.009
R25477 vss.n18442 vss.n18441 0.009
R25478 vss.n18373 vss.n18189 0.009
R25479 vss.n18319 vss.n18239 0.009
R25480 vss.n20248 vss.n19063 0.009
R25481 vss.n20194 vss.n19113 0.009
R25482 vss.n20119 vss.n19167 0.009
R25483 vss.n20070 vss.n20069 0.009
R25484 vss.n20001 vss.n19270 0.009
R25485 vss.n19947 vss.n19320 0.009
R25486 vss.n19872 vss.n19374 0.009
R25487 vss.n19823 vss.n19822 0.009
R25488 vss.n19754 vss.n19477 0.009
R25489 vss.n19700 vss.n19527 0.009
R25490 vss.n19625 vss.n19581 0.009
R25491 vss.n20474 vss.n20472 0.009
R25492 vss.n20799 vss.n20798 0.009
R25493 vss.n21547 vss.n21546 0.009
R25494 vss.n21500 vss.n21488 0.009
R25495 vss.n21339 vss.n21338 0.009
R25496 vss.n21292 vss.n21280 0.009
R25497 vss.n21131 vss.n21130 0.009
R25498 vss.n21084 vss.n21072 0.009
R25499 vss.n20923 vss.n20922 0.009
R25500 vss.n22011 vss.n22009 0.009
R25501 vss.n21793 vss.n21685 0.009
R25502 vss.n21793 vss.n21792 0.009
R25503 vss.n21758 vss.n21757 0.009
R25504 vss.n22065 vss.n22063 0.009
R25505 vss.n10187 vss.n10186 0.009
R25506 vss.n10409 vss.n10408 0.009
R25507 vss.n15059 vss.n15041 0.009
R25508 vss.n12593 vss.n12592 0.009
R25509 vss.n11316 vss.n11305 0.009
R25510 vss.n11817 vss.n11806 0.009
R25511 vss.n14532 vss.n14529 0.009
R25512 vss.n14881 vss.n14869 0.009
R25513 vss.n3960 vss.n3958 0.009
R25514 vss.n3742 vss.n3634 0.009
R25515 vss.n3742 vss.n3741 0.009
R25516 vss.n3707 vss.n3706 0.009
R25517 vss.n5583 vss.n4270 0.009
R25518 vss.n5534 vss.n5533 0.009
R25519 vss.n5465 vss.n4373 0.009
R25520 vss.n5411 vss.n4423 0.009
R25521 vss.n5343 vss.n5342 0.009
R25522 vss.n5293 vss.n5292 0.009
R25523 vss.n5224 vss.n4586 0.009
R25524 vss.n5170 vss.n4636 0.009
R25525 vss.n5102 vss.n5101 0.009
R25526 vss.n5052 vss.n5051 0.009
R25527 vss.n4983 vss.n4799 0.009
R25528 vss.n4929 vss.n4849 0.009
R25529 vss.n6858 vss.n5673 0.009
R25530 vss.n6804 vss.n5723 0.009
R25531 vss.n6729 vss.n5777 0.009
R25532 vss.n6680 vss.n6679 0.009
R25533 vss.n6611 vss.n5880 0.009
R25534 vss.n6557 vss.n5930 0.009
R25535 vss.n6482 vss.n5984 0.009
R25536 vss.n6433 vss.n6432 0.009
R25537 vss.n6364 vss.n6087 0.009
R25538 vss.n6310 vss.n6137 0.009
R25539 vss.n6235 vss.n6191 0.009
R25540 vss.n7084 vss.n7082 0.009
R25541 vss.n7409 vss.n7408 0.009
R25542 vss.n8199 vss.n8187 0.009
R25543 vss.n8158 vss.n8157 0.009
R25544 vss.n8111 vss.n8099 0.009
R25545 vss.n8070 vss.n8069 0.009
R25546 vss.n7991 vss.n7979 0.009
R25547 vss.n7950 vss.n7949 0.009
R25548 vss.n7903 vss.n7891 0.009
R25549 vss.n7862 vss.n7861 0.009
R25550 vss.n7782 vss.n7770 0.009
R25551 vss.n7741 vss.n7740 0.009
R25552 vss.n7694 vss.n7682 0.009
R25553 vss.n7653 vss.n7652 0.009
R25554 vss.n7574 vss.n7562 0.009
R25555 vss.n7533 vss.n7532 0.009
R25556 vss.n4014 vss.n4012 0.009
R25557 vss.n8782 vss.n8781 0.009
R25558 vss.n8735 vss.n8723 0.009
R25559 vss.n8574 vss.n8573 0.009
R25560 vss.n8527 vss.n8515 0.009
R25561 vss.n8366 vss.n8365 0.009
R25562 vss.n8319 vss.n8307 0.009
R25563 vss.n1875 vss.n1874 0.009
R25564 vss.n1878 vss.n1876 0.009
R25565 vss.n2120 vss.n2119 0.009
R25566 vss.n2123 vss.n2121 0.009
R25567 vss.n2364 vss.n2363 0.009
R25568 vss.n2367 vss.n2365 0.009
R25569 vss.n2608 vss.n2607 0.009
R25570 vss.n2612 vss.n2610 0.009
R25571 vss.n2847 vss.n2846 0.009
R25572 vss.n2850 vss.n2848 0.009
R25573 vss.n3091 vss.n3090 0.009
R25574 vss.n3094 vss.n3092 0.009
R25575 vss.n3336 vss.n3335 0.009
R25576 vss.n3339 vss.n3337 0.009
R25577 vss.n15195 vss.n15194 0.009
R25578 vss.n15194 vss.n15190 0.009
R25579 vss.n15156 vss.n15155 0.009
R25580 vss.n17073 vss.n17072 0.009
R25581 vss.n17208 vss.n17207 0.009
R25582 vss.n22619 vss.n22618 0.009
R25583 vss.n22572 vss.n22560 0.009
R25584 vss.n22411 vss.n22410 0.009
R25585 vss.n22364 vss.n22352 0.009
R25586 vss.n22203 vss.n22202 0.009
R25587 vss.n22156 vss.n22144 0.009
R25588 vss.n336 vss.n335 0.009
R25589 vss.n339 vss.n337 0.009
R25590 vss.n581 vss.n580 0.009
R25591 vss.n584 vss.n582 0.009
R25592 vss.n825 vss.n824 0.009
R25593 vss.n828 vss.n826 0.009
R25594 vss.n1069 vss.n1068 0.009
R25595 vss.n1073 vss.n1071 0.009
R25596 vss.n23411 vss.n23409 0.009
R25597 vss.n23408 vss.n23407 0.009
R25598 vss.n23168 vss.n23166 0.009
R25599 vss.n23165 vss.n23164 0.009
R25600 vss.n22923 vss.n22921 0.009
R25601 vss.n22920 vss.n22919 0.009
R25602 vss.n22829 vss.n22828 0.009
R25603 vss.n22828 vss.n22824 0.009
R25604 vss.n22790 vss.n22789 0.009
R25605 vss.n12735 vss.n10457 0.009
R25606 vss.n21895 vss.n21893 0.009
R25607 vss.n3844 vss.n3842 0.009
R25608 vss.n21893 vss.n21892 0.008
R25609 vss.n3842 vss.n3841 0.008
R25610 vss.n18984 vss.n18983 0.008
R25611 vss.n17713 vss.n17705 0.008
R25612 vss.n18857 vss.n18856 0.008
R25613 vss.n18800 vss.n17814 0.008
R25614 vss.n17875 vss.n17863 0.008
R25615 vss.n17926 vss.n17918 0.008
R25616 vss.n18616 vss.n18615 0.008
R25617 vss.n18559 vss.n18027 0.008
R25618 vss.n18088 vss.n18076 0.008
R25619 vss.n18139 vss.n18131 0.008
R25620 vss.n18375 vss.n18374 0.008
R25621 vss.n18318 vss.n18240 0.008
R25622 vss.n20250 vss.n20249 0.008
R25623 vss.n20193 vss.n19114 0.008
R25624 vss.n20130 vss.n20129 0.008
R25625 vss.n19220 vss.n19212 0.008
R25626 vss.n20003 vss.n20002 0.008
R25627 vss.n19946 vss.n19321 0.008
R25628 vss.n19883 vss.n19882 0.008
R25629 vss.n19427 vss.n19419 0.008
R25630 vss.n19756 vss.n19755 0.008
R25631 vss.n19699 vss.n19528 0.008
R25632 vss.n19636 vss.n19635 0.008
R25633 vss.n19617 vss.n19589 0.008
R25634 vss.n20487 vss.n20485 0.008
R25635 vss.n21577 vss.n21576 0.008
R25636 vss.n21459 vss.n21458 0.008
R25637 vss.n21380 vss.n21368 0.008
R25638 vss.n21251 vss.n21250 0.008
R25639 vss.n21172 vss.n21160 0.008
R25640 vss.n21043 vss.n21042 0.008
R25641 vss.n20964 vss.n20952 0.008
R25642 vss.n22048 vss.n22046 0.008
R25643 vss.n21856 vss.n21854 0.008
R25644 vss.n21820 vss.n21810 0.008
R25645 vss.n22049 vss.n21990 0.008
R25646 vss.n21674 vss.n21672 0.008
R25647 vss.n21752 vss.n21747 0.008
R25648 vss.n21777 vss.n21776 0.008
R25649 vss.n21800 vss.n21799 0.008
R25650 vss.n10445 vss.n10444 0.008
R25651 vss.n12776 vss.n12775 0.008
R25652 vss.n11924 vss.n11914 0.008
R25653 vss.n11204 vss.n11203 0.008
R25654 vss.n11200 vss.n11199 0.008
R25655 vss.n11832 vss.n11677 0.008
R25656 vss.n14557 vss.n14547 0.008
R25657 vss.n14882 vss.n14881 0.008
R25658 vss.n3997 vss.n3995 0.008
R25659 vss.n3805 vss.n3803 0.008
R25660 vss.n3769 vss.n3759 0.008
R25661 vss.n3998 vss.n3939 0.008
R25662 vss.n3623 vss.n3621 0.008
R25663 vss.n3701 vss.n3696 0.008
R25664 vss.n3726 vss.n3725 0.008
R25665 vss.n3749 vss.n3748 0.008
R25666 vss.n5594 vss.n5593 0.008
R25667 vss.n4323 vss.n4315 0.008
R25668 vss.n5467 vss.n5466 0.008
R25669 vss.n5410 vss.n4424 0.008
R25670 vss.n4485 vss.n4473 0.008
R25671 vss.n4536 vss.n4528 0.008
R25672 vss.n5226 vss.n5225 0.008
R25673 vss.n5169 vss.n4637 0.008
R25674 vss.n4698 vss.n4686 0.008
R25675 vss.n4749 vss.n4741 0.008
R25676 vss.n4985 vss.n4984 0.008
R25677 vss.n4928 vss.n4850 0.008
R25678 vss.n6860 vss.n6859 0.008
R25679 vss.n6803 vss.n5724 0.008
R25680 vss.n6740 vss.n6739 0.008
R25681 vss.n5830 vss.n5822 0.008
R25682 vss.n6613 vss.n6612 0.008
R25683 vss.n6556 vss.n5931 0.008
R25684 vss.n6493 vss.n6492 0.008
R25685 vss.n6037 vss.n6029 0.008
R25686 vss.n6366 vss.n6365 0.008
R25687 vss.n6309 vss.n6138 0.008
R25688 vss.n6246 vss.n6245 0.008
R25689 vss.n6227 vss.n6199 0.008
R25690 vss.n7097 vss.n7095 0.008
R25691 vss.n8172 vss.n8171 0.008
R25692 vss.n8097 vss.n8085 0.008
R25693 vss.n7964 vss.n7963 0.008
R25694 vss.n7889 vss.n7877 0.008
R25695 vss.n7755 vss.n7754 0.008
R25696 vss.n7680 vss.n7668 0.008
R25697 vss.n7547 vss.n7546 0.008
R25698 vss.n8902 vss.n8901 0.008
R25699 vss.n8823 vss.n8811 0.008
R25700 vss.n8694 vss.n8693 0.008
R25701 vss.n8615 vss.n8603 0.008
R25702 vss.n8486 vss.n8485 0.008
R25703 vss.n8407 vss.n8395 0.008
R25704 vss.n8278 vss.n8277 0.008
R25705 vss.n1861 vss.n1859 0.008
R25706 vss.n1879 vss.n1878 0.008
R25707 vss.n1895 vss.n1893 0.008
R25708 vss.n1993 vss.n1991 0.008
R25709 vss.n2020 vss.n2004 0.008
R25710 vss.n2103 vss.n2101 0.008
R25711 vss.n2105 vss.n2103 0.008
R25712 vss.n2139 vss.n2137 0.008
R25713 vss.n2238 vss.n2236 0.008
R25714 vss.n2264 vss.n2248 0.008
R25715 vss.n2349 vss.n2347 0.008
R25716 vss.n2383 vss.n2381 0.008
R25717 vss.n2482 vss.n2480 0.008
R25718 vss.n2508 vss.n2492 0.008
R25719 vss.n2593 vss.n2591 0.008
R25720 vss.n2628 vss.n2626 0.008
R25721 vss.n2727 vss.n2725 0.008
R25722 vss.n2753 vss.n2737 0.008
R25723 vss.n2833 vss.n2832 0.008
R25724 vss.n2834 bandgapmd_0.otam_1.pdiffaloadm_0.vss 0.008
R25725 vss.n2866 vss.n2864 0.008
R25726 vss.n2965 vss.n2963 0.008
R25727 vss.n2991 vss.n2975 0.008
R25728 vss.n3076 vss.n3074 0.008
R25729 vss.n3110 vss.n3108 0.008
R25730 vss.n3209 vss.n3207 0.008
R25731 vss.n3236 vss.n3220 0.008
R25732 vss.n3320 vss.n3318 0.008
R25733 vss.n3354 vss.n3352 0.008
R25734 vss.n15383 vss.n15373 0.008
R25735 vss.n15476 vss.n15474 0.008
R25736 vss.n15619 vss.n15609 0.008
R25737 vss.n15712 vss.n15710 0.008
R25738 vss.n15847 vss.n15837 0.008
R25739 vss.n15909 vss.n15908 0.008
R25740 vss.n16003 vss.n15991 0.008
R25741 vss.n16145 vss.n16144 0.008
R25742 vss.n16239 vss.n16227 0.008
R25743 vss.n15275 vss.n15273 0.008
R25744 vss.n16330 vss.n16320 0.008
R25745 vss.n16423 vss.n16421 0.008
R25746 vss.n16566 vss.n16556 0.008
R25747 vss.n16659 vss.n16657 0.008
R25748 vss.n16727 vss.n16726 0.008
R25749 vss.n16849 vss.n16837 0.008
R25750 vss.n16863 vss.n16851 0.008
R25751 vss.n16957 vss.n16956 0.008
R25752 vss.n17099 vss.n17087 0.008
R25753 vss.n17193 vss.n17192 0.008
R25754 vss.n22739 vss.n22738 0.008
R25755 vss.n22660 vss.n22648 0.008
R25756 vss.n22531 vss.n22530 0.008
R25757 vss.n22452 vss.n22440 0.008
R25758 vss.n22323 vss.n22322 0.008
R25759 vss.n22244 vss.n22232 0.008
R25760 vss.n22115 vss.n22114 0.008
R25761 vss.n322 vss.n320 0.008
R25762 vss.n340 vss.n339 0.008
R25763 vss.n356 vss.n354 0.008
R25764 vss.n454 vss.n452 0.008
R25765 vss.n481 vss.n465 0.008
R25766 vss.n564 vss.n562 0.008
R25767 vss.n566 vss.n564 0.008
R25768 vss.n600 vss.n598 0.008
R25769 vss.n699 vss.n697 0.008
R25770 vss.n725 vss.n709 0.008
R25771 vss.n810 vss.n808 0.008
R25772 vss.n844 vss.n842 0.008
R25773 vss.n943 vss.n941 0.008
R25774 vss.n969 vss.n953 0.008
R25775 vss.n1054 vss.n1052 0.008
R25776 vss.n1089 vss.n1087 0.008
R25777 vss.n1188 vss.n1186 0.008
R25778 vss.n1214 vss.n1198 0.008
R25779 vss.n1299 vss.n1297 0.008
R25780 ldomc_0.otaldom_0.pdiffaloadm_0.vss vss.n1311 0.008
R25781 vss.n23393 vss.n23391 0.008
R25782 vss.n23309 vss.n23293 0.008
R25783 vss.n23283 vss.n23281 0.008
R25784 vss.n23184 vss.n23182 0.008
R25785 vss.n23150 vss.n23148 0.008
R25786 vss.n23065 vss.n23049 0.008
R25787 vss.n23038 vss.n23036 0.008
R25788 vss.n22940 vss.n22938 0.008
R25789 vss.n22906 vss.n22904 0.008
R25790 vss.n21915 vss.n21914 0.008
R25791 vss.n3864 vss.n3863 0.008
R25792 vss.n10347 vss.n10346 0.008
R25793 vss.n9010 vss.n9007 0.008
R25794 vss.n21906 vss.n21822 0.007
R25795 vss.n3855 vss.n3771 0.007
R25796 vss.n14375 vss.n14365 0.007
R25797 vss.n20405 vss.n17551 0.007
R25798 vss.n18985 vss.n18984 0.007
R25799 vss.n18914 vss.n17713 0.007
R25800 vss.n18857 vss.n17757 0.007
R25801 vss.n17817 vss.n17814 0.007
R25802 vss.n18742 vss.n17863 0.007
R25803 vss.n18673 vss.n17926 0.007
R25804 vss.n18616 vss.n17970 0.007
R25805 vss.n18030 vss.n18027 0.007
R25806 vss.n18501 vss.n18076 0.007
R25807 vss.n18432 vss.n18139 0.007
R25808 vss.n18375 vss.n18183 0.007
R25809 vss.n18243 vss.n18240 0.007
R25810 vss.n20250 vss.n19057 0.007
R25811 vss.n19117 vss.n19114 0.007
R25812 vss.n20131 vss.n20130 0.007
R25813 vss.n20060 vss.n19220 0.007
R25814 vss.n20003 vss.n19264 0.007
R25815 vss.n19324 vss.n19321 0.007
R25816 vss.n19884 vss.n19883 0.007
R25817 vss.n19813 vss.n19427 0.007
R25818 vss.n19756 vss.n19471 0.007
R25819 vss.n19531 vss.n19528 0.007
R25820 vss.n19637 vss.n19636 0.007
R25821 vss.n20382 vss.n20381 0.007
R25822 vss.n20489 vss.n20487 0.007
R25823 vss.n20654 vss.n20653 0.007
R25824 vss.n20657 vss.n20656 0.007
R25825 vss.n20763 vss.n20749 0.007
R25826 vss.n20764 vss.n20763 0.007
R25827 vss.n20783 vss.n20769 0.007
R25828 vss.n21574 vss.n21562 0.007
R25829 vss.n21561 vss.n21560 0.007
R25830 vss.n21486 vss.n21474 0.007
R25831 vss.n21473 vss.n21472 0.007
R25832 vss.n21366 vss.n21354 0.007
R25833 vss.n21353 vss.n21352 0.007
R25834 vss.n21278 vss.n21266 0.007
R25835 vss.n21265 vss.n21264 0.007
R25836 vss.n21158 vss.n21146 0.007
R25837 vss.n21145 vss.n21144 0.007
R25838 vss.n21070 vss.n21058 0.007
R25839 vss.n21057 vss.n21056 0.007
R25840 vss.n20950 vss.n20938 0.007
R25841 vss.n20937 vss.n20936 0.007
R25842 vss.n22004 vss.n22002 0.007
R25843 vss.n21973 vss.n21970 0.007
R25844 vss.n21781 vss.n21776 0.007
R25845 vss.n21668 vss.n21642 0.007
R25846 vss.n21626 vss.n21622 0.007
R25847 vss.n22058 vss.n22056 0.007
R25848 vss.n10187 bandgapmd_0.bg_trimmup_0.vss 0.007
R25849 vss.n12589 vss.n12588 0.007
R25850 vss.n14700 vss.n13467 0.007
R25851 vss.n12303 vss.n12301 0.007
R25852 vss.n12734 vss.n12733 0.007
R25853 vss.n12714 vss.n12713 0.007
R25854 vss.n12642 vss.n12641 0.007
R25855 vss.n12639 vss.n12638 0.007
R25856 vss.n14974 vss.n14973 0.007
R25857 vss.n12845 vss.n12844 0.007
R25858 vss.n3953 vss.n3951 0.007
R25859 vss.n3922 vss.n3919 0.007
R25860 vss.n3730 vss.n3725 0.007
R25861 vss.n3617 vss.n3591 0.007
R25862 vss.n3575 vss.n3571 0.007
R25863 vss.n7015 vss.n4161 0.007
R25864 vss.n5595 vss.n5594 0.007
R25865 vss.n5524 vss.n4323 0.007
R25866 vss.n5467 vss.n4367 0.007
R25867 vss.n4427 vss.n4424 0.007
R25868 vss.n5352 vss.n4473 0.007
R25869 vss.n5283 vss.n4536 0.007
R25870 vss.n5226 vss.n4580 0.007
R25871 vss.n4640 vss.n4637 0.007
R25872 vss.n5111 vss.n4686 0.007
R25873 vss.n5042 vss.n4749 0.007
R25874 vss.n4985 vss.n4793 0.007
R25875 vss.n4853 vss.n4850 0.007
R25876 vss.n6860 vss.n5667 0.007
R25877 vss.n5727 vss.n5724 0.007
R25878 vss.n6741 vss.n6740 0.007
R25879 vss.n6670 vss.n5830 0.007
R25880 vss.n6613 vss.n5874 0.007
R25881 vss.n5934 vss.n5931 0.007
R25882 vss.n6494 vss.n6493 0.007
R25883 vss.n6423 vss.n6037 0.007
R25884 vss.n6366 vss.n6081 0.007
R25885 vss.n6141 vss.n6138 0.007
R25886 vss.n6247 vss.n6246 0.007
R25887 vss.n6992 vss.n6991 0.007
R25888 vss.n7099 vss.n7097 0.007
R25889 vss.n7264 vss.n7263 0.007
R25890 vss.n7267 vss.n7266 0.007
R25891 vss.n7373 vss.n7359 0.007
R25892 vss.n7374 vss.n7373 0.007
R25893 vss.n7393 vss.n7379 0.007
R25894 vss.n8185 vss.n8173 0.007
R25895 vss.n8084 vss.n8083 0.007
R25896 vss.n7977 vss.n7965 0.007
R25897 vss.n7876 vss.n7875 0.007
R25898 vss.n7849 vss.n7848 0.007
R25899 vss.n7768 vss.n7756 0.007
R25900 vss.n7667 vss.n7666 0.007
R25901 vss.n7560 vss.n7548 0.007
R25902 vss.n4007 vss.n4005 0.007
R25903 vss.n8916 vss.n8915 0.007
R25904 vss.n8809 vss.n8797 0.007
R25905 vss.n8796 vss.n8795 0.007
R25906 vss.n8721 vss.n8709 0.007
R25907 vss.n8708 vss.n8707 0.007
R25908 vss.n8601 vss.n8589 0.007
R25909 vss.n8588 vss.n8587 0.007
R25910 vss.n8513 vss.n8501 0.007
R25911 vss.n8500 vss.n8499 0.007
R25912 vss.n8393 vss.n8381 0.007
R25913 vss.n8380 vss.n8379 0.007
R25914 vss.n8305 vss.n8293 0.007
R25915 vss.n8292 vss.n8291 0.007
R25916 vss.n8250 vss.n8249 0.007
R25917 vss.n1973 vss.n1971 0.007
R25918 vss.n2036 vss.n2024 0.007
R25919 vss.n2218 vss.n2216 0.007
R25920 vss.n2280 vss.n2268 0.007
R25921 vss.n2462 vss.n2460 0.007
R25922 vss.n2525 vss.n2513 0.007
R25923 vss.n2706 vss.n2704 0.007
R25924 vss.n2769 vss.n2757 0.007
R25925 vss.n2945 vss.n2943 0.007
R25926 vss.n3007 vss.n2995 0.007
R25927 vss.n3189 vss.n3187 0.007
R25928 vss.n3252 vss.n3240 0.007
R25929 vss.n15189 vss.n15175 0.007
R25930 vss.n15175 vss.n15174 0.007
R25931 vss.n15173 vss.n15172 0.007
R25932 vss.n15168 vss.n15157 0.007
R25933 vss.n15506 vss.n15504 0.007
R25934 vss.n15581 vss.n15579 0.007
R25935 vss.n15742 vss.n15740 0.007
R25936 vss.n16032 vss.n16031 0.007
R25937 vss.n16116 vss.n16104 0.007
R25938 vss.n16453 vss.n16451 0.007
R25939 vss.n16528 vss.n16526 0.007
R25940 vss.n16756 vss.n16755 0.007
R25941 vss.n16986 vss.n16985 0.007
R25942 vss.n17059 vss.n17058 0.007
R25943 vss.n17222 vss.n17221 0.007
R25944 vss.n22753 vss.n22752 0.007
R25945 vss.n22646 vss.n22634 0.007
R25946 vss.n22633 vss.n22632 0.007
R25947 vss.n22558 vss.n22546 0.007
R25948 vss.n22545 vss.n22544 0.007
R25949 vss.n22438 vss.n22426 0.007
R25950 vss.n22425 vss.n22424 0.007
R25951 vss.n22350 vss.n22338 0.007
R25952 vss.n22337 vss.n22336 0.007
R25953 vss.n22230 vss.n22218 0.007
R25954 vss.n22217 vss.n22216 0.007
R25955 vss.n22142 vss.n22130 0.007
R25956 vss.n22129 vss.n22128 0.007
R25957 vss.n22087 vss.n22086 0.007
R25958 vss.n434 vss.n432 0.007
R25959 vss.n497 vss.n485 0.007
R25960 vss.n679 vss.n677 0.007
R25961 vss.n741 vss.n729 0.007
R25962 vss.n923 vss.n921 0.007
R25963 vss.n986 vss.n974 0.007
R25964 vss.n1167 vss.n1165 0.007
R25965 vss.n1230 vss.n1218 0.007
R25966 vss.n23325 vss.n23313 0.007
R25967 vss.n23263 vss.n23261 0.007
R25968 vss.n23081 vss.n23069 0.007
R25969 vss.n23018 vss.n23016 0.007
R25970 vss.n22823 vss.n22809 0.007
R25971 vss.n22809 vss.n22808 0.007
R25972 vss.n22807 vss.n22806 0.007
R25973 vss.n22802 vss.n22791 0.007
R25974 vss.n12637 vss.n12632 0.007
R25975 vss.n9714 vss.n9713 0.007
R25976 vss.n10447 vss.n10442 0.006
R25977 vss.n9672 vss.n9671 0.006
R25978 vss.n18973 vss.n18972 0.006
R25979 vss.n18925 vss.n18924 0.006
R25980 vss.n17775 vss.n17763 0.006
R25981 vss.n17813 vss.n17805 0.006
R25982 vss.n18732 vss.n18731 0.006
R25983 vss.n18684 vss.n18683 0.006
R25984 vss.n17988 vss.n17976 0.006
R25985 vss.n18026 vss.n18018 0.006
R25986 vss.n18491 vss.n18490 0.006
R25987 vss.n18443 vss.n18442 0.006
R25988 vss.n18201 vss.n18189 0.006
R25989 vss.n18239 vss.n18231 0.006
R25990 vss.n19075 vss.n19063 0.006
R25991 vss.n19113 vss.n19105 0.006
R25992 vss.n20119 vss.n20118 0.006
R25993 vss.n20071 vss.n20070 0.006
R25994 vss.n19282 vss.n19270 0.006
R25995 vss.n19320 vss.n19312 0.006
R25996 vss.n19872 vss.n19871 0.006
R25997 vss.n19824 vss.n19823 0.006
R25998 vss.n19489 vss.n19477 0.006
R25999 vss.n19527 vss.n19519 0.006
R26000 vss.n19625 vss.n19624 0.006
R26001 vss.n19613 vss.n19593 0.006
R26002 vss.n20360 vss.n17585 0.006
R26003 vss.n20379 vss.n17558 0.006
R26004 vss.n20361 vss.n17584 0.006
R26005 vss.n17570 vss.n17562 0.006
R26006 vss.n20457 vss.n20456 0.006
R26007 vss.n20472 vss.n20470 0.006
R26008 vss.n20591 vss.n20580 0.006
R26009 vss.n20640 vss.n20638 0.006
R26010 vss.n20673 vss.n20671 0.006
R26011 vss.n20746 vss.n20744 0.006
R26012 vss.n20798 vss.n20787 0.006
R26013 vss.n21575 vss.n21574 0.006
R26014 vss.n21472 vss.n21460 0.006
R26015 vss.n21367 vss.n21366 0.006
R26016 vss.n21264 vss.n21252 0.006
R26017 vss.n21159 vss.n21158 0.006
R26018 vss.n21056 vss.n21044 0.006
R26019 vss.n20951 vss.n20950 0.006
R26020 vss.n22060 vss.n22058 0.006
R26021 vss.n9686 vss.n9685 0.006
R26022 vss.n9662 vss.n9661 0.006
R26023 vss.n15060 vss.n15059 0.006
R26024 vss.n12204 vss.n12202 0.006
R26025 vss.n12230 vss.n12229 0.006
R26026 vss.n12244 vss.n12243 0.006
R26027 vss.n12265 vss.n12264 0.006
R26028 vss.n10722 vss.n10721 0.006
R26029 vss.n13012 vss.n13011 0.006
R26030 vss.n12381 vss.n12380 0.006
R26031 vss.n12719 vss.n12718 0.006
R26032 vss.n12694 vss.n12693 0.006
R26033 vss.n11541 vss.n11540 0.006
R26034 vss.n14340 vss.n14330 0.006
R26035 vss.n13884 vss.n13882 0.006
R26036 vss.n13917 vss.n13916 0.006
R26037 vss.n13931 vss.n13930 0.006
R26038 vss.n13951 vss.n13950 0.006
R26039 vss.n14776 vss.n14766 0.006
R26040 vss.n14743 vss.n14733 0.006
R26041 vss.n14729 vss.n14728 0.006
R26042 vss.n14723 vss.n14703 0.006
R26043 vss.n14820 bandgapmd_0.pnp_groupm_0.vss 0.006
R26044 vss.n14975 vss.n14974 0.006
R26045 vss.n14897 vss.n14896 0.006
R26046 vss.n5583 vss.n5582 0.006
R26047 vss.n5535 vss.n5534 0.006
R26048 vss.n4385 vss.n4373 0.006
R26049 vss.n4423 vss.n4415 0.006
R26050 vss.n5342 vss.n5341 0.006
R26051 vss.n5294 vss.n5293 0.006
R26052 vss.n4598 vss.n4586 0.006
R26053 vss.n4636 vss.n4628 0.006
R26054 vss.n5101 vss.n5100 0.006
R26055 vss.n5053 vss.n5052 0.006
R26056 vss.n4811 vss.n4799 0.006
R26057 vss.n4849 vss.n4841 0.006
R26058 vss.n5685 vss.n5673 0.006
R26059 vss.n5723 vss.n5715 0.006
R26060 vss.n6729 vss.n6728 0.006
R26061 vss.n6681 vss.n6680 0.006
R26062 vss.n5892 vss.n5880 0.006
R26063 vss.n5930 vss.n5922 0.006
R26064 vss.n6482 vss.n6481 0.006
R26065 vss.n6434 vss.n6433 0.006
R26066 vss.n6099 vss.n6087 0.006
R26067 vss.n6137 vss.n6129 0.006
R26068 vss.n6235 vss.n6234 0.006
R26069 vss.n6223 vss.n6203 0.006
R26070 vss.n6970 vss.n4195 0.006
R26071 vss.n6989 vss.n4168 0.006
R26072 vss.n6971 vss.n4194 0.006
R26073 vss.n4180 vss.n4172 0.006
R26074 vss.n7067 vss.n7066 0.006
R26075 vss.n7082 vss.n7080 0.006
R26076 vss.n7201 vss.n7190 0.006
R26077 vss.n7250 vss.n7248 0.006
R26078 vss.n7283 vss.n7281 0.006
R26079 vss.n7356 vss.n7354 0.006
R26080 vss.n7408 vss.n7397 0.006
R26081 vss.n8186 vss.n8185 0.006
R26082 vss.n8083 vss.n8071 0.006
R26083 vss.n7978 vss.n7977 0.006
R26084 vss.n7875 vss.n7863 0.006
R26085 vss.n7769 vss.n7768 0.006
R26086 vss.n7666 vss.n7654 0.006
R26087 vss.n7561 vss.n7560 0.006
R26088 vss.n4009 vss.n4007 0.006
R26089 vss.n4017 vss.n4016 0.006
R26090 vss.n8915 vss.n8903 0.006
R26091 vss.n8810 vss.n8809 0.006
R26092 vss.n8707 vss.n8695 0.006
R26093 vss.n8602 vss.n8601 0.006
R26094 vss.n8499 vss.n8487 0.006
R26095 vss.n8394 vss.n8393 0.006
R26096 vss.n8291 vss.n8279 0.006
R26097 vss.n1812 vss.n1801 0.006
R26098 vss.n1846 vss.n1844 0.006
R26099 vss.n1911 vss.n1909 0.006
R26100 vss.n1957 vss.n1955 0.006
R26101 vss.n2052 vss.n2040 0.006
R26102 vss.n2088 vss.n2086 0.006
R26103 vss.n2155 vss.n2153 0.006
R26104 vss.n2202 vss.n2200 0.006
R26105 vss.n2296 vss.n2284 0.006
R26106 vss.n2333 vss.n2331 0.006
R26107 vss.n2400 vss.n2397 0.006
R26108 vss.n2446 vss.n2444 0.006
R26109 vss.n2509 vss.n2508 0.006
R26110 vss.n2541 vss.n2529 0.006
R26111 vss.n2577 vss.n2575 0.006
R26112 vss.n2644 vss.n2642 0.006
R26113 vss.n2690 vss.n2688 0.006
R26114 vss.n2785 vss.n2773 0.006
R26115 vss.n2882 vss.n2880 0.006
R26116 vss.n2929 vss.n2927 0.006
R26117 vss.n3060 vss.n3058 0.006
R26118 vss.n3111 vss.n3110 0.006
R26119 vss.n3127 vss.n3125 0.006
R26120 vss.n3173 vss.n3171 0.006
R26121 vss.n3268 vss.n3256 0.006
R26122 vss.n3304 vss.n3302 0.006
R26123 vss.n3335 vss.n3333 0.006
R26124 vss.n3369 vss.n3367 0.006
R26125 vss.n3412 vss.n3410 0.006
R26126 vss.n15397 vss.n15387 0.006
R26127 vss.n15462 vss.n15460 0.006
R26128 vss.n15633 vss.n15623 0.006
R26129 vss.n15698 vss.n15696 0.006
R26130 vss.n15309 vss.n15308 0.006
R26131 vss.n15324 vss.n15323 0.006
R26132 vss.n15861 vss.n15851 0.006
R26133 vss.n15923 vss.n15922 0.006
R26134 vss.n15989 vss.n15977 0.006
R26135 vss.n16159 vss.n16158 0.006
R26136 vss.n16225 vss.n16213 0.006
R26137 vss.n15261 vss.n15259 0.006
R26138 vss.n16344 vss.n16334 0.006
R26139 vss.n16409 vss.n16407 0.006
R26140 vss.n16580 vss.n16570 0.006
R26141 vss.n16645 vss.n16643 0.006
R26142 vss.n16713 vss.n16712 0.006
R26143 vss.n16779 vss.n16778 0.006
R26144 vss.n16796 vss.n16784 0.006
R26145 vss.n16877 vss.n16865 0.006
R26146 vss.n16943 vss.n16942 0.006
R26147 vss.n17113 vss.n17101 0.006
R26148 vss.n17179 vss.n17178 0.006
R26149 vss.n22752 vss.n22740 0.006
R26150 vss.n22647 vss.n22646 0.006
R26151 vss.n22544 vss.n22532 0.006
R26152 vss.n22439 vss.n22438 0.006
R26153 vss.n22336 vss.n22324 0.006
R26154 vss.n22231 vss.n22230 0.006
R26155 vss.n22128 vss.n22116 0.006
R26156 vss.n273 vss.n262 0.006
R26157 vss.n307 vss.n305 0.006
R26158 vss.n372 vss.n370 0.006
R26159 vss.n418 vss.n416 0.006
R26160 vss.n513 vss.n501 0.006
R26161 vss.n549 vss.n547 0.006
R26162 vss.n616 vss.n614 0.006
R26163 vss.n663 vss.n661 0.006
R26164 vss.n757 vss.n745 0.006
R26165 vss.n794 vss.n792 0.006
R26166 vss.n861 vss.n858 0.006
R26167 vss.n907 vss.n905 0.006
R26168 vss.n970 vss.n969 0.006
R26169 vss.n1002 vss.n990 0.006
R26170 vss.n1038 vss.n1036 0.006
R26171 vss.n1105 vss.n1103 0.006
R26172 vss.n1151 vss.n1149 0.006
R26173 vss.n1246 vss.n1234 0.006
R26174 vss.n23377 vss.n23375 0.006
R26175 vss.n23341 vss.n23329 0.006
R26176 vss.n23200 vss.n23198 0.006
R26177 vss.n23148 vss.n23146 0.006
R26178 vss.n23133 vss.n23131 0.006
R26179 vss.n23097 vss.n23085 0.006
R26180 vss.n23002 vss.n23000 0.006
R26181 vss.n22956 vss.n22954 0.006
R26182 vss.n22924 vss.n22923 0.006
R26183 vss.n22891 vss.n22889 0.006
R26184 vss.n22857 vss.n22846 0.006
R26185 vss.n21948 vss.n21947 0.006
R26186 vss.n21947 vss.n21919 0.006
R26187 vss.n3897 vss.n3896 0.006
R26188 vss.n3896 vss.n3868 0.006
R26189 vss.n21910 vss.n21909 0.005
R26190 vss.n21909 vss.n21908 0.005
R26191 vss.n3859 vss.n3858 0.005
R26192 vss.n3858 vss.n3857 0.005
R26193 vss.n13407 vss.n13406 0.005
R26194 vss.n21801 vss.n21640 0.005
R26195 vss.n3750 vss.n3589 0.005
R26196 vss.n17657 vss.n17651 0.005
R26197 vss.n17717 vss.n17714 0.005
R26198 vss.n18869 vss.n18868 0.005
R26199 vss.n18788 vss.n18787 0.005
R26200 vss.n18744 vss.n17857 0.005
R26201 vss.n17930 vss.n17927 0.005
R26202 vss.n18628 vss.n18627 0.005
R26203 vss.n18547 vss.n18546 0.005
R26204 vss.n18503 vss.n18070 0.005
R26205 vss.n18143 vss.n18140 0.005
R26206 vss.n18387 vss.n18386 0.005
R26207 vss.n18306 vss.n18305 0.005
R26208 vss.n20262 vss.n20261 0.005
R26209 vss.n20181 vss.n20180 0.005
R26210 vss.n19164 vss.n19158 0.005
R26211 vss.n19224 vss.n19221 0.005
R26212 vss.n20015 vss.n20014 0.005
R26213 vss.n19934 vss.n19933 0.005
R26214 vss.n19371 vss.n19365 0.005
R26215 vss.n19431 vss.n19428 0.005
R26216 vss.n19768 vss.n19767 0.005
R26217 vss.n19687 vss.n19686 0.005
R26218 vss.n19578 vss.n19572 0.005
R26219 vss.n19593 vss.n19592 0.005
R26220 vss.n20504 vss.n20502 0.005
R26221 vss.n20580 vss.n20578 0.005
R26222 vss.n20625 vss.n20623 0.005
R26223 vss.n20688 vss.n20686 0.005
R26224 vss.n20731 vss.n20729 0.005
R26225 vss.n20814 vss.n20803 0.005
R26226 vss.n20849 vss.n20847 0.005
R26227 vss.n21560 vss.n21548 0.005
R26228 vss.n21487 vss.n21486 0.005
R26229 vss.n21352 vss.n21340 0.005
R26230 vss.n21279 vss.n21278 0.005
R26231 vss.n21144 vss.n21132 0.005
R26232 vss.n21071 vss.n21070 0.005
R26233 vss.n20936 vss.n20924 0.005
R26234 vss.n21887 vss.n21886 0.005
R26235 vss.n21810 vss.n21809 0.005
R26236 vss.n21939 vss.n21938 0.005
R26237 vss.n21966 vss.n21965 0.005
R26238 vss.n21739 vss.n21705 0.005
R26239 vss.n21711 vss.n21705 0.005
R26240 vss.n21785 vss.n21784 0.005
R26241 vss.n21650 vss.n21644 0.005
R26242 vss.n21639 vss.n21637 0.005
R26243 vss.n22067 vss.n22065 0.005
R26244 vss.n9640 vss.n9203 0.005
R26245 vss.n9662 vss.n9657 0.005
R26246 vss.n10192 bandgapmd_0.bg_trimmup_0.vss 0.005
R26247 vss.n8933 vss.n8930 0.005
R26248 vss.n12822 vss.n12819 0.005
R26249 vss.n15010 vss.n12818 0.005
R26250 vss.n12490 vss.n12489 0.005
R26251 vss.n12589 vss.n12562 0.005
R26252 vss.n14547 vss.n14164 0.005
R26253 vss.n11914 vss.n11913 0.005
R26254 vss.n12730 vss.n12729 0.005
R26255 vss.n12712 vss.n12711 0.005
R26256 vss.n14410 vss.n14385 0.005
R26257 vss.n12860 vss.n12859 0.005
R26258 vss.n3836 vss.n3835 0.005
R26259 vss.n3759 vss.n3758 0.005
R26260 vss.n3888 vss.n3887 0.005
R26261 vss.n3915 vss.n3914 0.005
R26262 vss.n3688 vss.n3654 0.005
R26263 vss.n3660 vss.n3654 0.005
R26264 vss.n3734 vss.n3733 0.005
R26265 vss.n3599 vss.n3593 0.005
R26266 vss.n4267 vss.n4261 0.005
R26267 vss.n4327 vss.n4324 0.005
R26268 vss.n5479 vss.n5478 0.005
R26269 vss.n5398 vss.n5397 0.005
R26270 vss.n5354 vss.n4467 0.005
R26271 vss.n4540 vss.n4537 0.005
R26272 vss.n5238 vss.n5237 0.005
R26273 vss.n5157 vss.n5156 0.005
R26274 vss.n5113 vss.n4680 0.005
R26275 vss.n4753 vss.n4750 0.005
R26276 vss.n4997 vss.n4996 0.005
R26277 vss.n4916 vss.n4915 0.005
R26278 vss.n6872 vss.n6871 0.005
R26279 vss.n6791 vss.n6790 0.005
R26280 vss.n5774 vss.n5768 0.005
R26281 vss.n5834 vss.n5831 0.005
R26282 vss.n6625 vss.n6624 0.005
R26283 vss.n6544 vss.n6543 0.005
R26284 vss.n5981 vss.n5975 0.005
R26285 vss.n6041 vss.n6038 0.005
R26286 vss.n6378 vss.n6377 0.005
R26287 vss.n6297 vss.n6296 0.005
R26288 vss.n6188 vss.n6182 0.005
R26289 vss.n6203 vss.n6202 0.005
R26290 vss.n7114 vss.n7112 0.005
R26291 vss.n7190 vss.n7188 0.005
R26292 vss.n7235 vss.n7233 0.005
R26293 vss.n7298 vss.n7296 0.005
R26294 vss.n7341 vss.n7339 0.005
R26295 vss.n7424 vss.n7413 0.005
R26296 vss.n7459 vss.n7457 0.005
R26297 vss.n8171 vss.n8159 0.005
R26298 vss.n8098 vss.n8097 0.005
R26299 vss.n7963 vss.n7951 0.005
R26300 vss.n7890 vss.n7889 0.005
R26301 vss.n7754 vss.n7742 0.005
R26302 vss.n7681 vss.n7680 0.005
R26303 vss.n7546 vss.n7534 0.005
R26304 vss.n3588 vss.n3586 0.005
R26305 vss.n4016 vss.n4014 0.005
R26306 vss.n8795 vss.n8783 0.005
R26307 vss.n8722 vss.n8721 0.005
R26308 vss.n8587 vss.n8575 0.005
R26309 vss.n8514 vss.n8513 0.005
R26310 vss.n8379 vss.n8367 0.005
R26311 vss.n8306 vss.n8305 0.005
R26312 vss.n1760 vss.n1746 0.005
R26313 vss.n1761 vss.n1760 0.005
R26314 vss.n1780 vss.n1766 0.005
R26315 vss.n1827 vss.n1816 0.005
R26316 vss.n1831 vss.n1829 0.005
R26317 vss.n1927 vss.n1925 0.005
R26318 vss.n1941 vss.n1939 0.005
R26319 vss.n2068 vss.n2056 0.005
R26320 vss.n2072 vss.n2070 0.005
R26321 vss.n2171 vss.n2169 0.005
R26322 vss.n2185 vss.n2183 0.005
R26323 vss.n2313 vss.n2301 0.005
R26324 vss.n2317 vss.n2315 0.005
R26325 vss.n2416 vss.n2414 0.005
R26326 vss.n2430 vss.n2428 0.005
R26327 vss.n2557 vss.n2545 0.005
R26328 vss.n2561 vss.n2559 0.005
R26329 vss.n2660 vss.n2658 0.005
R26330 vss.n2674 vss.n2672 0.005
R26331 vss.n2801 vss.n2789 0.005
R26332 vss.n2805 vss.n2803 0.005
R26333 vss.n2898 vss.n2896 0.005
R26334 vss.n2912 vss.n2910 0.005
R26335 vss.n3012 vss.n3011 0.005
R26336 vss.n3040 vss.n3028 0.005
R26337 vss.n3044 vss.n3042 0.005
R26338 vss.n3143 vss.n3141 0.005
R26339 vss.n3157 vss.n3155 0.005
R26340 vss.n3284 vss.n3272 0.005
R26341 vss.n3288 vss.n3286 0.005
R26342 vss.n3384 vss.n3382 0.005
R26343 vss.n3397 vss.n3395 0.005
R26344 vss.n15359 vss.n15357 0.005
R26345 vss.n15520 vss.n15518 0.005
R26346 vss.n15567 vss.n15565 0.005
R26347 vss.n15756 vss.n15754 0.005
R26348 vss.n15307 vss.n15306 0.005
R26349 vss.n15326 vss.n15325 0.005
R26350 vss.n16046 vss.n16045 0.005
R26351 vss.n16102 vss.n16090 0.005
R26352 vss.n16467 vss.n16465 0.005
R26353 vss.n16514 vss.n16512 0.005
R26354 vss.n16768 vss.n16766 0.005
R26355 vss.n16807 vss.n16797 0.005
R26356 vss.n17000 vss.n16999 0.005
R26357 vss.n22632 vss.n22620 0.005
R26358 vss.n22559 vss.n22558 0.005
R26359 vss.n22424 vss.n22412 0.005
R26360 vss.n22351 vss.n22350 0.005
R26361 vss.n22216 vss.n22204 0.005
R26362 vss.n22143 vss.n22142 0.005
R26363 vss.n221 vss.n207 0.005
R26364 vss.n222 vss.n221 0.005
R26365 vss.n241 vss.n227 0.005
R26366 vss.n288 vss.n277 0.005
R26367 vss.n292 vss.n290 0.005
R26368 vss.n388 vss.n386 0.005
R26369 vss.n402 vss.n400 0.005
R26370 vss.n529 vss.n517 0.005
R26371 vss.n533 vss.n531 0.005
R26372 vss.n632 vss.n630 0.005
R26373 vss.n646 vss.n644 0.005
R26374 vss.n774 vss.n762 0.005
R26375 vss.n778 vss.n776 0.005
R26376 vss.n877 vss.n875 0.005
R26377 vss.n891 vss.n889 0.005
R26378 vss.n1018 vss.n1006 0.005
R26379 vss.n1022 vss.n1020 0.005
R26380 vss.n1121 vss.n1119 0.005
R26381 vss.n1135 vss.n1133 0.005
R26382 vss.n1262 vss.n1250 0.005
R26383 vss.n1266 vss.n1264 0.005
R26384 vss.n23361 vss.n23359 0.005
R26385 vss.n23357 vss.n23345 0.005
R26386 vss.n23247 vss.n23245 0.005
R26387 vss.n23230 vss.n23228 0.005
R26388 vss.n23216 vss.n23214 0.005
R26389 vss.n23117 vss.n23115 0.005
R26390 vss.n23113 vss.n23101 0.005
R26391 vss.n22986 vss.n22984 0.005
R26392 vss.n22972 vss.n22970 0.005
R26393 vss.n22876 vss.n22874 0.005
R26394 vss.n22872 vss.n22861 0.005
R26395 vss.n21650 vss.n21640 0.005
R26396 vss.n3599 vss.n3589 0.005
R26397 vss.n21987 vss.n21986 0.005
R26398 vss.n3936 vss.n3935 0.005
R26399 vss.n12288 vss.n12280 0.004
R26400 vss.n13487 vss.n13479 0.004
R26401 vss.n20384 vss.n17573 0.004
R26402 vss.n6994 vss.n4183 0.004
R26403 vss.n10262 vss.n10261 0.004
R26404 vss.n17678 vss.n17666 0.004
R26405 vss.n18936 vss.n17692 0.004
R26406 vss.n18845 vss.n18844 0.004
R26407 vss.n18812 vss.n18811 0.004
R26408 vss.n18721 vss.n18720 0.004
R26409 vss.n18695 vss.n17905 0.004
R26410 vss.n18604 vss.n18603 0.004
R26411 vss.n18571 vss.n18570 0.004
R26412 vss.n18480 vss.n18479 0.004
R26413 vss.n18454 vss.n18118 0.004
R26414 vss.n18363 vss.n18362 0.004
R26415 vss.n18330 vss.n18329 0.004
R26416 vss.n20238 vss.n20237 0.004
R26417 vss.n20205 vss.n20204 0.004
R26418 vss.n19185 vss.n19173 0.004
R26419 vss.n20082 vss.n19199 0.004
R26420 vss.n19991 vss.n19990 0.004
R26421 vss.n19958 vss.n19957 0.004
R26422 vss.n19392 vss.n19380 0.004
R26423 vss.n19835 vss.n19406 0.004
R26424 vss.n19744 vss.n19743 0.004
R26425 vss.n19711 vss.n19710 0.004
R26426 vss.n20359 vss.n17586 0.004
R26427 vss.n17589 vss.n17583 0.004
R26428 vss.n20456 vss.n20454 0.004
R26429 vss.n20459 vss.n20457 0.004
R26430 vss.n20606 vss.n20595 0.004
R26431 vss.n20610 vss.n20608 0.004
R26432 vss.n20703 vss.n20701 0.004
R26433 vss.n20716 vss.n20714 0.004
R26434 vss.n20829 vss.n20818 0.004
R26435 vss.n20833 vss.n20831 0.004
R26436 vss.n21606 vss.n21579 0.004
R26437 vss.n21578 vss.n21577 0.004
R26438 vss.n21458 vss.n21446 0.004
R26439 vss.n21381 vss.n21380 0.004
R26440 vss.n21250 vss.n21238 0.004
R26441 vss.n21173 vss.n21172 0.004
R26442 vss.n21042 vss.n21030 0.004
R26443 vss.n20965 vss.n20964 0.004
R26444 vss.n21908 vss.n21907 0.004
R26445 vss.n10378 vss.n10376 0.004
R26446 vss.n8999 vss.n8988 0.004
R26447 vss.n9091 vss.n9080 0.004
R26448 vss.n9140 vss.n9129 0.004
R26449 vss.n12591 vss.n12590 0.004
R26450 vss.n12150 vss.n12149 0.004
R26451 vss.n11914 vss.n11330 0.004
R26452 vss.n11290 vss.n11289 0.004
R26453 vss.n11264 vss.n11263 0.004
R26454 vss.n11226 vss.n11224 0.004
R26455 vss.n12733 vss.n12732 0.004
R26456 vss.n12729 vss.n12728 0.004
R26457 vss.n12718 vss.n12717 0.004
R26458 vss.n12715 vss.n12714 0.004
R26459 vss.n12710 vss.n12709 0.004
R26460 vss.n12677 vss.n12676 0.004
R26461 vss.n12661 vss.n12660 0.004
R26462 vss.n12644 vss.n12643 0.004
R26463 vss.n12641 vss.n12640 0.004
R26464 vss.n12638 vss.n12637 0.004
R26465 vss.n11832 vss.n11831 0.004
R26466 vss.n11791 vss.n11790 0.004
R26467 vss.n11754 vss.n11753 0.004
R26468 vss.n11727 vss.n11725 0.004
R26469 vss.n11148 vss.n11147 0.004
R26470 vss.n13310 vss.n13309 0.004
R26471 vss.n14547 vss.n14546 0.004
R26472 vss.n14514 vss.n14513 0.004
R26473 vss.n14476 vss.n14475 0.004
R26474 vss.n14450 vss.n14448 0.004
R26475 vss.n14422 vss.n14421 0.004
R26476 vss.n13234 vss.n13233 0.004
R26477 vss.n14968 vss.n14967 0.004
R26478 vss.n15009 vss.n15008 0.004
R26479 vss.n14911 vss.n14867 0.004
R26480 vss.n3857 vss.n3856 0.004
R26481 vss.n4288 vss.n4276 0.004
R26482 vss.n5546 vss.n4302 0.004
R26483 vss.n5455 vss.n5454 0.004
R26484 vss.n5422 vss.n5421 0.004
R26485 vss.n5331 vss.n5330 0.004
R26486 vss.n5305 vss.n4515 0.004
R26487 vss.n5214 vss.n5213 0.004
R26488 vss.n5181 vss.n5180 0.004
R26489 vss.n5090 vss.n5089 0.004
R26490 vss.n5064 vss.n4728 0.004
R26491 vss.n4973 vss.n4972 0.004
R26492 vss.n4940 vss.n4939 0.004
R26493 vss.n6848 vss.n6847 0.004
R26494 vss.n6815 vss.n6814 0.004
R26495 vss.n5795 vss.n5783 0.004
R26496 vss.n6692 vss.n5809 0.004
R26497 vss.n6601 vss.n6600 0.004
R26498 vss.n6568 vss.n6567 0.004
R26499 vss.n6002 vss.n5990 0.004
R26500 vss.n6445 vss.n6016 0.004
R26501 vss.n6354 vss.n6353 0.004
R26502 vss.n6321 vss.n6320 0.004
R26503 vss.n6969 vss.n4196 0.004
R26504 vss.n4199 vss.n4193 0.004
R26505 vss.n7066 vss.n7064 0.004
R26506 vss.n7069 vss.n7067 0.004
R26507 vss.n7216 vss.n7205 0.004
R26508 vss.n7220 vss.n7218 0.004
R26509 vss.n7313 vss.n7311 0.004
R26510 vss.n7326 vss.n7324 0.004
R26511 vss.n7439 vss.n7428 0.004
R26512 vss.n7443 vss.n7441 0.004
R26513 vss.n8200 vss.n8199 0.004
R26514 vss.n8157 vss.n8145 0.004
R26515 vss.n8112 vss.n8111 0.004
R26516 vss.n8069 vss.n8057 0.004
R26517 vss.n7992 vss.n7991 0.004
R26518 vss.n7949 vss.n7937 0.004
R26519 vss.n7904 vss.n7903 0.004
R26520 vss.n7861 vss.n7849 0.004
R26521 vss.n7783 vss.n7782 0.004
R26522 vss.n7740 vss.n7728 0.004
R26523 vss.n7695 vss.n7694 0.004
R26524 vss.n7652 vss.n7640 0.004
R26525 vss.n7575 vss.n7574 0.004
R26526 vss.n7532 vss.n7520 0.004
R26527 vss.n8901 vss.n8889 0.004
R26528 vss.n8824 vss.n8823 0.004
R26529 vss.n8693 vss.n8681 0.004
R26530 vss.n8616 vss.n8615 0.004
R26531 vss.n8485 vss.n8473 0.004
R26532 vss.n8408 vss.n8407 0.004
R26533 vss.n8277 vss.n8265 0.004
R26534 vss.n1743 vss.n1653 0.004
R26535 vss.n1740 vss.n1738 0.004
R26536 vss.n1797 vss.n1784 0.004
R26537 vss.n1816 vss.n1814 0.004
R26538 vss.n1842 vss.n1831 0.004
R26539 vss.n1925 vss.n1923 0.004
R26540 vss.n1943 vss.n1941 0.004
R26541 vss.n2056 vss.n2054 0.004
R26542 vss.n2084 vss.n2072 0.004
R26543 vss.n2169 vss.n2167 0.004
R26544 vss.n2187 vss.n2185 0.004
R26545 vss.n2301 vss.n2299 0.004
R26546 vss.n2329 vss.n2317 0.004
R26547 vss.n2414 vss.n2412 0.004
R26548 vss.n2432 vss.n2430 0.004
R26549 vss.n2545 vss.n2543 0.004
R26550 vss.n2573 vss.n2561 0.004
R26551 vss.n2658 vss.n2656 0.004
R26552 vss.n2676 vss.n2674 0.004
R26553 vss.n2789 vss.n2787 0.004
R26554 vss.n2816 vss.n2805 0.004
R26555 vss.n2819 vss.n2818 0.004
R26556 vss.n2896 vss.n2894 0.004
R26557 vss.n2915 vss.n2912 0.004
R26558 vss.n3028 vss.n3026 0.004
R26559 vss.n3056 vss.n3044 0.004
R26560 vss.n3141 vss.n3139 0.004
R26561 vss.n3159 vss.n3157 0.004
R26562 vss.n3272 vss.n3270 0.004
R26563 vss.n3300 vss.n3288 0.004
R26564 vss.n3382 vss.n3380 0.004
R26565 vss.n3399 vss.n3397 0.004
R26566 vss.n3450 vss.n3449 0.004
R26567 vss.n15124 vss.n15123 0.004
R26568 vss.n15340 vss.n15330 0.004
R26569 vss.n16821 vss.n16809 0.004
R26570 vss.n17045 vss.n17044 0.004
R26571 vss.n17236 vss.n17235 0.004
R26572 vss.n22738 vss.n22726 0.004
R26573 vss.n22661 vss.n22660 0.004
R26574 vss.n22530 vss.n22518 0.004
R26575 vss.n22453 vss.n22452 0.004
R26576 vss.n22322 vss.n22310 0.004
R26577 vss.n22245 vss.n22244 0.004
R26578 vss.n22114 vss.n22102 0.004
R26579 vss.n204 vss.n114 0.004
R26580 vss.n201 vss.n199 0.004
R26581 vss.n258 vss.n245 0.004
R26582 vss.n277 vss.n275 0.004
R26583 vss.n303 vss.n292 0.004
R26584 vss.n386 vss.n384 0.004
R26585 vss.n404 vss.n402 0.004
R26586 vss.n517 vss.n515 0.004
R26587 vss.n545 vss.n533 0.004
R26588 vss.n630 vss.n628 0.004
R26589 vss.n648 vss.n646 0.004
R26590 vss.n762 vss.n760 0.004
R26591 vss.n790 vss.n778 0.004
R26592 vss.n875 vss.n873 0.004
R26593 vss.n893 vss.n891 0.004
R26594 vss.n1006 vss.n1004 0.004
R26595 vss.n1034 vss.n1022 0.004
R26596 vss.n1119 vss.n1117 0.004
R26597 vss.n1137 vss.n1135 0.004
R26598 vss.n1250 vss.n1248 0.004
R26599 vss.n1278 vss.n1266 0.004
R26600 vss.n1281 vss.n1280 0.004
R26601 vss.n23373 vss.n23361 0.004
R26602 vss.n23345 vss.n23343 0.004
R26603 vss.n23232 vss.n23230 0.004
R26604 vss.n23214 vss.n23212 0.004
R26605 vss.n23129 vss.n23117 0.004
R26606 vss.n23101 vss.n23099 0.004
R26607 vss.n22988 vss.n22986 0.004
R26608 vss.n22970 vss.n22968 0.004
R26609 vss.n22887 vss.n22876 0.004
R26610 vss.n22861 vss.n22859 0.004
R26611 vss.n1425 vss.n1424 0.004
R26612 vss.n22759 vss.n22758 0.004
R26613 vss.n10566 vss.n10560 0.004
R26614 vss.n10567 vss.n10566 0.004
R26615 vss.n12972 vss.n12971 0.004
R26616 vss.n12971 vss.n12963 0.004
R26617 vss.n21637 vss.n21636 0.004
R26618 vss.n3586 vss.n3585 0.004
R26619 vss.n21907 vss.n21906 0.004
R26620 vss.n3856 vss.n3855 0.004
R26621 vss.n9010 vss.n9009 0.004
R26622 vss.n10348 vss.n10347 0.004
R26623 vss.n10395 vss.n10394 0.004
R26624 vss.n10779 vss.n10778 0.003
R26625 vss.n12289 vss.n12288 0.003
R26626 vss.n10778 vss.n10770 0.003
R26627 vss.n13488 vss.n13487 0.003
R26628 vss.n12941 vss.n12940 0.003
R26629 vss.n13182 vss.n13181 0.003
R26630 vss.n13181 vss.n13173 0.003
R26631 vss.n12940 vss.n12932 0.003
R26632 vss.n12351 vss.n12345 0.003
R26633 vss.n12352 vss.n12351 0.003
R26634 vss.n13775 vss.n13769 0.003
R26635 vss.n13815 vss.n13814 0.003
R26636 vss.n13816 vss.n13815 0.003
R26637 vss.n13776 vss.n13775 0.003
R26638 vss.n11511 vss.n11505 0.003
R26639 vss.n11512 vss.n11511 0.003
R26640 vss.n9160 vss.t327 0.003
R26641 vss.n11786 vss.n11776 0.003
R26642 vss.n12663 vss.n12662 0.003
R26643 vss.n17649 vss.n17641 0.003
R26644 vss.n18901 vss.n18900 0.003
R26645 vss.n18878 vss.n17742 0.003
R26646 vss.n18778 vss.n17832 0.003
R26647 vss.n18756 vss.n18755 0.003
R26648 vss.n18660 vss.n18659 0.003
R26649 vss.n18637 vss.n17955 0.003
R26650 vss.n18537 vss.n18045 0.003
R26651 vss.n18515 vss.n18514 0.003
R26652 vss.n18419 vss.n18418 0.003
R26653 vss.n18396 vss.n18168 0.003
R26654 vss.n18296 vss.n18258 0.003
R26655 vss.n19054 vss.n19048 0.003
R26656 vss.n20171 vss.n19132 0.003
R26657 vss.n19156 vss.n19148 0.003
R26658 vss.n20047 vss.n20046 0.003
R26659 vss.n20024 vss.n19249 0.003
R26660 vss.n19924 vss.n19339 0.003
R26661 vss.n19363 vss.n19355 0.003
R26662 vss.n19800 vss.n19799 0.003
R26663 vss.n19777 vss.n19456 0.003
R26664 vss.n19677 vss.n19546 0.003
R26665 vss.n19570 vss.n19562 0.003
R26666 vss.n20376 vss.n17576 0.003
R26667 vss.n20520 vss.n20518 0.003
R26668 vss.n20565 vss.n20563 0.003
R26669 vss.n20595 vss.n20593 0.003
R26670 vss.n20621 vss.n20610 0.003
R26671 vss.n20701 vss.n20699 0.003
R26672 vss.n20718 vss.n20716 0.003
R26673 vss.n20818 vss.n20816 0.003
R26674 vss.n20844 vss.n20833 0.003
R26675 vss.n21546 vss.n21534 0.003
R26676 vss.n21501 vss.n21500 0.003
R26677 vss.n21444 vss.n21432 0.003
R26678 vss.n21395 vss.n21394 0.003
R26679 vss.n21338 vss.n21326 0.003
R26680 vss.n21293 vss.n21292 0.003
R26681 vss.n21236 vss.n21224 0.003
R26682 vss.n21187 vss.n21186 0.003
R26683 vss.n21130 vss.n21118 0.003
R26684 vss.n21085 vss.n21084 0.003
R26685 vss.n21028 vss.n21016 0.003
R26686 vss.n20979 vss.n20978 0.003
R26687 vss.n20922 vss.n20910 0.003
R26688 vss.n9029 vss.n9018 0.003
R26689 vss.n9060 vss.n9049 0.003
R26690 vss.n9111 vss.n9099 0.003
R26691 vss.n12592 vss.n12591 0.003
R26692 vss.n12243 vss.n12242 0.003
R26693 vss.n12245 vss.n12244 0.003
R26694 vss.n12248 vss.n12247 0.003
R26695 vss.n12267 vss.n12265 0.003
R26696 vss.n11978 vss.n11968 0.003
R26697 vss.n11952 vss.n11951 0.003
R26698 vss.n11951 vss.n11950 0.003
R26699 vss.n11940 vss.n11924 0.003
R26700 vss.n11326 vss.n11316 0.003
R26701 vss.n11301 vss.n11291 0.003
R26702 vss.n11291 vss.n11290 0.003
R26703 vss.n11224 vss.n11222 0.003
R26704 vss.n11221 vss.n11219 0.003
R26705 vss.n14094 vss.n14093 0.003
R26706 vss.n13757 vss.n13756 0.003
R26707 vss.n11454 vss.n11453 0.003
R26708 vss.n11850 vss.n11849 0.003
R26709 vss.n13452 vss.n13451 0.003
R26710 vss.n13096 vss.n13095 0.003
R26711 vss.n10649 vss.n10648 0.003
R26712 vss.n12318 vss.n12317 0.003
R26713 vss.n12717 vss.n12716 0.003
R26714 vss.n12716 vss.n12715 0.003
R26715 vss.n12696 vss.n12695 0.003
R26716 vss.n12680 vss.n12679 0.003
R26717 vss.n12643 vss.n12642 0.003
R26718 vss.n12640 vss.n12639 0.003
R26719 vss.n14421 vss.n14411 0.003
R26720 vss.n14377 vss.n14376 0.003
R26721 vss.n14376 vss.n14375 0.003
R26722 vss.n14341 vss.n14340 0.003
R26723 vss.n13930 vss.n13929 0.003
R26724 vss.n13932 vss.n13931 0.003
R26725 vss.n13935 vss.n13934 0.003
R26726 vss.n13953 vss.n13951 0.003
R26727 vss.n11629 vss.n11628 0.003
R26728 vss.n11656 vss.n11655 0.003
R26729 vss.n11666 vss.n11656 0.003
R26730 vss.n11677 vss.n11667 0.003
R26731 vss.n11827 vss.n11817 0.003
R26732 vss.n11802 vss.n11792 0.003
R26733 vss.n11792 vss.n11791 0.003
R26734 vss.n11725 vss.n11723 0.003
R26735 vss.n11133 vss.n11132 0.003
R26736 vss.n14731 vss.n14729 0.003
R26737 vss.n14728 vss.n14727 0.003
R26738 vss.n14726 vss.n14724 0.003
R26739 vss.n14703 vss.n14702 0.003
R26740 vss.n14617 vss.n14607 0.003
R26741 vss.n14600 vss.n14599 0.003
R26742 vss.n14599 vss.n14597 0.003
R26743 vss.n14587 vss.n14557 0.003
R26744 vss.n14542 vss.n14532 0.003
R26745 vss.n14525 vss.n14515 0.003
R26746 vss.n14515 vss.n14514 0.003
R26747 vss.n14448 vss.n14446 0.003
R26748 vss.n14445 vss.n14443 0.003
R26749 vss.n12875 vss.n12874 0.003
R26750 vss.n4259 vss.n4251 0.003
R26751 vss.n5511 vss.n5510 0.003
R26752 vss.n5488 vss.n4352 0.003
R26753 vss.n5388 vss.n4442 0.003
R26754 vss.n5366 vss.n5365 0.003
R26755 vss.n5270 vss.n5269 0.003
R26756 vss.n5247 vss.n4565 0.003
R26757 vss.n5147 vss.n4655 0.003
R26758 vss.n5125 vss.n5124 0.003
R26759 vss.n5029 vss.n5028 0.003
R26760 vss.n5006 vss.n4778 0.003
R26761 vss.n4906 vss.n4868 0.003
R26762 vss.n5664 vss.n5658 0.003
R26763 vss.n6781 vss.n5742 0.003
R26764 vss.n5766 vss.n5758 0.003
R26765 vss.n6657 vss.n6656 0.003
R26766 vss.n6634 vss.n5859 0.003
R26767 vss.n6534 vss.n5949 0.003
R26768 vss.n5973 vss.n5965 0.003
R26769 vss.n6410 vss.n6409 0.003
R26770 vss.n6387 vss.n6066 0.003
R26771 vss.n6287 vss.n6156 0.003
R26772 vss.n6180 vss.n6172 0.003
R26773 vss.n6986 vss.n4186 0.003
R26774 vss.n7130 vss.n7128 0.003
R26775 vss.n7175 vss.n7173 0.003
R26776 vss.n7205 vss.n7203 0.003
R26777 vss.n7231 vss.n7220 0.003
R26778 vss.n7311 vss.n7309 0.003
R26779 vss.n7328 vss.n7326 0.003
R26780 vss.n7428 vss.n7426 0.003
R26781 vss.n7454 vss.n7443 0.003
R26782 vss.n8214 vss.n8213 0.003
R26783 vss.n8055 vss.n8043 0.003
R26784 vss.n8006 vss.n8005 0.003
R26785 vss.n7846 vss.n7834 0.003
R26786 vss.n7797 vss.n7796 0.003
R26787 vss.n7638 vss.n7626 0.003
R26788 vss.n7589 vss.n7588 0.003
R26789 vss.n8249 vss.n8230 0.003
R26790 vss.n8887 vss.n8875 0.003
R26791 vss.n8838 vss.n8837 0.003
R26792 vss.n8781 vss.n8769 0.003
R26793 vss.n8736 vss.n8735 0.003
R26794 vss.n8679 vss.n8667 0.003
R26795 vss.n8630 vss.n8629 0.003
R26796 vss.n8573 vss.n8561 0.003
R26797 vss.n8528 vss.n8527 0.003
R26798 vss.n8471 vss.n8459 0.003
R26799 vss.n8422 vss.n8421 0.003
R26800 vss.n8365 vss.n8353 0.003
R26801 vss.n8320 vss.n8319 0.003
R26802 vss.n8263 vss.n8251 0.003
R26803 vss.n1697 vss.n1695 0.003
R26804 vss.n1710 vss.n1708 0.003
R26805 vss.n1725 vss.n1723 0.003
R26806 vss.n1801 vss.n1799 0.003
R26807 vss.n1959 vss.n1957 0.003
R26808 vss.n2040 vss.n2038 0.003
R26809 vss.n2204 vss.n2202 0.003
R26810 vss.n2284 vss.n2282 0.003
R26811 vss.n2448 vss.n2446 0.003
R26812 vss.n2529 vss.n2527 0.003
R26813 vss.n2692 vss.n2690 0.003
R26814 vss.n2725 vss.n2709 0.003
R26815 vss.n2773 vss.n2771 0.003
R26816 vss.n2931 vss.n2929 0.003
R26817 vss.n3011 vss.n3009 0.003
R26818 vss.n3175 vss.n3173 0.003
R26819 vss.n3256 vss.n3254 0.003
R26820 vss.n3414 vss.n3412 0.003
R26821 vss.n15411 vss.n15401 0.003
R26822 vss.n15448 vss.n15446 0.003
R26823 vss.n15647 vss.n15637 0.003
R26824 vss.n15684 vss.n15682 0.003
R26825 vss.n15354 vss.n15344 0.003
R26826 vss.n15865 vss.n15864 0.003
R26827 vss.n15937 vss.n15936 0.003
R26828 vss.n15975 vss.n15963 0.003
R26829 vss.n16173 vss.n16172 0.003
R26830 vss.n16211 vss.n16199 0.003
R26831 vss.n16282 vss.n16272 0.003
R26832 vss.n16358 vss.n16348 0.003
R26833 vss.n16395 vss.n16393 0.003
R26834 vss.n16594 vss.n16584 0.003
R26835 vss.n16631 vss.n16629 0.003
R26836 vss.n16699 vss.n16698 0.003
R26837 vss.n16835 vss.n16823 0.003
R26838 vss.n16837 vss.n16836 0.003
R26839 vss.n16891 vss.n16879 0.003
R26840 vss.n16929 vss.n16928 0.003
R26841 vss.n17127 vss.n17115 0.003
R26842 vss.n17165 vss.n17164 0.003
R26843 vss.n16266 vss.n16265 0.003
R26844 vss.n22724 vss.n22712 0.003
R26845 vss.n22675 vss.n22674 0.003
R26846 vss.n22618 vss.n22606 0.003
R26847 vss.n22573 vss.n22572 0.003
R26848 vss.n22516 vss.n22504 0.003
R26849 vss.n22467 vss.n22466 0.003
R26850 vss.n22410 vss.n22398 0.003
R26851 vss.n22365 vss.n22364 0.003
R26852 vss.n22308 vss.n22296 0.003
R26853 vss.n22259 vss.n22258 0.003
R26854 vss.n22202 vss.n22190 0.003
R26855 vss.n22157 vss.n22156 0.003
R26856 vss.n22100 vss.n22088 0.003
R26857 vss.n158 vss.n156 0.003
R26858 vss.n171 vss.n169 0.003
R26859 vss.n186 vss.n184 0.003
R26860 vss.n262 vss.n260 0.003
R26861 vss.n420 vss.n418 0.003
R26862 vss.n501 vss.n499 0.003
R26863 vss.n665 vss.n663 0.003
R26864 vss.n745 vss.n743 0.003
R26865 vss.n909 vss.n907 0.003
R26866 vss.n990 vss.n988 0.003
R26867 vss.n1153 vss.n1151 0.003
R26868 vss.n1186 vss.n1170 0.003
R26869 vss.n1234 vss.n1232 0.003
R26870 vss.n23329 vss.n23327 0.003
R26871 vss.n23249 vss.n23247 0.003
R26872 vss.n23085 vss.n23083 0.003
R26873 vss.n23004 vss.n23002 0.003
R26874 vss.n22846 vss.n22844 0.003
R26875 vss.n14509 vss.n14499 0.003
R26876 vss.n13406 vss.n13397 0.003
R26877 vss.n9041 vss.n9040 0.003
R26878 vss.n9201 vss.n9200 0.003
R26879 vss.n9200 vss.t217 0.003
R26880 vss.n9199 vss.n9198 0.003
R26881 vss.t217 vss.n9199 0.003
R26882 vss.n17327 vss.n17317 0.002
R26883 vss.n17328 vss.n17327 0.002
R26884 vss.n20379 vss.n20378 0.002
R26885 vss.n6989 vss.n6988 0.002
R26886 vss.n9040 vss.n9038 0.002
R26887 vss.n21989 vss.n21987 0.002
R26888 vss.n3938 vss.n3936 0.002
R26889 vss.n15096 vss.n15062 0.002
R26890 vss.n18961 vss.n18960 0.002
R26891 vss.n18938 vss.n17686 0.002
R26892 vss.n18834 vss.n18833 0.002
R26893 vss.n18823 vss.n17795 0.002
R26894 vss.n17894 vss.n17882 0.002
R26895 vss.n18697 vss.n17896 0.002
R26896 vss.n18593 vss.n18592 0.002
R26897 vss.n18582 vss.n18008 0.002
R26898 vss.n18107 vss.n18095 0.002
R26899 vss.n18456 vss.n18109 0.002
R26900 vss.n18352 vss.n18351 0.002
R26901 vss.n18341 vss.n18221 0.002
R26902 vss.n20227 vss.n20226 0.002
R26903 vss.n20216 vss.n19095 0.002
R26904 vss.n20107 vss.n20106 0.002
R26905 vss.n20084 vss.n19193 0.002
R26906 vss.n19980 vss.n19979 0.002
R26907 vss.n19969 vss.n19302 0.002
R26908 vss.n19860 vss.n19859 0.002
R26909 vss.n19837 vss.n19399 0.002
R26910 vss.n19733 vss.n19732 0.002
R26911 vss.n19722 vss.n19509 0.002
R26912 vss.n19621 vss.n19587 0.002
R26913 vss.n20370 vss.n17581 0.002
R26914 vss.n20561 vss.n20547 0.002
R26915 vss.n20636 vss.n20625 0.002
R26916 vss.n20686 vss.n20684 0.002
R26917 vss.n20733 vss.n20731 0.002
R26918 vss.n20803 vss.n20801 0.002
R26919 vss.n20847 vss.n20845 0.002
R26920 vss.n20860 vss.n20849 0.002
R26921 vss.n21532 vss.n21520 0.002
R26922 vss.n21515 vss.n21514 0.002
R26923 vss.n21324 vss.n21312 0.002
R26924 vss.n21307 vss.n21306 0.002
R26925 vss.n21116 vss.n21104 0.002
R26926 vss.n21099 vss.n21098 0.002
R26927 vss.n20908 vss.n20896 0.002
R26928 vss.n22037 vss.n22036 0.002
R26929 vss.n22041 vss.n22039 0.002
R26930 vss.n22049 vss.n22048 0.002
R26931 vss.n21835 vss.n21828 0.002
R26932 vss.n21844 vss.n21842 0.002
R26933 vss.n21892 vss.n21889 0.002
R26934 vss.n22024 vss.n22022 0.002
R26935 vss.n22020 vss.n22018 0.002
R26936 vss.n21946 vss.n21922 0.002
R26937 vss.n21683 vss.n21680 0.002
R26938 vss.n21679 vss.n21665 0.002
R26939 vss.n21724 vss.n21723 0.002
R26940 vss.n21717 vss.n21715 0.002
R26941 vss.n21752 vss.n21709 0.002
R26942 vss.n21752 vss.n21707 0.002
R26943 vss.n21766 vss.n21762 0.002
R26944 vss.n21769 vss.n21768 0.002
R26945 vss.n9691 vss.n9690 0.002
R26946 vss.n9714 vss.n9696 0.002
R26947 vss.n10186 vss.n9676 0.002
R26948 vss.n10453 vss.n10452 0.002
R26949 vss.n15041 vss.n12778 0.002
R26950 vss.n15010 vss.n12824 0.002
R26951 vss.n14976 vss.n12903 0.002
R26952 vss.n12608 vss.n12486 0.002
R26953 vss.n12589 vss.n12534 0.002
R26954 vss.n12542 vss.n12541 0.002
R26955 vss.n12148 vss.n12106 0.002
R26956 vss.n12608 vss.n12607 0.002
R26957 vss.n12174 vss.n12164 0.002
R26958 vss.n12188 vss.n12178 0.002
R26959 vss.n12192 vss.n12190 0.002
R26960 vss.n12219 vss.n12217 0.002
R26961 vss.n12247 vss.n12245 0.002
R26962 vss.n12036 vss.n12025 0.002
R26963 vss.n12013 vss.n12011 0.002
R26964 vss.n11992 vss.n11982 0.002
R26965 vss.n11328 vss.n11326 0.002
R26966 vss.n11303 vss.n11301 0.002
R26967 vss.n11289 vss.n11287 0.002
R26968 vss.n11285 vss.n11275 0.002
R26969 vss.n11263 vss.n11261 0.002
R26970 vss.n11259 vss.n11249 0.002
R26971 vss.n11218 vss.n11217 0.002
R26972 vss.n11186 vss.n11184 0.002
R26973 vss.n11173 vss.n11171 0.002
R26974 vss.n11171 vss.n11169 0.002
R26975 vss.n11162 vss.n11152 0.002
R26976 vss.n11150 vss.n11148 0.002
R26977 vss.n12735 vss.n12734 0.002
R26978 vss.n12713 vss.n12712 0.002
R26979 vss.n12711 vss.n12710 0.002
R26980 vss.n12708 vss.n12696 0.002
R26981 vss.n12695 vss.n12694 0.002
R26982 vss.n12692 vss.n12680 0.002
R26983 vss.n12679 vss.n12678 0.002
R26984 vss.n12676 vss.n12675 0.002
R26985 vss.n12660 vss.n12659 0.002
R26986 vss.n12647 vss.n12646 0.002
R26987 vss.n14316 vss.n14314 0.002
R26988 vss.n14302 vss.n14300 0.002
R26989 vss.n13872 vss.n13870 0.002
R26990 vss.n13906 vss.n13904 0.002
R26991 vss.n13934 vss.n13932 0.002
R26992 vss.n14077 vss.n14056 0.002
R26993 vss.n14044 vss.n14043 0.002
R26994 vss.n11616 vss.n11614 0.002
R26995 vss.n11829 vss.n11827 0.002
R26996 vss.n11804 vss.n11802 0.002
R26997 vss.n11790 vss.n11788 0.002
R26998 vss.n11753 vss.n11751 0.002
R26999 vss.n11749 vss.n11739 0.002
R27000 vss.n11136 vss.n11134 0.002
R27001 vss.n14806 vss.n14804 0.002
R27002 vss.n14792 vss.n14790 0.002
R27003 vss.n14780 vss.n14778 0.002
R27004 vss.n14746 vss.n14745 0.002
R27005 vss.n14727 vss.n14726 0.002
R27006 vss.n14699 vss.n14686 0.002
R27007 vss.n14674 vss.n14672 0.002
R27008 vss.n14631 vss.n14621 0.002
R27009 vss.n14544 vss.n14542 0.002
R27010 vss.n14527 vss.n14525 0.002
R27011 vss.n14513 vss.n14511 0.002
R27012 vss.n14475 vss.n14473 0.002
R27013 vss.n14471 vss.n14461 0.002
R27014 vss.n14442 vss.n14441 0.002
R27015 vss.n14911 vss.n13249 0.002
R27016 vss.n14841 vss.n14840 0.002
R27017 vss.n14855 vss.n14852 0.002
R27018 vss.n15097 vss.n15096 0.002
R27019 vss.n3986 vss.n3985 0.002
R27020 vss.n3990 vss.n3988 0.002
R27021 vss.n3998 vss.n3997 0.002
R27022 vss.n3784 vss.n3777 0.002
R27023 vss.n3793 vss.n3791 0.002
R27024 vss.n3841 vss.n3838 0.002
R27025 vss.n3973 vss.n3971 0.002
R27026 vss.n3969 vss.n3967 0.002
R27027 vss.n3895 vss.n3871 0.002
R27028 vss.n3632 vss.n3629 0.002
R27029 vss.n3628 vss.n3614 0.002
R27030 vss.n3673 vss.n3672 0.002
R27031 vss.n3666 vss.n3664 0.002
R27032 vss.n3701 vss.n3658 0.002
R27033 vss.n3701 vss.n3656 0.002
R27034 vss.n3715 vss.n3711 0.002
R27035 vss.n3718 vss.n3717 0.002
R27036 vss.n5571 vss.n5570 0.002
R27037 vss.n5548 vss.n4296 0.002
R27038 vss.n5444 vss.n5443 0.002
R27039 vss.n5433 vss.n4405 0.002
R27040 vss.n4504 vss.n4492 0.002
R27041 vss.n5307 vss.n4506 0.002
R27042 vss.n5203 vss.n5202 0.002
R27043 vss.n5192 vss.n4618 0.002
R27044 vss.n4717 vss.n4705 0.002
R27045 vss.n5066 vss.n4719 0.002
R27046 vss.n4962 vss.n4961 0.002
R27047 vss.n4951 vss.n4831 0.002
R27048 vss.n6837 vss.n6836 0.002
R27049 vss.n6826 vss.n5705 0.002
R27050 vss.n6717 vss.n6716 0.002
R27051 vss.n6694 vss.n5803 0.002
R27052 vss.n6590 vss.n6589 0.002
R27053 vss.n6579 vss.n5912 0.002
R27054 vss.n6470 vss.n6469 0.002
R27055 vss.n6447 vss.n6009 0.002
R27056 vss.n6343 vss.n6342 0.002
R27057 vss.n6332 vss.n6119 0.002
R27058 vss.n6231 vss.n6197 0.002
R27059 vss.n6980 vss.n4191 0.002
R27060 vss.n7171 vss.n7157 0.002
R27061 vss.n7246 vss.n7235 0.002
R27062 vss.n7296 vss.n7294 0.002
R27063 vss.n7343 vss.n7341 0.002
R27064 vss.n7413 vss.n7411 0.002
R27065 vss.n7457 vss.n7455 0.002
R27066 vss.n7470 vss.n7459 0.002
R27067 vss.n8143 vss.n8131 0.002
R27068 vss.n8126 vss.n8125 0.002
R27069 vss.n7935 vss.n7923 0.002
R27070 vss.n7918 vss.n7917 0.002
R27071 vss.n7726 vss.n7714 0.002
R27072 vss.n7709 vss.n7708 0.002
R27073 vss.n7518 vss.n7506 0.002
R27074 vss.n8767 vss.n8755 0.002
R27075 vss.n8750 vss.n8749 0.002
R27076 vss.n8559 vss.n8547 0.002
R27077 vss.n8542 vss.n8541 0.002
R27078 vss.n8351 vss.n8339 0.002
R27079 vss.n8334 vss.n8333 0.002
R27080 vss.n1695 vss.n1693 0.002
R27081 vss.n1712 vss.n1710 0.002
R27082 vss.n1727 vss.n1725 0.002
R27083 vss.n1746 vss.n1743 0.002
R27084 vss.n1857 vss.n1846 0.002
R27085 vss.n1909 vss.n1907 0.002
R27086 vss.n1975 vss.n1973 0.002
R27087 vss.n2024 vss.n2022 0.002
R27088 vss.n2100 vss.n2088 0.002
R27089 vss.n2153 vss.n2151 0.002
R27090 vss.n2220 vss.n2218 0.002
R27091 vss.n2268 vss.n2266 0.002
R27092 vss.n2345 vss.n2333 0.002
R27093 vss.n2397 vss.n2395 0.002
R27094 vss.n2464 vss.n2462 0.002
R27095 vss.n2513 vss.n2511 0.002
R27096 vss.n2589 vss.n2577 0.002
R27097 vss.n2642 vss.n2640 0.002
R27098 vss.n2708 vss.n2706 0.002
R27099 vss.n2757 vss.n2755 0.002
R27100 vss.n2821 vss.n2819 0.002
R27101 vss.n2831 vss.n2821 0.002
R27102 vss.n2880 vss.n2878 0.002
R27103 vss.n2947 vss.n2945 0.002
R27104 vss.n2995 vss.n2993 0.002
R27105 vss.n3072 vss.n3060 0.002
R27106 vss.n3125 vss.n3123 0.002
R27107 vss.n3191 vss.n3189 0.002
R27108 vss.n3240 vss.n3238 0.002
R27109 vss.n3316 vss.n3304 0.002
R27110 vss.n3367 vss.n3365 0.002
R27111 vss.n3441 vss.n3439 0.002
R27112 vss.n15209 vss.n15195 0.002
R27113 vss.n15190 vss.n15189 0.002
R27114 vss.n15217 vss.n15216 0.002
R27115 vss.n15534 vss.n15532 0.002
R27116 vss.n15553 vss.n15551 0.002
R27117 vss.n15770 vss.n15768 0.002
R27118 vss.n15305 vss.n15303 0.002
R27119 vss.n15344 vss.n15342 0.002
R27120 vss.n15819 vss.n15816 0.002
R27121 vss.n16060 vss.n16059 0.002
R27122 vss.n16088 vss.n16076 0.002
R27123 vss.n16481 vss.n16479 0.002
R27124 vss.n16500 vss.n16498 0.002
R27125 vss.n16823 vss.n16822 0.002
R27126 vss.n17014 vss.n17013 0.002
R27127 vss.n17031 vss.n17030 0.002
R27128 vss.n17250 vss.n17249 0.002
R27129 vss.n17317 vss.n16266 0.002
R27130 vss.n22604 vss.n22592 0.002
R27131 vss.n22587 vss.n22586 0.002
R27132 vss.n22396 vss.n22384 0.002
R27133 vss.n22379 vss.n22378 0.002
R27134 vss.n22188 vss.n22176 0.002
R27135 vss.n22171 vss.n22170 0.002
R27136 vss.n156 vss.n154 0.002
R27137 vss.n173 vss.n171 0.002
R27138 vss.n188 vss.n186 0.002
R27139 vss.n207 vss.n204 0.002
R27140 vss.n318 vss.n307 0.002
R27141 vss.n370 vss.n368 0.002
R27142 vss.n436 vss.n434 0.002
R27143 vss.n485 vss.n483 0.002
R27144 vss.n561 vss.n549 0.002
R27145 vss.n614 vss.n612 0.002
R27146 vss.n681 vss.n679 0.002
R27147 vss.n729 vss.n727 0.002
R27148 vss.n806 vss.n794 0.002
R27149 vss.n858 vss.n856 0.002
R27150 vss.n925 vss.n923 0.002
R27151 vss.n974 vss.n972 0.002
R27152 vss.n1050 vss.n1038 0.002
R27153 vss.n1103 vss.n1101 0.002
R27154 vss.n1169 vss.n1167 0.002
R27155 vss.n1218 vss.n1216 0.002
R27156 vss.n1283 vss.n1281 0.002
R27157 vss.n1295 vss.n1283 0.002
R27158 vss.n23389 vss.n23377 0.002
R27159 vss.n23313 vss.n23311 0.002
R27160 vss.n23265 vss.n23263 0.002
R27161 vss.n23198 vss.n23196 0.002
R27162 vss.n23145 vss.n23133 0.002
R27163 vss.n23069 vss.n23067 0.002
R27164 vss.n23020 vss.n23018 0.002
R27165 vss.n22954 vss.n22952 0.002
R27166 vss.n22902 vss.n22891 0.002
R27167 vss.n1416 vss.n1414 0.002
R27168 vss.n22842 vss.n22829 0.002
R27169 vss.n22824 vss.n22823 0.002
R27170 vss.n10263 vss.n10262 0.002
R27171 vss.n10425 vss.n10423 0.002
R27172 vss.n21821 vss.n21806 0.001
R27173 vss.n21821 vss.n21820 0.001
R27174 vss.n3770 vss.n3755 0.001
R27175 vss.n3770 vss.n3769 0.001
R27176 vss.n10423 vss.n10422 0.001
R27177 vss.n10394 vss.n10393 0.001
R27178 vss.n9146 vss.n9145 0.001
R27179 vss.n14040 vss.n14039 0.001
R27180 vss.n14499 vss.n14498 0.001
R27181 vss.n14668 vss.n14667 0.001
R27182 vss.n17549 vss.n17548 0.001
R27183 vss.n4159 vss.n4158 0.001
R27184 vss.n10225 vss.n10222 0.001
R27185 vss.n19023 vss.n19022 0.001
R27186 vss.n19006 vss.n19005 0.001
R27187 vss.n18891 vss.n17732 0.001
R27188 vss.n18880 vss.n17733 0.001
R27189 vss.n17836 vss.n17833 0.001
R27190 vss.n18765 vss.n17843 0.001
R27191 vss.n18650 vss.n17945 0.001
R27192 vss.n18639 vss.n17946 0.001
R27193 vss.n18049 vss.n18046 0.001
R27194 vss.n18524 vss.n18056 0.001
R27195 vss.n18409 vss.n18158 0.001
R27196 vss.n18398 vss.n18159 0.001
R27197 vss.n18262 vss.n18259 0.001
R27198 vss.n18283 vss.n18269 0.001
R27199 vss.n20289 vss.n20288 0.001
R27200 vss.n19046 vss.n19044 0.001
R27201 vss.n19136 vss.n19133 0.001
R27202 vss.n20152 vss.n20151 0.001
R27203 vss.n20037 vss.n19239 0.001
R27204 vss.n20026 vss.n19240 0.001
R27205 vss.n19343 vss.n19340 0.001
R27206 vss.n19905 vss.n19904 0.001
R27207 vss.n19790 vss.n19446 0.001
R27208 vss.n19779 vss.n19447 0.001
R27209 vss.n19550 vss.n19547 0.001
R27210 vss.n19658 vss.n19657 0.001
R27211 vss.n20374 vss.n17577 0.001
R27212 vss.n17537 vss.n17535 0.001
R27213 vss.n17542 vss.n17540 0.001
R27214 vss.n20538 vss.n20536 0.001
R27215 vss.n20546 vss.n20544 0.001
R27216 vss.n17492 vss.n17490 0.001
R27217 vss.n17497 vss.n17495 0.001
R27218 vss.n20651 vss.n20640 0.001
R27219 vss.n20671 vss.n20669 0.001
R27220 vss.n20748 vss.n20746 0.001
R27221 vss.n20787 vss.n20785 0.001
R27222 vss.n21430 vss.n21416 0.001
R27223 vss.n21411 vss.n21410 0.001
R27224 vss.n21222 vss.n21208 0.001
R27225 vss.n21203 vss.n21202 0.001
R27226 vss.n21014 vss.n21000 0.001
R27227 vss.n20995 vss.n20994 0.001
R27228 vss.n21902 vss.n21901 0.001
R27229 vss.n21919 vss.n21918 0.001
R27230 vss.n9661 vss.n9658 0.001
R27231 vss.n10228 vss.n9674 0.001
R27232 vss.n10445 vss.n10443 0.001
R27233 vss.n8930 vss.n8929 0.001
R27234 vss.n8967 vss.n8966 0.001
R27235 vss.n8979 vss.n8978 0.001
R27236 vss.n9000 vss.n8999 0.001
R27237 vss.n9030 vss.n9029 0.001
R27238 vss.n9061 vss.n9060 0.001
R27239 vss.n9092 vss.n9091 0.001
R27240 vss.n9112 vss.n9111 0.001
R27241 vss.n9141 vss.n9140 0.001
R27242 vss.n13173 vss.n13172 0.001
R27243 vss.n12775 vss.n12770 0.001
R27244 vss.n12901 vss.n12898 0.001
R27245 vss.n14976 vss.n12923 0.001
R27246 vss.n12637 vss.n12636 0.001
R27247 vss.n12608 vss.n12510 0.001
R27248 vss.n12632 vss.n12630 0.001
R27249 vss.n12630 vss.n12621 0.001
R27250 vss.n12621 vss.n12619 0.001
R27251 vss.n12619 vss.n12609 0.001
R27252 vss.n12607 vss.n12605 0.001
R27253 vss.n12605 vss.n12604 0.001
R27254 vss.n12604 vss.n12602 0.001
R27255 vss.n12602 vss.n12593 0.001
R27256 vss.n12158 vss.n12150 0.001
R27257 vss.n12160 vss.n12158 0.001
R27258 vss.n12162 vss.n12160 0.001
R27259 vss.n12164 vss.n12162 0.001
R27260 vss.n12178 vss.n12176 0.001
R27261 vss.n12202 vss.n12192 0.001
R27262 vss.n12206 vss.n12204 0.001
R27263 vss.n12215 vss.n12206 0.001
R27264 vss.n12217 vss.n12215 0.001
R27265 vss.n12229 vss.n12219 0.001
R27266 vss.n12240 vss.n12230 0.001
R27267 vss.n12242 vss.n12240 0.001
R27268 vss.n12301 vss.n12267 0.001
R27269 vss.n12023 vss.n12013 0.001
R27270 vss.n12011 vss.n12009 0.001
R27271 vss.n12008 vss.n12007 0.001
R27272 vss.n12007 vss.n11996 0.001
R27273 vss.n11995 vss.n11994 0.001
R27274 vss.n11994 vss.n11993 0.001
R27275 vss.n11982 vss.n11980 0.001
R27276 vss.n11967 vss.n11966 0.001
R27277 vss.n11966 vss.n11956 0.001
R27278 vss.n11955 vss.n11954 0.001
R27279 vss.n11954 vss.n11953 0.001
R27280 vss.n11330 vss.n11328 0.001
R27281 vss.n11305 vss.n11303 0.001
R27282 vss.n11287 vss.n11285 0.001
R27283 vss.n11275 vss.n11274 0.001
R27284 vss.n11274 vss.n11264 0.001
R27285 vss.n11261 vss.n11259 0.001
R27286 vss.n11249 vss.n11248 0.001
R27287 vss.n11248 vss.n11239 0.001
R27288 vss.n11239 vss.n11226 0.001
R27289 vss.n11217 vss.n11215 0.001
R27290 vss.n11215 vss.n11213 0.001
R27291 vss.n11213 vss.n11204 0.001
R27292 vss.n11203 vss.n11202 0.001
R27293 vss.n11202 vss.n11201 0.001
R27294 vss.n11201 vss.n11200 0.001
R27295 vss.n11199 vss.n11189 0.001
R27296 vss.n11189 vss.n11187 0.001
R27297 vss.n11187 vss.n11186 0.001
R27298 vss.n11183 vss.n11173 0.001
R27299 vss.n11152 vss.n11150 0.001
R27300 vss.n14164 vss.n14163 0.001
R27301 vss.n14163 vss.n14153 0.001
R27302 vss.n14153 vss.n14151 0.001
R27303 vss.n14151 vss.n14143 0.001
R27304 vss.n14141 vss.n14139 0.001
R27305 vss.n14139 vss.n14122 0.001
R27306 vss.n14122 vss.n14120 0.001
R27307 vss.n14120 vss.n14110 0.001
R27308 vss.n14109 vss.n14107 0.001
R27309 vss.n14107 vss.n14106 0.001
R27310 vss.n14106 vss.n14104 0.001
R27311 vss.n14104 vss.n14095 0.001
R27312 vss.n13755 vss.n13754 0.001
R27313 vss.n13754 vss.n13745 0.001
R27314 vss.n13745 vss.n13743 0.001
R27315 vss.n13743 vss.n13742 0.001
R27316 vss.n13740 vss.n13739 0.001
R27317 vss.n13739 vss.n13729 0.001
R27318 vss.n13729 vss.n13727 0.001
R27319 vss.n13727 vss.n13726 0.001
R27320 vss.n11424 vss.n11407 0.001
R27321 vss.n11426 vss.n11424 0.001
R27322 vss.n11436 vss.n11426 0.001
R27323 vss.n11437 vss.n11436 0.001
R27324 vss.n11440 vss.n11439 0.001
R27325 vss.n11442 vss.n11440 0.001
R27326 vss.n11451 vss.n11442 0.001
R27327 vss.n11452 vss.n11451 0.001
R27328 vss.n11860 vss.n11851 0.001
R27329 vss.n11862 vss.n11860 0.001
R27330 vss.n11863 vss.n11862 0.001
R27331 vss.n11865 vss.n11863 0.001
R27332 vss.n11876 vss.n11866 0.001
R27333 vss.n11878 vss.n11876 0.001
R27334 vss.n11879 vss.n11878 0.001
R27335 vss.n11881 vss.n11879 0.001
R27336 vss.n11900 vss.n11883 0.001
R27337 vss.n11902 vss.n11900 0.001
R27338 vss.n11912 vss.n11902 0.001
R27339 vss.n11913 vss.n11912 0.001
R27340 vss.n13467 vss.n13465 0.001
R27341 vss.n13465 vss.n13464 0.001
R27342 vss.n13464 vss.n13462 0.001
R27343 vss.n13462 vss.n13453 0.001
R27344 vss.n14975 vss.n13111 0.001
R27345 vss.n13094 vss.n13093 0.001
R27346 vss.n13093 vss.n13084 0.001
R27347 vss.n13084 vss.n13082 0.001
R27348 vss.n13082 vss.n13081 0.001
R27349 vss.n13079 vss.n13078 0.001
R27350 vss.n13078 vss.n13068 0.001
R27351 vss.n13068 vss.n13066 0.001
R27352 vss.n13066 vss.n13065 0.001
R27353 vss.n10619 vss.n10601 0.001
R27354 vss.n10621 vss.n10619 0.001
R27355 vss.n10631 vss.n10621 0.001
R27356 vss.n10632 vss.n10631 0.001
R27357 vss.n10635 vss.n10634 0.001
R27358 vss.n10637 vss.n10635 0.001
R27359 vss.n10646 vss.n10637 0.001
R27360 vss.n10647 vss.n10646 0.001
R27361 vss.n12710 vss.n10725 0.001
R27362 vss.n12316 vss.n12315 0.001
R27363 vss.n12315 vss.n12306 0.001
R27364 vss.n12306 vss.n12304 0.001
R27365 vss.n12304 vss.n12303 0.001
R27366 vss.n12732 vss.n12731 0.001
R27367 vss.n12731 vss.n12730 0.001
R27368 vss.n12728 vss.n12727 0.001
R27369 vss.n12727 vss.n12719 0.001
R27370 vss.n12709 vss.n12708 0.001
R27371 vss.n12693 vss.n12692 0.001
R27372 vss.n12678 vss.n12677 0.001
R27373 vss.n12675 vss.n12663 0.001
R27374 vss.n12659 vss.n12647 0.001
R27375 vss.n12646 vss.n12645 0.001
R27376 vss.n12645 vss.n12644 0.001
R27377 vss.n13814 vss.n13813 0.001
R27378 vss.n14364 vss.n14341 0.001
R27379 vss.n14330 vss.n14329 0.001
R27380 vss.n14329 vss.n14320 0.001
R27381 vss.n14320 vss.n14318 0.001
R27382 vss.n14318 vss.n14316 0.001
R27383 vss.n14304 vss.n14302 0.001
R27384 vss.n13882 vss.n13872 0.001
R27385 vss.n13893 vss.n13884 0.001
R27386 vss.n13902 vss.n13893 0.001
R27387 vss.n13904 vss.n13902 0.001
R27388 vss.n13916 vss.n13906 0.001
R27389 vss.n13927 vss.n13917 0.001
R27390 vss.n13929 vss.n13927 0.001
R27391 vss.n14078 vss.n13953 0.001
R27392 vss.n14054 vss.n14044 0.001
R27393 vss.n14043 vss.n14041 0.001
R27394 vss.n14029 vss.n14028 0.001
R27395 vss.n14027 vss.n14026 0.001
R27396 vss.n14026 vss.n14025 0.001
R27397 vss.n11618 vss.n11616 0.001
R27398 vss.n11641 vss.n11639 0.001
R27399 vss.n11642 vss.n11641 0.001
R27400 vss.n11653 vss.n11643 0.001
R27401 vss.n11654 vss.n11653 0.001
R27402 vss.n11831 vss.n11829 0.001
R27403 vss.n11806 vss.n11804 0.001
R27404 vss.n11788 vss.n11786 0.001
R27405 vss.n11767 vss.n11754 0.001
R27406 vss.n11751 vss.n11749 0.001
R27407 vss.n11739 vss.n11738 0.001
R27408 vss.n11738 vss.n11729 0.001
R27409 vss.n11729 vss.n11727 0.001
R27410 vss.n11138 vss.n11136 0.001
R27411 vss.n11146 vss.n11138 0.001
R27412 vss.n11147 vss.n11146 0.001
R27413 vss.n13318 vss.n13310 0.001
R27414 vss.n13320 vss.n13318 0.001
R27415 vss.n14807 vss.n13320 0.001
R27416 vss.n14807 vss.n14806 0.001
R27417 vss.n14794 vss.n14792 0.001
R27418 vss.n14778 vss.n14776 0.001
R27419 vss.n14766 vss.n14764 0.001
R27420 vss.n14764 vss.n14755 0.001
R27421 vss.n14755 vss.n14746 0.001
R27422 vss.n14745 vss.n14743 0.001
R27423 vss.n14733 vss.n14732 0.001
R27424 vss.n14732 vss.n14731 0.001
R27425 vss.n14702 vss.n14700 0.001
R27426 vss.n14684 vss.n14674 0.001
R27427 vss.n14672 vss.n14670 0.001
R27428 vss.n14667 vss.n14646 0.001
R27429 vss.n14645 vss.n14644 0.001
R27430 vss.n14644 vss.n14632 0.001
R27431 vss.n14621 vss.n14619 0.001
R27432 vss.n14606 vss.n14605 0.001
R27433 vss.n14605 vss.n14604 0.001
R27434 vss.n14603 vss.n14602 0.001
R27435 vss.n14602 vss.n14601 0.001
R27436 vss.n14546 vss.n14544 0.001
R27437 vss.n14529 vss.n14527 0.001
R27438 vss.n14511 vss.n14509 0.001
R27439 vss.n14498 vss.n14476 0.001
R27440 vss.n14473 vss.n14471 0.001
R27441 vss.n14461 vss.n14460 0.001
R27442 vss.n14460 vss.n14451 0.001
R27443 vss.n14451 vss.n14450 0.001
R27444 vss.n14441 vss.n14439 0.001
R27445 vss.n14439 vss.n14430 0.001
R27446 vss.n14430 vss.n14422 0.001
R27447 vss.n13244 vss.n13235 0.001
R27448 vss.n13246 vss.n13244 0.001
R27449 vss.n13247 vss.n13246 0.001
R27450 vss.n13249 vss.n13247 0.001
R27451 vss.n14922 vss.n14912 0.001
R27452 vss.n14924 vss.n14922 0.001
R27453 vss.n14925 vss.n14924 0.001
R27454 vss.n14927 vss.n14925 0.001
R27455 vss.n14938 vss.n14929 0.001
R27456 vss.n14940 vss.n14938 0.001
R27457 vss.n14950 vss.n14940 0.001
R27458 vss.n14951 vss.n14950 0.001
R27459 vss.n14954 vss.n14953 0.001
R27460 vss.n14956 vss.n14954 0.001
R27461 vss.n14965 vss.n14956 0.001
R27462 vss.n14966 vss.n14965 0.001
R27463 vss.n15006 vss.n14976 0.001
R27464 vss.n15008 vss.n15007 0.001
R27465 vss.n15019 vss.n15010 0.001
R27466 vss.n15021 vss.n15019 0.001
R27467 vss.n15022 vss.n15021 0.001
R27468 vss.n15024 vss.n15022 0.001
R27469 vss.n15035 vss.n15025 0.001
R27470 vss.n15037 vss.n15035 0.001
R27471 vss.n15038 vss.n15037 0.001
R27472 vss.n15040 vss.n15038 0.001
R27473 vss.n12896 vss.n12895 0.001
R27474 vss.n3851 vss.n3850 0.001
R27475 vss.n3868 vss.n3867 0.001
R27476 vss.n5633 vss.n5632 0.001
R27477 vss.n5616 vss.n5615 0.001
R27478 vss.n5501 vss.n4342 0.001
R27479 vss.n5490 vss.n4343 0.001
R27480 vss.n4446 vss.n4443 0.001
R27481 vss.n5375 vss.n4453 0.001
R27482 vss.n5260 vss.n4555 0.001
R27483 vss.n5249 vss.n4556 0.001
R27484 vss.n4659 vss.n4656 0.001
R27485 vss.n5134 vss.n4666 0.001
R27486 vss.n5019 vss.n4768 0.001
R27487 vss.n5008 vss.n4769 0.001
R27488 vss.n4872 vss.n4869 0.001
R27489 vss.n4893 vss.n4879 0.001
R27490 vss.n6899 vss.n6898 0.001
R27491 vss.n5656 vss.n5654 0.001
R27492 vss.n5746 vss.n5743 0.001
R27493 vss.n6762 vss.n6761 0.001
R27494 vss.n6647 vss.n5849 0.001
R27495 vss.n6636 vss.n5850 0.001
R27496 vss.n5953 vss.n5950 0.001
R27497 vss.n6515 vss.n6514 0.001
R27498 vss.n6400 vss.n6056 0.001
R27499 vss.n6389 vss.n6057 0.001
R27500 vss.n6160 vss.n6157 0.001
R27501 vss.n6268 vss.n6267 0.001
R27502 vss.n6984 vss.n4187 0.001
R27503 vss.n4147 vss.n4145 0.001
R27504 vss.n4152 vss.n4150 0.001
R27505 vss.n7148 vss.n7146 0.001
R27506 vss.n7156 vss.n7154 0.001
R27507 vss.n4102 vss.n4100 0.001
R27508 vss.n4107 vss.n4105 0.001
R27509 vss.n7261 vss.n7250 0.001
R27510 vss.n7281 vss.n7279 0.001
R27511 vss.n7358 vss.n7356 0.001
R27512 vss.n7397 vss.n7395 0.001
R27513 vss.n8041 vss.n8027 0.001
R27514 vss.n8022 vss.n8021 0.001
R27515 vss.n7832 vss.n7818 0.001
R27516 vss.n7813 vss.n7812 0.001
R27517 vss.n7624 vss.n7610 0.001
R27518 vss.n7605 vss.n7604 0.001
R27519 vss.n8873 vss.n8859 0.001
R27520 vss.n8854 vss.n8853 0.001
R27521 vss.n8665 vss.n8651 0.001
R27522 vss.n8646 vss.n8645 0.001
R27523 vss.n8457 vss.n8443 0.001
R27524 vss.n8438 vss.n8437 0.001
R27525 vss.n1742 vss.n1740 0.001
R27526 vss.n1784 vss.n1782 0.001
R27527 vss.n1872 vss.n1861 0.001
R27528 vss.n1893 vss.n1891 0.001
R27529 vss.n1995 vss.n1993 0.001
R27530 vss.n2004 vss.n2002 0.001
R27531 vss.n2117 vss.n2105 0.001
R27532 vss.n2137 vss.n2135 0.001
R27533 vss.n2200 vss.n2188 0.001
R27534 vss.n2240 vss.n2238 0.001
R27535 vss.n2248 vss.n2246 0.001
R27536 vss.n2361 vss.n2349 0.001
R27537 vss.n2381 vss.n2379 0.001
R27538 vss.n2484 vss.n2482 0.001
R27539 vss.n2492 vss.n2490 0.001
R27540 vss.n2605 vss.n2593 0.001
R27541 vss.n2626 vss.n2624 0.001
R27542 vss.n2729 vss.n2727 0.001
R27543 vss.n2737 vss.n2735 0.001
R27544 vss.n2834 vss.n2833 0.001
R27545 vss.n2864 vss.n2862 0.001
R27546 vss.n2967 vss.n2965 0.001
R27547 vss.n2975 vss.n2973 0.001
R27548 vss.n3024 vss.n3012 0.001
R27549 vss.n3088 vss.n3076 0.001
R27550 vss.n3108 vss.n3106 0.001
R27551 vss.n3211 vss.n3209 0.001
R27552 vss.n3220 vss.n3218 0.001
R27553 vss.n3332 vss.n3320 0.001
R27554 vss.n3352 vss.n3350 0.001
R27555 vss.n3446 vss.n3444 0.001
R27556 vss.n3435 vss.n3433 0.001
R27557 vss.n15174 vss.n15173 0.001
R27558 vss.n15172 vss.n15170 0.001
R27559 vss.n15170 vss.n15168 0.001
R27560 vss.n15157 vss.n15156 0.001
R27561 vss.n15422 vss.n15415 0.001
R27562 vss.n15434 vss.n15432 0.001
R27563 vss.n15658 vss.n15651 0.001
R27564 vss.n15670 vss.n15668 0.001
R27565 vss.n15330 vss.n15328 0.001
R27566 vss.n15357 vss.n15356 0.001
R27567 vss.n15948 vss.n15947 0.001
R27568 vss.n15961 vss.n15949 0.001
R27569 vss.n16184 vss.n16183 0.001
R27570 vss.n16197 vss.n16185 0.001
R27571 vss.n16293 vss.n16286 0.001
R27572 vss.n16369 vss.n16362 0.001
R27573 vss.n16381 vss.n16379 0.001
R27574 vss.n16605 vss.n16598 0.001
R27575 vss.n16617 vss.n16615 0.001
R27576 vss.n16685 vss.n16684 0.001
R27577 vss.n16809 vss.n16808 0.001
R27578 vss.n16902 vss.n16893 0.001
R27579 vss.n16915 vss.n16914 0.001
R27580 vss.n17138 vss.n17129 0.001
R27581 vss.n17151 vss.n17150 0.001
R27582 vss.n16253 vss.n16252 0.001
R27583 vss.n22710 vss.n22696 0.001
R27584 vss.n22691 vss.n22690 0.001
R27585 vss.n22502 vss.n22488 0.001
R27586 vss.n22483 vss.n22482 0.001
R27587 vss.n22294 vss.n22280 0.001
R27588 vss.n22275 vss.n22274 0.001
R27589 vss.n203 vss.n201 0.001
R27590 vss.n245 vss.n243 0.001
R27591 vss.n333 vss.n322 0.001
R27592 vss.n354 vss.n352 0.001
R27593 vss.n456 vss.n454 0.001
R27594 vss.n465 vss.n463 0.001
R27595 vss.n578 vss.n566 0.001
R27596 vss.n598 vss.n596 0.001
R27597 vss.n661 vss.n649 0.001
R27598 vss.n701 vss.n699 0.001
R27599 vss.n709 vss.n707 0.001
R27600 vss.n822 vss.n810 0.001
R27601 vss.n842 vss.n840 0.001
R27602 vss.n945 vss.n943 0.001
R27603 vss.n953 vss.n951 0.001
R27604 vss.n1066 vss.n1054 0.001
R27605 vss.n1087 vss.n1085 0.001
R27606 vss.n1190 vss.n1188 0.001
R27607 vss.n1198 vss.n1196 0.001
R27608 vss.n1311 vss.n1299 0.001
R27609 vss.n23405 vss.n23393 0.001
R27610 vss.n23293 vss.n23291 0.001
R27611 vss.n23285 vss.n23283 0.001
R27612 vss.n23245 vss.n23244 0.001
R27613 vss.n23182 vss.n23180 0.001
R27614 vss.n23162 vss.n23150 0.001
R27615 vss.n23049 vss.n23047 0.001
R27616 vss.n23040 vss.n23038 0.001
R27617 vss.n22938 vss.n22936 0.001
R27618 vss.n22917 vss.n22906 0.001
R27619 vss.n1421 vss.n1419 0.001
R27620 vss.n1410 vss.n1408 0.001
R27621 vss.n22808 vss.n22807 0.001
R27622 vss.n22806 vss.n22804 0.001
R27623 vss.n22804 vss.n22802 0.001
R27624 vss.n22791 vss.n22790 0.001
R27625 vss.n12280 vss.n12270 0.001
R27626 vss.n13479 vss.n13470 0.001
R27627 vss.n10721 vss.n10720 0.001
R27628 vss.n13011 vss.n13010 0.001
R27629 vss.n12380 vss.n12379 0.001
R27630 vss.n11540 vss.n11539 0.001
R27631 vss.n10228 vss.n10225 0.001
R27632 vss.n9170 vss.n9169 0.001
R27633 vss.n9162 vss.n9161 0.001
R27634 vss.n10235 vss.n10234 0.001
R27635 vss.n10261 vss.n10260 0.001
R27636 vss.n10280 vss.n10279 0.001
R27637 vss.n10303 vss.n10302 0.001
R27638 vss.n10346 vss.n10345 0.001
R27639 vss.n10362 vss.n10361 0.001
R27640 vss.n10393 vss.n10392 0.001
R27641 vss.n10422 vss.n10421 0.001
R27642 vss.n8929 vss.n8928 0.001
R27643 vss.n8966 vss.n8965 0.001
R27644 vss.n8978 vss.n8977 0.001
R27645 vss.n9007 vss.n9006 0.001
R27646 vss.n9038 vss.n9037 0.001
R27647 vss.n9069 vss.n9068 0.001
R27648 vss.n9117 vss.n9116 0.001
R27649 vss.n9145 vss.n9144 0.001
R27650 vss.n9169 vss.n9168 0.001
R27651 vss.n9173 vss.n9172 0.001
R27652 vss.n20374 vss.n17578 0.001
R27653 vss.n6984 vss.n4188 0.001
R27654 vss.n12662 vss.n12661 0.001
R27655 vss.n14365 vss.n14364 0.001
R27656 vss.n14669 vss.n14668 0.001
R27657 vss.n14039 vss.n14029 0.001
R27658 vss.n11776 vss.n11767 0.001
R27659 vss.n10221 vss.n10220 0.001
R27660 vss.n15062 vss.n15061 0.001
R27661 vss.n9174 vss.n9173 0.001
R27662 vss.n10236 vss.n10235 0.001
R27663 vss.n10281 vss.n10280 0.001
R27664 vss.t166 vss.n14019 0.001
R27665 vss.t174 vss.n11229 0.001
R27666 vss.t110 vss.n10863 0.001
R27667 vss.n10865 vss.n10864 0.001
R27668 vss.n10864 vss.t110 0.001
R27669 vss.t147 vss.n12782 0.001
R27670 vss.t168 vss.n13206 0.001
R27671 vss.n12782 vss.n12781 0.001
R27672 vss.n13206 vss.n13205 0.001
R27673 vss.t176 vss.n13059 0.001
R27674 vss.n13059 vss.n13058 0.001
R27675 vss.n10863 vss.n10862 0.001
R27676 vss.n14019 vss.n14018 0.001
R27677 vss.n11229 vss.n11228 0.001
R27678 vss.n15122 vss.n10456 0.001
R27679 vss.n7 vss.n4235 806.541
R27680 vss.n5 vss.n4227 806.541
R27681 vss.n3 vss.n17625 806.541
R27682 vss.n1 vss.n17617 806.541
R27683 bandgapmd_0.otam_1.nmosrm_0.outn.n49 bandgapmd_0.otam_1.nmosrm_0.outn.n48 99.753
R27684 bandgapmd_0.otam_1.nmosrm_0.outn.n142 bandgapmd_0.otam_1.nmosrm_0.outn.n141 99.753
R27685 bandgapmd_0.otam_1.nmosrm_0.outn.n78 bandgapmd_0.otam_1.nmosrm_0.outn.n77 98.624
R27686 bandgapmd_0.otam_1.nmosrm_0.outn.n36 bandgapmd_0.otam_1.nmosrm_0.outn.n34 98.248
R27687 bandgapmd_0.otam_1.nmosrm_0.outn.n127 bandgapmd_0.otam_1.nmosrm_0.outn.n125 98.248
R27688 bandgapmd_0.otam_1.nmosrm_0.outn.n97 bandgapmd_0.otam_1.nmosrm_0.outn.n95 95.953
R27689 bandgapmd_0.otam_1.nmosrm_0.outn.n48 bandgapmd_0.otam_1.nmosrm_0.outn.t7 16.53
R27690 bandgapmd_0.otam_1.nmosrm_0.outn.n48 bandgapmd_0.otam_1.nmosrm_0.outn.t4 16.53
R27691 bandgapmd_0.otam_1.nmosrm_0.outn.n34 bandgapmd_0.otam_1.nmosrm_0.outn.t10 16.53
R27692 bandgapmd_0.otam_1.nmosrm_0.outn.n34 bandgapmd_0.otam_1.nmosrm_0.outn.t12 16.53
R27693 bandgapmd_0.otam_1.nmosrm_0.outn.n59 bandgapmd_0.otam_1.nmosrm_0.outn.t6 16.53
R27694 bandgapmd_0.otam_1.nmosrm_0.outn.n59 bandgapmd_0.otam_1.nmosrm_0.outn.t8 16.53
R27695 bandgapmd_0.otam_1.nmosrm_0.outn.n77 bandgapmd_0.otam_1.nmosrm_0.outn.t15 16.53
R27696 bandgapmd_0.otam_1.nmosrm_0.outn.n77 bandgapmd_0.otam_1.nmosrm_0.outn.t1 16.53
R27697 bandgapmd_0.otam_1.nmosrm_0.outn.n95 bandgapmd_0.otam_1.nmosrm_0.outn.t2 16.53
R27698 bandgapmd_0.otam_1.nmosrm_0.outn.n95 bandgapmd_0.otam_1.nmosrm_0.outn.t9 16.53
R27699 bandgapmd_0.otam_1.nmosrm_0.outn.n102 bandgapmd_0.otam_1.nmosrm_0.outn.t0 16.53
R27700 bandgapmd_0.otam_1.nmosrm_0.outn.n102 bandgapmd_0.otam_1.nmosrm_0.outn.t13 16.53
R27701 bandgapmd_0.otam_1.nmosrm_0.outn.n141 bandgapmd_0.otam_1.nmosrm_0.outn.t3 16.53
R27702 bandgapmd_0.otam_1.nmosrm_0.outn.n141 bandgapmd_0.otam_1.nmosrm_0.outn.t5 16.53
R27703 bandgapmd_0.otam_1.nmosrm_0.outn.n125 bandgapmd_0.otam_1.nmosrm_0.outn.t11 16.53
R27704 bandgapmd_0.otam_1.nmosrm_0.outn.n125 bandgapmd_0.otam_1.nmosrm_0.outn.t14 16.53
R27705 bandgapmd_0.otam_1.nmosrm_0.outn.n58 bandgapmd_0.otam_1.nmosrm_0.outn.n57 13.176
R27706 bandgapmd_0.otam_1.nmosrm_0.outn.n107 bandgapmd_0.otam_1.nmosrm_0.outn.n105 12.423
R27707 bandgapmd_0.otam_1.nmosrm_0.outn.n28 bandgapmd_0.otam_1.nmosrm_0.outn.n26 10.541
R27708 bandgapmd_0.otam_1.nmosrm_0.outn.n119 bandgapmd_0.otam_1.nmosrm_0.outn.n117 10.541
R27709 bandgapmd_0.otam_1.nmosrm_0.outn.n70 bandgapmd_0.otam_1.nmosrm_0.outn.n68 10.164
R27710 bandgapmd_0.otam_1.nmosrm_0.outn.n14 bandgapmd_0.otam_1.nmosrm_0.outn.n156 9.321
R27711 bandgapmd_0.otam_1.nmosrm_0.outn.n24 bandgapmd_0.otam_1.nmosrm_0.outn.n31 9.3
R27712 bandgapmd_0.otam_1.nmosrm_0.outn.n66 bandgapmd_0.otam_1.nmosrm_0.outn.n73 9.3
R27713 bandgapmd_0.otam_1.nmosrm_0.outn.n21 bandgapmd_0.otam_1.nmosrm_0.outn.n104 9.3
R27714 bandgapmd_0.otam_1.nmosrm_0.outn.n21 bandgapmd_0.otam_1.nmosrm_0.outn.n103 9.3
R27715 bandgapmd_0.otam_1.nmosrm_0.outn.n115 bandgapmd_0.otam_1.nmosrm_0.outn.n122 9.3
R27716 bandgapmd_0.otam_1.nmosrm_0.outn.n155 bandgapmd_0.otam_1.nmosrm_0.outn.n154 9.3
R27717 bandgapmd_0.otam_1.nmosrm_0.outn.n15 bandgapmd_0.otam_1.nmosrm_0.outn.n158 9.3
R27718 bandgapmd_0.otam_1.nmosrm_0.outn.n15 bandgapmd_0.otam_1.nmosrm_0.outn.n157 9.3
R27719 bandgapmd_0.otam_1.nmosrm_0.outn.n60 bandgapmd_0.otam_1.nmosrm_0.outn.n59 8.5
R27720 bandgapmd_0.otam_1.nmosrm_0.outn.n103 bandgapmd_0.otam_1.nmosrm_0.outn.n102 8.5
R27721 bandgapmd_0.otam_1.nmosrm_0.outn.n160 bandgapmd_0.otam_1.nmosrm_0.outn.t18 8.265
R27722 bandgapmd_0.otam_1.nmosrm_0.outn.n160 bandgapmd_0.otam_1.nmosrm_0.outn.t17 8.265
R27723 bandgapmd_0.otam_1.nmosrm_0.outn.n165 bandgapmd_0.otam_1.nmosrm_0.outn.t19 8.265
R27724 bandgapmd_0.otam_1.nmosrm_0.outn.n165 bandgapmd_0.otam_1.nmosrm_0.outn.t21 8.265
R27725 bandgapmd_0.otam_1.nmosrm_0.outn.n164 bandgapmd_0.otam_1.nmosrm_0.outn.t20 8.265
R27726 bandgapmd_0.otam_1.nmosrm_0.outn.n164 bandgapmd_0.otam_1.nmosrm_0.outn.t22 8.265
R27727 bandgapmd_0.otam_1.nmosrm_0.outn.n180 bandgapmd_0.otam_1.nmosrm_0.outn.t23 8.265
R27728 bandgapmd_0.otam_1.nmosrm_0.outn.n180 bandgapmd_0.otam_1.nmosrm_0.outn.t16 8.265
R27729 bandgapmd_0.otam_1.nmosrm_0.outn.n43 bandgapmd_0.otam_1.nmosrm_0.outn.n42 7.905
R27730 bandgapmd_0.otam_1.nmosrm_0.outn.n136 bandgapmd_0.otam_1.nmosrm_0.outn.n135 7.905
R27731 bandgapmd_0.otam_1.nmosrm_0.outn.n92 bandgapmd_0.otam_1.nmosrm_0.outn.n91 7.529
R27732 bandgapmd_0.otam_1.nmosrm_0.outn.n195 bandgapmd_0.otam_1.nmosrm_0.outn.n194 7.072
R27733 bandgapmd_0.otam_1.nmosrm_0.outn.n229 bandgapmd_0.otam_1.nmosrm_0.outn.n228 7.072
R27734 bandgapmd_0.otam_1.nmosrm_0.outn.n215 bandgapmd_0.otam_1.nmosrm_0.outn.t30 6.923
R27735 bandgapmd_0.otam_1.nmosrm_0.outn.n215 bandgapmd_0.otam_1.nmosrm_0.outn.t31 6.923
R27736 bandgapmd_0.otam_1.nmosrm_0.outn.n224 bandgapmd_0.otam_1.nmosrm_0.outn.t29 6.923
R27737 bandgapmd_0.otam_1.nmosrm_0.outn.n224 bandgapmd_0.otam_1.nmosrm_0.outn.t27 6.923
R27738 bandgapmd_0.otam_1.nmosrm_0.outn.n234 bandgapmd_0.otam_1.nmosrm_0.outn.t26 6.923
R27739 bandgapmd_0.otam_1.nmosrm_0.outn.n234 bandgapmd_0.otam_1.nmosrm_0.outn.t33 6.923
R27740 bandgapmd_0.otam_1.nmosrm_0.outn.n190 bandgapmd_0.otam_1.nmosrm_0.outn.t28 6.923
R27741 bandgapmd_0.otam_1.nmosrm_0.outn.n190 bandgapmd_0.otam_1.nmosrm_0.outn.t25 6.923
R27742 bandgapmd_0.otam_1.nmosrm_0.outn.n204 bandgapmd_0.otam_1.nmosrm_0.outn.t24 6.923
R27743 bandgapmd_0.otam_1.nmosrm_0.outn.n204 bandgapmd_0.otam_1.nmosrm_0.outn.t32 6.923
R27744 bandgapmd_0.otam_1.nmosrm_0.outn.n205 bandgapmd_0.otam_1.nmosrm_0.outn.n203 6.865
R27745 bandgapmd_0.otam_1.nmosrm_0.outn.n216 bandgapmd_0.otam_1.nmosrm_0.outn.n214 6.843
R27746 bandgapmd_0.otam_1.nmosrm_0.outn.n166 bandgapmd_0.otam_1.nmosrm_0.outn.n165 6.641
R27747 bandgapmd_0.otam_1.nmosrm_0.outn.n181 bandgapmd_0.otam_1.nmosrm_0.outn.n180 5.852
R27748 bandgapmd_0.otam_1.nmosrm_0.outn.n161 bandgapmd_0.otam_1.nmosrm_0.outn.n160 5.845
R27749 bandgapmd_0.otam_1.nmosrm_0.outn.n150 bandgapmd_0.otam_1.nmosrm_0.outn.n149 5.27
R27750 bandgapmd_0.otam_1.nmosrm_0.outn.n151 bandgapmd_0.otam_1.nmosrm_0.outn.n150 4.894
R27751 bandgapmd_0.otam_1.nmosrm_0.outn.n16 bandgapmd_0.otam_1.nmosrm_0.outn.n60 4.669
R27752 bandgapmd_0.otam_1.nmosrm_0.outn.n3 bandgapmd_0.otam_1.nmosrm_0.outn.n45 4.65
R27753 bandgapmd_0.otam_1.nmosrm_0.outn.n4 bandgapmd_0.otam_1.nmosrm_0.outn.n138 4.65
R27754 bandgapmd_0.otam_1.nmosrm_0.outn.n2 bandgapmd_0.otam_1.nmosrm_0.outn.n169 4.521
R27755 bandgapmd_0.otam_1.nmosrm_0.outn.n50 bandgapmd_0.otam_1.nmosrm_0.outn.n49 4.5
R27756 bandgapmd_0.otam_1.nmosrm_0.outn.n3 bandgapmd_0.otam_1.nmosrm_0.outn.n44 4.5
R27757 bandgapmd_0.otam_1.nmosrm_0.outn.n9 bandgapmd_0.otam_1.nmosrm_0.outn.n43 4.5
R27758 bandgapmd_0.otam_1.nmosrm_0.outn.n40 bandgapmd_0.otam_1.nmosrm_0.outn.n47 4.5
R27759 bandgapmd_0.otam_1.nmosrm_0.outn.n37 bandgapmd_0.otam_1.nmosrm_0.outn.n36 4.5
R27760 bandgapmd_0.otam_1.nmosrm_0.outn.n30 bandgapmd_0.otam_1.nmosrm_0.outn.n28 4.5
R27761 bandgapmd_0.otam_1.nmosrm_0.outn.n25 bandgapmd_0.otam_1.nmosrm_0.outn.n33 4.5
R27762 bandgapmd_0.otam_1.nmosrm_0.outn.n22 bandgapmd_0.otam_1.nmosrm_0.outn.n56 4.5
R27763 bandgapmd_0.otam_1.nmosrm_0.outn.n79 bandgapmd_0.otam_1.nmosrm_0.outn.n78 4.5
R27764 bandgapmd_0.otam_1.nmosrm_0.outn.n72 bandgapmd_0.otam_1.nmosrm_0.outn.n70 4.5
R27765 bandgapmd_0.otam_1.nmosrm_0.outn.n67 bandgapmd_0.otam_1.nmosrm_0.outn.n75 4.5
R27766 bandgapmd_0.otam_1.nmosrm_0.outn.n143 bandgapmd_0.otam_1.nmosrm_0.outn.n142 4.5
R27767 bandgapmd_0.otam_1.nmosrm_0.outn.n4 bandgapmd_0.otam_1.nmosrm_0.outn.n137 4.5
R27768 bandgapmd_0.otam_1.nmosrm_0.outn.n10 bandgapmd_0.otam_1.nmosrm_0.outn.n136 4.5
R27769 bandgapmd_0.otam_1.nmosrm_0.outn.n133 bandgapmd_0.otam_1.nmosrm_0.outn.n140 4.5
R27770 bandgapmd_0.otam_1.nmosrm_0.outn.n128 bandgapmd_0.otam_1.nmosrm_0.outn.n127 4.5
R27771 bandgapmd_0.otam_1.nmosrm_0.outn.n121 bandgapmd_0.otam_1.nmosrm_0.outn.n119 4.5
R27772 bandgapmd_0.otam_1.nmosrm_0.outn.n116 bandgapmd_0.otam_1.nmosrm_0.outn.n124 4.5
R27773 bandgapmd_0.otam_1.nmosrm_0.outn.n167 bandgapmd_0.otam_1.nmosrm_0.outn.n2 4.5
R27774 bandgapmd_0.otam_1.nmosrm_0.outn.n177 bandgapmd_0.otam_1.nmosrm_0.outn.n176 4.5
R27775 bandgapmd_0.otam_1.nmosrm_0.outn.n99 bandgapmd_0.otam_1.nmosrm_0.outn.n98 4.141
R27776 bandgapmd_0.otam_1.nmosrm_0.outn.n5 bandgapmd_0.otam_1.nmosrm_0.outn.n164 4.06
R27777 bandgapmd_0.otam_1.nmosrm_0.outn.n94 bandgapmd_0.otam_1.nmosrm_0.outn.n93 3.764
R27778 bandgapmd_0.otam_1.nmosrm_0.outn.n175 bandgapmd_0.otam_1.nmosrm_0.outn.n174 3.688
R27779 bandgapmd_0.otam_1.nmosrm_0.outn.n47 bandgapmd_0.otam_1.nmosrm_0.outn.n46 3.388
R27780 bandgapmd_0.otam_1.nmosrm_0.outn.n78 bandgapmd_0.otam_1.nmosrm_0.outn.n76 3.388
R27781 bandgapmd_0.otam_1.nmosrm_0.outn.n140 bandgapmd_0.otam_1.nmosrm_0.outn.n139 3.388
R27782 bandgapmd_0.otam_1.nmosrm_0.outn.n13 bandgapmd_0.otam_1.nmosrm_0.outn.n94 3.111
R27783 bandgapmd_0.otam_1.nmosrm_0.outn.n16 bandgapmd_0.otam_1.nmosrm_0.outn.n58 3.033
R27784 bandgapmd_0.otam_1.nmosrm_0.outn.n100 bandgapmd_0.otam_1.nmosrm_0.outn.n99 3.033
R27785 bandgapmd_0.otam_1.nmosrm_0.outn.n13 bandgapmd_0.otam_1.nmosrm_0.outn.n92 3.033
R27786 bandgapmd_0.otam_1.nmosrm_0.outn.n89 bandgapmd_0.otam_1.nmosrm_0.outn.n97 3.033
R27787 bandgapmd_0.otam_1.nmosrm_0.outn.n20 bandgapmd_0.otam_1.nmosrm_0.outn.n107 3.033
R27788 bandgapmd_0.otam_1.nmosrm_0.outn.n23 bandgapmd_0.otam_1.nmosrm_0.outn.n112 3.033
R27789 bandgapmd_0.otam_1.nmosrm_0.outn.n0 bandgapmd_0.otam_1.nmosrm_0.outn.n151 3.029
R27790 bandgapmd_0.otam_1.nmosrm_0.outn.n43 bandgapmd_0.otam_1.nmosrm_0.outn.n41 3.011
R27791 bandgapmd_0.otam_1.nmosrm_0.outn.n36 bandgapmd_0.otam_1.nmosrm_0.outn.n35 3.011
R27792 bandgapmd_0.otam_1.nmosrm_0.outn.n70 bandgapmd_0.otam_1.nmosrm_0.outn.n69 3.011
R27793 bandgapmd_0.otam_1.nmosrm_0.outn.n97 bandgapmd_0.otam_1.nmosrm_0.outn.n96 3.011
R27794 bandgapmd_0.otam_1.nmosrm_0.outn.n136 bandgapmd_0.otam_1.nmosrm_0.outn.n134 3.011
R27795 bandgapmd_0.otam_1.nmosrm_0.outn.n127 bandgapmd_0.otam_1.nmosrm_0.outn.n126 3.011
R27796 bandgapmd_0.otam_1.nmosrm_0.outn.n131 bandgapmd_0.otam_1.nmosrm_0.outn.n130 2.748
R27797 bandgapmd_0.otam_1.nmosrm_0.outn.n28 bandgapmd_0.otam_1.nmosrm_0.outn.n27 2.635
R27798 bandgapmd_0.otam_1.nmosrm_0.outn.n92 bandgapmd_0.otam_1.nmosrm_0.outn.n90 2.635
R27799 bandgapmd_0.otam_1.nmosrm_0.outn.n119 bandgapmd_0.otam_1.nmosrm_0.outn.n118 2.635
R27800 bandgapmd_0.otam_1.pdiffm_0.outn bandgapmd_0.otam_1.nmosrm_0.outn.n237 2.345
R27801 bandgapmd_0.otam_1.nmosrm_0.outn.n199 bandgapmd_0.otam_1.nmosrm_0.outn.n198 2.328
R27802 bandgapmd_0.otam_1.nmosrm_0.outn.n211 bandgapmd_0.otam_1.nmosrm_0.outn.n189 2.31
R27803 bandgapmd_0.otam_1.nmosrm_0.outn.n223 bandgapmd_0.otam_1.nmosrm_0.outn.n222 2.304
R27804 bandgapmd_0.otam_1.nmosrm_0.outn.n191 bandgapmd_0.otam_1.nmosrm_0.outn.n190 2.302
R27805 bandgapmd_0.otam_1.nmosrm_0.outn.n205 bandgapmd_0.otam_1.nmosrm_0.outn.n204 2.288
R27806 bandgapmd_0.otam_1.nmosrm_0.outn.n216 bandgapmd_0.otam_1.nmosrm_0.outn.n215 2.288
R27807 bandgapmd_0.otam_1.nmosrm_0.outn.n171 bandgapmd_0.otam_1.nmosrm_0.outn.n170 2.286
R27808 bandgapmd_0.otam_1.nmosrm_0.outn.n88 bandgapmd_0.otam_1.nmosrm_0.outn.n39 3.062
R27809 bandgapmd_0.otam_1.nmosrm_0.outn.n85 bandgapmd_0.otam_1.nmosrm_0.outn.n51 3.059
R27810 bandgapmd_0.otam_1.nmosrm_0.outn.n168 bandgapmd_0.otam_1.nmosrm_0.outn.n166 2.272
R27811 bandgapmd_0.otam_1.nmosrm_0.outn.n65 bandgapmd_0.otam_1.nmosrm_0.outn.n62 3.062
R27812 bandgapmd_0.otam_1.nmosrm_0.outn.n221 bandgapmd_0.otam_1.nmosrm_0.outn.n220 2.259
R27813 bandgapmd_0.otam_1.nmosrm_0.outn.n210 bandgapmd_0.otam_1.nmosrm_0.outn.n209 2.259
R27814 bandgapmd_0.otam_1.nmosrm_0.outn.n233 bandgapmd_0.otam_1.nmosrm_0.outn.n232 2.258
R27815 bandgapmd_0.otam_1.nmosrm_0.outn.n75 bandgapmd_0.otam_1.nmosrm_0.outn.n74 2.258
R27816 bandgapmd_0.otam_1.nmosrm_0.outn.n185 bandgapmd_0.otam_1.nmosrm_0.outn.n184 2.254
R27817 bandgapmd_0.otam_1.nmosrm_0.outn.n145 bandgapmd_0.otam_1.nmosrm_0.outn.n144 3.035
R27818 bandgapmd_0.otam_1.nmosrm_0.outn.n188 bandgapmd_0.otam_1.nmosrm_0.outn.n187 2.389
R27819 bandgapmd_0.otam_1.nmosrm_0.outn.n8 bandgapmd_0.otam_1.nmosrm_0.outn.n178 2.25
R27820 bandgapmd_0.otam_1.nmosrm_0.outn.n33 bandgapmd_0.otam_1.nmosrm_0.outn.n32 1.882
R27821 bandgapmd_0.otam_1.nmosrm_0.outn.n124 bandgapmd_0.otam_1.nmosrm_0.outn.n123 1.882
R27822 bandgapmd_0.otam_1.nmosrm_0.outn.n187 bandgapmd_0.otam_1.nmosrm_0.outn.n186 1.782
R27823 bandgapmd_0.otam_1.nmosrm_0.outn.n63 bandgapmd_0.otam_1.pdiffaloadm_0.outn 1.649
R27824 bandgapmd_0.otam_1.nmosrm_0.outn.n225 bandgapmd_0.otam_1.nmosrm_0.outn.n224 1.577
R27825 bandgapmd_0.otam_1.nmosrm_0.outn.n82 bandgapmd_0.otam_1.nmosrm_0.outn.n81 1.513
R27826 bandgapmd_0.otam_1.nmosrm_0.outn.n146 bandgapmd_0.otam_1.nmosrm_0.outn.n114 1.505
R27827 bandgapmd_0.otam_1.nmosrm_0.outn.n147 bandgapmd_0.otam_1.nmosrm_0.outn.n101 1.491
R27828 bandgapmd_0.otam_1.nmosrm_0.outn.n186 bandgapmd_0.otam_1.nmosrm_0.outn.n163 1.597
R27829 bandgapmd_0.otam_1.nmosrm_0.outn.n12 bandgapmd_0.otam_1.nmosrm_0.outn.n234 1.452
R27830 bandgapmd_0.otam_1.nmosrm_0.outn.n171 bandgapmd_0.otam_1.nmosrm_0.outn 1.44
R27831 bandgapmd_0.otam_1.nmosrm_0.outn.n147 bandgapmd_0.otam_1.nmosrm_0.outn.n146 1.328
R27832 bandgapmd_0.otam_1.nmosrm_0.outn.n82 bandgapmd_0.otam_1.nmosrm_0.outn.n65 1.294
R27833 bandgapmd_0.otam_1.nmosrm_0.outn.n146 bandgapmd_0.otam_1.nmosrm_0.outn.n145 1.275
R27834 bandgapmd_0.otam_1.nmosrm_0.outn.n83 bandgapmd_0.otam_1.nmosrm_0.outn.n82 1.246
R27835 bandgapmd_0.otam_1.nmosrm_0.outn.n86 bandgapmd_0.otam_1.nmosrm_0.outn.n85 1.169
R27836 bandgapmd_0.otam_1.nmosrm_0.outn.n6 bandgapmd_0.otam_1.nmosrm_0.outn.n5 0.748
R27837 bandgapmd_0.otam_1.nmosrm_0.outn.n101 bandgapmd_0.otam_1.nmosrm_0.outn.n89 1.127
R27838 bandgapmd_0.otam_1.nmosrm_0.outn.n114 bandgapmd_0.otam_1.nmosrm_0.outn.n23 1.124
R27839 bandgapmd_0.otam_1.nmosrm_0.outn.n197 bandgapmd_0.otam_1.nmosrm_0.outn.n7 1.033
R27840 bandgapmd_0.otam_1.nmosrm_0.outn.n17 bandgapmd_0.otam_1.nmosrm_0.outn.n225 1.005
R27841 bandgapmd_0.otam_1.nmosrm_0.outn.n163 bandgapmd_0.otam_1.nmosrm_0.outn.n162 0.969
R27842 bandgapmd_0.otam_1.nmosrm_0.outn.n211 bandgapmd_0.otam_1.nmosrm_0.outn.n210 0.966
R27843 bandgapmd_0.otam_1.nmosrm_0.outn.n223 bandgapmd_0.otam_1.nmosrm_0.outn.n221 0.957
R27844 bandgapmd_0.otam_1.nmosrm_0.outn.n199 bandgapmd_0.otam_1.nmosrm_0.outn.n197 0.955
R27845 bandgapmd_0.otam_1.nmosrm_0.outn.n38 bandgapmd_0.otam_1.nmosrm_0.outn.n37 0.944
R27846 bandgapmd_0.otam_1.nmosrm_0.outn.n129 bandgapmd_0.otam_1.nmosrm_0.outn.n128 0.941
R27847 bandgapmd_0.otam_1.nmosrm_0.outn.n80 bandgapmd_0.otam_1.nmosrm_0.outn.n79 0.941
R27848 bandgapmd_0.otam_1.pdiffm_0.outn bandgapmd_0.otam_1.nmosrm_0.outn.n233 0.925
R27849 bandgapmd_0.otam_1.nmosrm_0.outn.n130 bandgapmd_0.otam_1.nmosrm_0.outn.n116 0.9
R27850 bandgapmd_0.otam_1.nmosrm_0.outn.n39 bandgapmd_0.otam_1.nmosrm_0.outn.n25 0.899
R27851 bandgapmd_0.otam_1.nmosrm_0.outn.n51 bandgapmd_0.otam_1.nmosrm_0.outn.n40 0.898
R27852 bandgapmd_0.otam_1.nmosrm_0.outn.n81 bandgapmd_0.otam_1.nmosrm_0.outn.n67 0.898
R27853 bandgapmd_0.otam_1.nmosrm_0.outn.n62 bandgapmd_0.otam_1.nmosrm_0.outn.n22 0.898
R27854 bandgapmd_0.otam_1.nmosrm_0.outn.n144 bandgapmd_0.otam_1.nmosrm_0.outn.n133 0.896
R27855 bandgapmd_0.otam_1.nmosrm_0.outn.n107 bandgapmd_0.otam_1.nmosrm_0.outn.n106 0.752
R27856 bandgapmd_0.otam_1.nmosrm_0.outn bandgapmd_0.otam_1.nmosrm_0.outn.n6 0.62
R27857 bandgapmd_0.otam_1.nmosrm_0.outn.n148 bandgapmd_0.otam_1.nmosrm_0.outn.n147 0.518
R27858 bandgapmd_0.otam_1.nmosrm_0.outn.n186 bandgapmd_0.otam_1.nmosrm_0.outn.n185 0.46
R27859 bandgapmd_0.otam_1.nmosrm_0.outn.n169 bandgapmd_0.otam_1.nmosrm_0.outn.n168 0.45
R27860 bandgapmd_0.otam_1.nmosrm_0.outn.n56 bandgapmd_0.otam_1.nmosrm_0.outn.n55 0.376
R27861 bandgapmd_0.otam_1.nmosrm_0.outn.n112 bandgapmd_0.otam_1.nmosrm_0.outn.n111 0.376
R27862 bandgapmd_0.otam_1.nmosrm_0.outn.n18 bandgapmd_0.otam_1.nmosrm_0.outn.n229 0.355
R27863 bandgapmd_0.otam_1.nmosrm_0.outn.n19 bandgapmd_0.otam_1.nmosrm_0.outn.n212 0.348
R27864 bandgapmd_0.otam_1.nmosrm_0.outn.n1 bandgapmd_0.otam_1.nmosrm_0.outn.n201 0.348
R27865 bandgapmd_0.otam_1.nmosrm_0.outn.n7 bandgapmd_0.otam_1.nmosrm_0.outn.n195 0.345
R27866 bandgapmd_0.otam_1.nmosrm_0.outn.n148 bandgapmd_0.otam_1.nmosrm_0.outn.n88 0.34
R27867 bandgapmd_0.otam_1.nmosrm_0.outn.n182 bandgapmd_0.otam_1.nmosrm_0.outn.n181 0.313
R27868 bandgapmd_0.otam_1.nmosrm_0.outn.n0 bandgapmd_0.otam_1.nmosrm_0.outn.n161 0.311
R27869 bandgapmd_0.otam_1.nmosrm_0.outn.n206 bandgapmd_0.otam_1.nmosrm_0.outn.n205 0.29
R27870 bandgapmd_0.otam_1.nmosrm_0.outn.n217 bandgapmd_0.otam_1.nmosrm_0.outn.n216 0.29
R27871 bandgapmd_0.otam_1.nmosrm_0.outn.n192 bandgapmd_0.otam_1.nmosrm_0.outn.n191 0.287
R27872 bandgapmd_0.otam_1.nmosrm_0.outn.n220 bandgapmd_0.otam_1.nmosrm_0.outn.n19 0.189
R27873 bandgapmd_0.otam_1.nmosrm_0.outn.n187 bandgapmd_0.otam_1.nmosrm_0.outn.n148 0.168
R27874 bandgapmd_0.otam_1.nmosrm_0.outn.n220 bandgapmd_0.otam_1.nmosrm_0.outn.n219 0.162
R27875 bandgapmd_0.otam_1.nmosrm_0.outn.n209 bandgapmd_0.otam_1.nmosrm_0.outn.n1 0.159
R27876 bandgapmd_0.otam_1.nmosrm_0.outn.n7 bandgapmd_0.otam_1.nmosrm_0.outn.n196 0.148
R27877 bandgapmd_0.otam_1.nmosrm_0.outn.n232 bandgapmd_0.otam_1.nmosrm_0.outn.n231 0.145
R27878 bandgapmd_0.otam_1.nmosrm_0.outn.n209 bandgapmd_0.otam_1.nmosrm_0.outn.n208 0.143
R27879 bandgapmd_0.otam_1.nmosrm_0.outn.n159 bandgapmd_0.otam_1.nmosrm_0.outn.n15 0.125
R27880 bandgapmd_0.otam_1.nmosrm_0.outn.n19 bandgapmd_0.otam_1.nmosrm_0.outn.n218 0.119
R27881 bandgapmd_0.otam_1.nmosrm_0.outn.n153 bandgapmd_0.otam_1.nmosrm_0.outn.n152 0.116
R27882 bandgapmd_0.otam_1.nmosrm_0.outn.n18 bandgapmd_0.otam_1.nmosrm_0.outn.n227 0.107
R27883 bandgapmd_0.otam_1.nmosrm_0.outn.n81 bandgapmd_0.otam_1.nmosrm_0.outn.n80 0.095
R27884 bandgapmd_0.otam_1.nmosrm_0.outn.n39 bandgapmd_0.otam_1.nmosrm_0.outn.n38 0.095
R27885 bandgapmd_0.otam_1.nmosrm_0.outn.n114 bandgapmd_0.otam_1.nmosrm_0.outn.n113 0.095
R27886 bandgapmd_0.otam_1.nmosrm_0.outn.n130 bandgapmd_0.otam_1.nmosrm_0.outn.n129 0.095
R27887 bandgapmd_0.otam_1.nmosrm_0.outn.n177 bandgapmd_0.otam_1.nmosrm_0.outn.n173 0.092
R27888 bandgapmd_0.otam_1.pdiffm_0.outn bandgapmd_0.otam_1.nmosrm_0.outn.n188 0.092
R27889 bandgapmd_0.otam_1.nmosrm_0.outn.n7 bandgapmd_0.otam_1.nmosrm_0.outn.n193 0.091
R27890 bandgapmd_0.otam_1.nmosrm_0.outn.n168 bandgapmd_0.otam_1.nmosrm_0.outn.n167 0.084
R27891 bandgapmd_0.otam_1.nmosrm_0.outn.n88 bandgapmd_0.otam_1.nmosrm_0.outn.n87 0.083
R27892 bandgapmd_0.otam_1.nmosrm_0.outn.n87 bandgapmd_0.otam_1.nmosrm_0.outn.n86 0.083
R27893 bandgapmd_0.otam_1.nmosrm_0.outn.n85 bandgapmd_0.otam_1.nmosrm_0.outn.n84 0.083
R27894 bandgapmd_0.otam_1.nmosrm_0.outn.n84 bandgapmd_0.otam_1.nmosrm_0.outn.n83 0.083
R27895 bandgapmd_0.otam_1.nmosrm_0.outn.n65 bandgapmd_0.otam_1.nmosrm_0.outn.n64 0.083
R27896 bandgapmd_0.otam_1.nmosrm_0.outn.n64 bandgapmd_0.otam_1.nmosrm_0.outn.n63 0.083
R27897 bandgapmd_0.otam_1.nmosrm_0.outn.n132 bandgapmd_0.otam_1.nmosrm_0.outn.n131 0.083
R27898 bandgapmd_0.otam_1.nmosrm_0.outn.n145 bandgapmd_0.otam_1.nmosrm_0.outn.n132 0.083
R27899 bandgapmd_0.otam_1.nmosrm_0.outn.n12 bandgapmd_0.otam_1.nmosrm_0.outn.n236 0.08
R27900 bandgapmd_0.otam_1.nmosrm_0.outn.n11 bandgapmd_0.otam_1.nmosrm_0.outn.n207 0.076
R27901 bandgapmd_0.otam_1.nmosrm_0.outn.n184 bandgapmd_0.otam_1.nmosrm_0.outn.n183 0.075
R27902 bandgapmd_0.otam_1.nmosrm_0.outn.n207 bandgapmd_0.otam_1.nmosrm_0.outn.n206 0.075
R27903 bandgapmd_0.otam_1.nmosrm_0.outn.n18 bandgapmd_0.otam_1.nmosrm_0.outn.n226 0.073
R27904 bandgapmd_0.otam_1.nmosrm_0.outn.n231 bandgapmd_0.otam_1.nmosrm_0.outn.n18 0.07
R27905 bandgapmd_0.otam_1.nmosrm_0.outn.n233 bandgapmd_0.otam_1.nmosrm_0.outn.n223 0.133
R27906 bandgapmd_0.otam_1.nmosrm_0.outn.n221 bandgapmd_0.otam_1.nmosrm_0.outn.n211 0.133
R27907 bandgapmd_0.otam_1.nmosrm_0.outn.n169 bandgapmd_0.otam_1.nmosrm_0.outn.n5 0.067
R27908 bandgapmd_0.otam_1.nmosrm_0.outn.n0 bandgapmd_0.otam_1.nmosrm_0.outn.n153 0.066
R27909 bandgapmd_0.otam_1.nmosrm_0.outn.n8 bandgapmd_0.otam_1.nmosrm_0.outn.n171 0.066
R27910 bandgapmd_0.otam_1.nmosrm_0.outn.n210 bandgapmd_0.otam_1.nmosrm_0.outn.n199 0.133
R27911 bandgapmd_0.otam_1.nmosrm_0.outn.n185 bandgapmd_0.otam_1.nmosrm_0.outn.n179 0.063
R27912 bandgapmd_0.otam_1.nmosrm_0.outn.n0 bandgapmd_0.otam_1.nmosrm_0.outn.n155 0.062
R27913 bandgapmd_0.otam_1.nmosrm_0.outn.n166 bandgapmd_0.otam_1.nmosrm_0.outn.n2 0.059
R27914 bandgapmd_0.otam_1.nmosrm_0.outn.n0 bandgapmd_0.otam_1.nmosrm_0.outn.n159 0.056
R27915 bandgapmd_0.otam_1.nmosrm_0.outn.n11 bandgapmd_0.otam_1.nmosrm_0.outn.n202 0.055
R27916 bandgapmd_0.otam_1.nmosrm_0.outn.n18 bandgapmd_0.otam_1.nmosrm_0.outn.n230 0.054
R27917 bandgapmd_0.otam_1.nmosrm_0.outn.n12 bandgapmd_0.otam_1.nmosrm_0.outn.n235 0.053
R27918 bandgapmd_0.otam_1.nmosrm_0.outn.n24 bandgapmd_0.otam_1.nmosrm_0.outn.n30 0.09
R27919 bandgapmd_0.otam_1.nmosrm_0.outn.n54 bandgapmd_0.otam_1.nmosrm_0.outn.n53 0.044
R27920 bandgapmd_0.otam_1.nmosrm_0.outn.n66 bandgapmd_0.otam_1.nmosrm_0.outn.n72 0.09
R27921 bandgapmd_0.otam_1.nmosrm_0.outn.n115 bandgapmd_0.otam_1.nmosrm_0.outn.n121 0.09
R27922 bandgapmd_0.otam_1.nmosrm_0.outn.n110 bandgapmd_0.otam_1.nmosrm_0.outn.n109 0.043
R27923 bandgapmd_0.otam_1.nmosrm_0.outn.n101 bandgapmd_0.otam_1.nmosrm_0.outn.n100 1.269
R27924 bandgapmd_0.otam_1.nmosrm_0.outn.n144 bandgapmd_0.otam_1.nmosrm_0.outn.n143 1.035
R27925 bandgapmd_0.otam_1.nmosrm_0.outn.n51 bandgapmd_0.otam_1.nmosrm_0.outn.n50 1.035
R27926 bandgapmd_0.otam_1.nmosrm_0.outn.n61 bandgapmd_0.otam_1.nmosrm_0.outn.n16 0.989
R27927 bandgapmd_0.otam_1.nmosrm_0.outn.n10 bandgapmd_0.otam_1.nmosrm_0.outn.n4 0.098
R27928 bandgapmd_0.otam_1.nmosrm_0.outn.n9 bandgapmd_0.otam_1.nmosrm_0.outn.n3 0.098
R27929 bandgapmd_0.otam_1.nmosrm_0.outn.n7 bandgapmd_0.otam_1.nmosrm_0.outn.n192 0.078
R27930 bandgapmd_0.otam_1.nmosrm_0.outn.n1 bandgapmd_0.otam_1.nmosrm_0.outn.n200 0.075
R27931 bandgapmd_0.otam_1.nmosrm_0.outn.n167 bandgapmd_0.otam_1.nmosrm_0.outn.n5 0.056
R27932 bandgapmd_0.otam_1.nmosrm_0.outn.n2 bandgapmd_0.otam_1.nmosrm_0.outn.n6 0.054
R27933 bandgapmd_0.otam_1.nmosrm_0.outn.n162 bandgapmd_0.otam_1.nmosrm_0.outn.n0 0.047
R27934 bandgapmd_0.otam_1.nmosrm_0.outn.n89 bandgapmd_0.otam_1.nmosrm_0.outn.n13 0.04
R27935 bandgapmd_0.otam_1.nmosrm_0.outn.n133 bandgapmd_0.otam_1.nmosrm_0.outn.n10 0.04
R27936 bandgapmd_0.otam_1.nmosrm_0.outn.n40 bandgapmd_0.otam_1.nmosrm_0.outn.n9 0.04
R27937 bandgapmd_0.otam_1.nmosrm_0.outn.n208 bandgapmd_0.otam_1.nmosrm_0.outn.n11 0.036
R27938 bandgapmd_0.otam_1.nmosrm_0.outn.n178 bandgapmd_0.otam_1.nmosrm_0.outn.n177 0.034
R27939 bandgapmd_0.otam_1.nmosrm_0.outn.n22 bandgapmd_0.otam_1.nmosrm_0.outn.n54 0.034
R27940 bandgapmd_0.otam_1.nmosrm_0.outn.n237 bandgapmd_0.otam_1.nmosrm_0.outn.n12 0.033
R27941 bandgapmd_0.otam_1.nmosrm_0.outn.n19 bandgapmd_0.otam_1.nmosrm_0.outn.n217 0.032
R27942 bandgapmd_0.otam_1.nmosrm_0.outn.n179 bandgapmd_0.otam_1.nmosrm_0.outn.n8 0.032
R27943 bandgapmd_0.otam_1.nmosrm_0.outn.n62 bandgapmd_0.otam_1.nmosrm_0.outn.n61 0.032
R27944 bandgapmd_0.otam_1.nmosrm_0.outn.n183 bandgapmd_0.otam_1.nmosrm_0.outn.n182 0.031
R27945 bandgapmd_0.otam_1.nmosrm_0.outn.n23 bandgapmd_0.otam_1.nmosrm_0.outn.n110 0.03
R27946 bandgapmd_0.otam_1.nmosrm_0.outn.n15 bandgapmd_0.otam_1.nmosrm_0.outn.n14 0.03
R27947 bandgapmd_0.otam_1.nmosrm_0.outn.n25 bandgapmd_0.otam_1.nmosrm_0.outn.n24 0.029
R27948 bandgapmd_0.otam_1.nmosrm_0.outn.n67 bandgapmd_0.otam_1.nmosrm_0.outn.n66 0.029
R27949 bandgapmd_0.otam_1.nmosrm_0.outn.n116 bandgapmd_0.otam_1.nmosrm_0.outn.n115 0.029
R27950 bandgapmd_0.otam_1.nmosrm_0.outn.n178 bandgapmd_0.otam_1.nmosrm_0.outn.n172 0.029
R27951 bandgapmd_0.otam_1.nmosrm_0.outn.n20 bandgapmd_0.otam_1.nmosrm_0.outn.n21 0.029
R27952 bandgapmd_0.otam_1.nmosrm_0.outn.n19 bandgapmd_0.otam_1.nmosrm_0.outn.n213 0.029
R27953 bandgapmd_0.otam_1.nmosrm_0.outn.n53 bandgapmd_0.otam_1.nmosrm_0.outn.n52 0.028
R27954 bandgapmd_0.otam_1.nmosrm_0.outn.n177 bandgapmd_0.otam_1.nmosrm_0.outn.n175 0.027
R27955 bandgapmd_0.otam_1.nmosrm_0.outn.n30 bandgapmd_0.otam_1.nmosrm_0.outn.n29 0.026
R27956 bandgapmd_0.otam_1.nmosrm_0.outn.n121 bandgapmd_0.otam_1.nmosrm_0.outn.n120 0.026
R27957 bandgapmd_0.otam_1.nmosrm_0.outn.n72 bandgapmd_0.otam_1.nmosrm_0.outn.n71 0.024
R27958 bandgapmd_0.otam_1.nmosrm_0.outn.n109 bandgapmd_0.otam_1.nmosrm_0.outn.n108 0.024
R27959 bandgapmd_0.otam_1.nmosrm_0.outn.n18 bandgapmd_0.otam_1.nmosrm_0.outn.n17 0.024
R27960 bandgapmd_0.otam_1.nmosrm_0.outn.n108 bandgapmd_0.otam_1.nmosrm_0.outn.n20 0.023
R27961 vdd.n8145 vdd.n8134 47025
R27962 vdd.n13082 vdd.n9287 19665.9
R27963 vdd.n12568 vdd.n10478 13311.6
R27964 vdd.n11601 vdd.n10517 13306.7
R27965 vdd.n13084 vdd.n13083 4529.64
R27966 vdd.n31150 vdd.t232 2454.41
R27967 vdd.n30323 vdd.t216 2454.31
R27968 vdd.n38138 vdd.t208 2454.26
R27969 vdd.n1731 vdd.t229 2454.26
R27970 vdd.n11739 vdd.n11726 585
R27971 vdd.n11741 vdd.n11740 585
R27972 vdd.n11823 vdd.n11821 585
R27973 vdd.n11825 vdd.n11824 585
R27974 vdd.n21914 vdd.n21912 585
R27975 vdd.n21916 vdd.n21915 585
R27976 vdd.n14501 vdd.n8198 416.689
R27977 vdd.n13116 vdd.n9273 416.689
R27978 vdd.n14657 vdd.n8144 408.826
R27979 vdd.n14943 vdd.n7988 408.826
R27980 vdd.n14528 vdd.n8211 395.068
R27981 vdd.n13108 vdd.n9272 395.068
R27982 vdd.n14616 vdd.n14615 389.171
R27983 vdd.n11630 vdd.n11629 389.171
R27984 vdd.n14642 vdd.n8168 387.206
R27985 vdd.n11656 vdd.n11575 387.206
R27986 vdd.n14600 vdd.n8147 385.24
R27987 vdd.n14971 vdd.n7985 385.24
R27988 vdd.n22359 vdd.n22356 299.702
R27989 vdd.n22225 vdd.n22222 299.702
R27990 vdd.n22251 vdd.n22248 299.702
R27991 vdd.n22265 vdd.n22262 299.702
R27992 vdd.n22088 vdd.n22085 299.702
R27993 vdd.n22101 vdd.n22098 299.702
R27994 vdd.n22127 vdd.n22124 299.702
R27995 vdd.n22150 vdd.n22147 299.702
R27996 vdd.n11911 vdd.n11910 299.681
R27997 vdd.n11732 vdd.n11730 292.5
R27998 vdd.n11715 vdd.n11714 292.5
R27999 vdd.n11715 vdd.n11693 292.5
R28000 vdd.n11832 vdd.n11813 292.5
R28001 vdd.n11854 vdd.n11837 292.5
R28002 vdd.n11840 vdd.n11837 292.5
R28003 vdd.n21923 vdd.n21904 292.5
R28004 vdd.n21945 vdd.n21928 292.5
R28005 vdd.n21931 vdd.n21928 292.5
R28006 vdd.n11733 vdd.t188 226.827
R28007 vdd.n21808 vdd.t179 226.827
R28008 vdd.n11834 vdd.n11833 226.827
R28009 vdd.n21925 vdd.n21924 226.827
R28010 vdd.n10240 vdd.n10228 189.131
R28011 vdd.n10237 vdd.n10228 188.642
R28012 vdd.n10488 vdd.n10482 188.09
R28013 vdd.n10482 vdd.n10121 187.18
R28014 vdd.n10390 vdd.n10389 185.005
R28015 vdd.n8133 vdd.n8131 185
R28016 vdd.n14673 vdd.n8133 185
R28017 vdd.n14694 vdd.n14693 185
R28018 vdd.n14695 vdd.n14694 185
R28019 vdd.n14683 vdd.n14682 185
R28020 vdd.n14684 vdd.n14683 185
R28021 vdd.n8112 vdd.n8111 185
R28022 vdd.n14713 vdd.n8112 185
R28023 vdd.n14740 vdd.n14739 185
R28024 vdd.n14741 vdd.n14740 185
R28025 vdd.n14723 vdd.n14722 185
R28026 vdd.n14730 vdd.n14723 185
R28027 vdd.n14750 vdd.n14749 185
R28028 vdd.n14749 vdd.n14748 185
R28029 vdd.n8093 vdd.n8092 185
R28030 vdd.n14759 vdd.n8093 185
R28031 vdd.n14772 vdd.n14771 185
R28032 vdd.n14773 vdd.n14772 185
R28033 vdd.n8070 vdd.n8069 185
R28034 vdd.n8072 vdd.n8070 185
R28035 vdd.n14786 vdd.n14785 185
R28036 vdd.n14787 vdd.n14786 185
R28037 vdd.n8079 vdd.n8078 185
R28038 vdd.n14780 vdd.n8079 185
R28039 vdd.n8063 vdd.n8061 185
R28040 vdd.n14801 vdd.n8063 185
R28041 vdd.n14827 vdd.n14826 185
R28042 vdd.n14828 vdd.n14827 185
R28043 vdd.n14810 vdd.n14809 185
R28044 vdd.n14817 vdd.n14810 185
R28045 vdd.n14836 vdd.n14835 185
R28046 vdd.n14835 vdd.n14834 185
R28047 vdd.n8043 vdd.n8041 185
R28048 vdd.n14845 vdd.n8043 185
R28049 vdd.n14868 vdd.n14867 185
R28050 vdd.n14869 vdd.n14868 185
R28051 vdd.n14857 vdd.n14853 185
R28052 vdd.n14858 vdd.n14857 185
R28053 vdd.n14905 vdd.n14904 185
R28054 vdd.n14906 vdd.n14905 185
R28055 vdd.n14885 vdd.n14884 185
R28056 vdd.n14895 vdd.n14885 185
R28057 vdd.n8015 vdd.n8014 185
R28058 vdd.n14913 vdd.n8015 185
R28059 vdd.n14925 vdd.n14924 185
R28060 vdd.n14926 vdd.n14925 185
R28061 vdd.n8008 vdd.n8006 185
R28062 vdd.n14931 vdd.n8008 185
R28063 vdd.n14929 vdd.n14928 185
R28064 vdd.n14930 vdd.n14929 185
R28065 vdd.n14916 vdd.n14915 185
R28066 vdd.n14915 vdd.n14914 185
R28067 vdd.n14903 vdd.n8023 185
R28068 vdd.n8023 vdd.n8021 185
R28069 vdd.n8038 vdd.n8036 185
R28070 vdd.n8036 vdd.n8034 185
R28071 vdd.n8049 vdd.n8048 185
R28072 vdd.n8050 vdd.n8049 185
R28073 vdd.n8058 vdd.n8056 185
R28074 vdd.n8056 vdd.n8054 185
R28075 vdd.n14783 vdd.n14782 185
R28076 vdd.n14782 vdd.n14781 185
R28077 vdd.n14784 vdd.n8075 185
R28078 vdd.n8075 vdd.n8073 185
R28079 vdd.n14770 vdd.n8085 185
R28080 vdd.n8085 vdd.n8083 185
R28081 vdd.n14751 vdd.n8095 185
R28082 vdd.n8095 vdd.n8094 185
R28083 vdd.n14738 vdd.n8107 185
R28084 vdd.n8107 vdd.n8105 185
R28085 vdd.n14687 vdd.n14686 185
R28086 vdd.n14686 vdd.n14685 185
R28087 vdd.n14671 vdd.n14670 185
R28088 vdd.n14672 vdd.n14671 185
R28089 vdd.n8128 vdd.n8126 185
R28090 vdd.n8126 vdd.n8124 185
R28091 vdd.n14716 vdd.n14715 185
R28092 vdd.n14715 vdd.n14714 185
R28093 vdd.n14728 vdd.n14727 185
R28094 vdd.n14729 vdd.n14728 185
R28095 vdd.n14762 vdd.n14761 185
R28096 vdd.n14761 vdd.n14760 185
R28097 vdd.n14791 vdd.n14790 185
R28098 vdd.n14790 vdd.n14789 185
R28099 vdd.n14799 vdd.n14798 185
R28100 vdd.n14800 vdd.n14799 185
R28101 vdd.n14820 vdd.n14819 185
R28102 vdd.n14819 vdd.n14818 185
R28103 vdd.n14843 vdd.n14842 185
R28104 vdd.n14844 vdd.n14843 185
R28105 vdd.n14861 vdd.n14860 185
R28106 vdd.n14860 vdd.n14859 185
R28107 vdd.n14893 vdd.n14892 185
R28108 vdd.n14894 vdd.n14893 185
R28109 vdd.n14923 vdd.n8007 185
R28110 vdd.n14927 vdd.n8007 185
R28111 vdd.n7985 vdd.n7983 185
R28112 vdd.n7987 vdd.n7985 185
R28113 vdd.n14941 vdd.n14940 185
R28114 vdd.n14942 vdd.n14941 185
R28115 vdd.n14655 vdd.n14654 185
R28116 vdd.n14656 vdd.n14655 185
R28117 vdd.n8154 vdd.n8153 185
R28118 vdd.n14645 vdd.n8154 185
R28119 vdd.n14664 vdd.n14663 185
R28120 vdd.n14663 vdd.n14662 185
R28121 vdd.n14648 vdd.n14647 185
R28122 vdd.n14647 vdd.n14646 185
R28123 vdd.n8149 vdd.n8147 185
R28124 vdd.n8173 vdd.n8147 185
R28125 vdd.n8139 vdd.n8138 185
R28126 vdd.n8140 vdd.n8139 185
R28127 vdd.n14359 vdd.n14358 185
R28128 vdd.n14360 vdd.n14359 185
R28129 vdd.n14329 vdd.n14328 185
R28130 vdd.n14328 vdd.n14327 185
R28131 vdd.n14282 vdd.n14281 185
R28132 vdd.n14283 vdd.n14282 185
R28133 vdd.n8406 vdd.n8404 185
R28134 vdd.n8408 vdd.n8406 185
R28135 vdd.n14072 vdd.n14071 185
R28136 vdd.n14071 vdd.n8541 185
R28137 vdd.n14054 vdd.n14053 185
R28138 vdd.n14053 vdd.n14052 185
R28139 vdd.n13991 vdd.n13990 185
R28140 vdd.n13992 vdd.n13991 185
R28141 vdd.n8628 vdd.n8626 185
R28142 vdd.n8631 vdd.n8628 185
R28143 vdd.n8772 vdd.n8771 185
R28144 vdd.n8772 vdd.n8754 185
R28145 vdd.n8779 vdd.n8777 185
R28146 vdd.n8777 vdd.n8776 185
R28147 vdd.n8820 vdd.n8819 185
R28148 vdd.n8820 vdd.n8801 185
R28149 vdd.n8828 vdd.n8826 185
R28150 vdd.n13669 vdd.n8826 185
R28151 vdd.n13474 vdd.n13473 185
R28152 vdd.n13473 vdd.n8988 185
R28153 vdd.n8996 vdd.n8994 185
R28154 vdd.n8994 vdd.n8992 185
R28155 vdd.n9041 vdd.n9040 185
R28156 vdd.n9041 vdd.n9021 185
R28157 vdd.n9049 vdd.n9047 185
R28158 vdd.n13377 vdd.n9047 185
R28159 vdd.n13248 vdd.n13247 185
R28160 vdd.n13247 vdd.n13246 185
R28161 vdd.n9177 vdd.n9175 185
R28162 vdd.n9178 vdd.n9177 185
R28163 vdd.n13268 vdd.n13267 185
R28164 vdd.n13267 vdd.n13266 185
R28165 vdd.n13269 vdd.n9160 185
R28166 vdd.n13265 vdd.n9160 185
R28167 vdd.n13289 vdd.n13288 185
R28168 vdd.n13288 vdd.n13287 185
R28169 vdd.n9149 vdd.n9148 185
R28170 vdd.n9150 vdd.n9149 185
R28171 vdd.n13302 vdd.n13301 185
R28172 vdd.n13303 vdd.n13302 185
R28173 vdd.n13300 vdd.n9144 185
R28174 vdd.n9144 vdd.n9142 185
R28175 vdd.n13338 vdd.n13337 185
R28176 vdd.n13337 vdd.n13336 185
R28177 vdd.n9102 vdd.n9101 185
R28178 vdd.n9103 vdd.n9102 185
R28179 vdd.n13347 vdd.n13346 185
R28180 vdd.n13348 vdd.n13347 185
R28181 vdd.n13345 vdd.n9096 185
R28182 vdd.n9096 vdd.n9094 185
R28183 vdd.n13368 vdd.n13367 185
R28184 vdd.n13367 vdd.n13366 185
R28185 vdd.n9068 vdd.n9067 185
R28186 vdd.n9070 vdd.n9068 185
R28187 vdd.n13358 vdd.n13357 185
R28188 vdd.n13359 vdd.n13358 185
R28189 vdd.n9064 vdd.n9063 185
R28190 vdd.n13355 vdd.n9063 185
R28191 vdd.n13403 vdd.n13402 185
R28192 vdd.n13404 vdd.n13403 185
R28193 vdd.n9054 vdd.n9051 185
R28194 vdd.n9055 vdd.n9054 185
R28195 vdd.n9053 vdd.n9052 185
R28196 vdd.n13390 vdd.n9053 185
R28197 vdd.n13412 vdd.n13411 185
R28198 vdd.n13411 vdd.n13410 185
R28199 vdd.n13425 vdd.n13424 185
R28200 vdd.n13426 vdd.n13425 185
R28201 vdd.n13423 vdd.n9035 185
R28202 vdd.n9035 vdd.n9033 185
R28203 vdd.n13491 vdd.n13490 185
R28204 vdd.n13492 vdd.n13491 185
R28205 vdd.n13484 vdd.n13483 185
R28206 vdd.n13483 vdd.n13482 185
R28207 vdd.n9001 vdd.n9000 185
R28208 vdd.n13481 vdd.n9001 185
R28209 vdd.n8987 vdd.n8986 185
R28210 vdd.n13498 vdd.n8987 185
R28211 vdd.n8983 vdd.n8982 185
R28212 vdd.n8982 vdd.n8981 185
R28213 vdd.n13508 vdd.n13507 185
R28214 vdd.n13509 vdd.n13508 185
R28215 vdd.n13540 vdd.n13539 185
R28216 vdd.n13539 vdd.n13538 185
R28217 vdd.n8956 vdd.n8955 185
R28218 vdd.n8957 vdd.n8956 185
R28219 vdd.n13560 vdd.n13559 185
R28220 vdd.n13559 vdd.n13558 185
R28221 vdd.n13561 vdd.n8938 185
R28222 vdd.n13557 vdd.n8938 185
R28223 vdd.n13581 vdd.n13580 185
R28224 vdd.n13580 vdd.n13579 185
R28225 vdd.n8928 vdd.n8927 185
R28226 vdd.n8929 vdd.n8928 185
R28227 vdd.n13594 vdd.n13593 185
R28228 vdd.n13595 vdd.n13594 185
R28229 vdd.n13592 vdd.n8923 185
R28230 vdd.n8923 vdd.n8921 185
R28231 vdd.n13630 vdd.n13629 185
R28232 vdd.n13629 vdd.n13628 185
R28233 vdd.n8881 vdd.n8880 185
R28234 vdd.n8882 vdd.n8881 185
R28235 vdd.n13639 vdd.n13638 185
R28236 vdd.n13640 vdd.n13639 185
R28237 vdd.n13637 vdd.n8876 185
R28238 vdd.n8876 vdd.n8874 185
R28239 vdd.n13660 vdd.n13659 185
R28240 vdd.n13659 vdd.n13658 185
R28241 vdd.n8848 vdd.n8847 185
R28242 vdd.n8850 vdd.n8848 185
R28243 vdd.n13650 vdd.n13649 185
R28244 vdd.n13651 vdd.n13650 185
R28245 vdd.n8844 vdd.n8843 185
R28246 vdd.n13647 vdd.n8843 185
R28247 vdd.n13696 vdd.n13695 185
R28248 vdd.n13697 vdd.n13696 185
R28249 vdd.n8834 vdd.n8830 185
R28250 vdd.n8835 vdd.n8834 185
R28251 vdd.n8833 vdd.n8832 185
R28252 vdd.n13682 vdd.n8833 185
R28253 vdd.n13706 vdd.n13705 185
R28254 vdd.n13705 vdd.n13704 185
R28255 vdd.n13717 vdd.n13716 185
R28256 vdd.n13718 vdd.n13717 185
R28257 vdd.n13715 vdd.n8814 185
R28258 vdd.n8814 vdd.n8812 185
R28259 vdd.n13771 vdd.n13770 185
R28260 vdd.n13772 vdd.n13771 185
R28261 vdd.n13764 vdd.n13763 185
R28262 vdd.n13763 vdd.n13762 185
R28263 vdd.n8784 vdd.n8783 185
R28264 vdd.n13761 vdd.n8784 185
R28265 vdd.n13780 vdd.n13779 185
R28266 vdd.n13779 vdd.n13778 185
R28267 vdd.n13790 vdd.n13789 185
R28268 vdd.n13791 vdd.n13790 185
R28269 vdd.n13788 vdd.n8768 185
R28270 vdd.n8768 vdd.n8766 185
R28271 vdd.n13825 vdd.n13824 185
R28272 vdd.n13824 vdd.n13823 185
R28273 vdd.n8737 vdd.n8736 185
R28274 vdd.n13821 vdd.n8737 185
R28275 vdd.n13842 vdd.n13841 185
R28276 vdd.n13841 vdd.n13840 185
R28277 vdd.n13843 vdd.n8720 185
R28278 vdd.n13839 vdd.n8720 185
R28279 vdd.n13849 vdd.n13848 185
R28280 vdd.n13848 vdd.n8707 185
R28281 vdd.n8724 vdd.n8722 185
R28282 vdd.n8722 vdd.n8721 185
R28283 vdd.n13898 vdd.n13897 185
R28284 vdd.n13899 vdd.n13898 185
R28285 vdd.n13896 vdd.n8684 185
R28286 vdd.n8684 vdd.n8682 185
R28287 vdd.n8690 vdd.n8676 185
R28288 vdd.n8694 vdd.n8676 185
R28289 vdd.n8692 vdd.n8691 185
R28290 vdd.n8695 vdd.n8692 185
R28291 vdd.n13906 vdd.n8675 185
R28292 vdd.n13906 vdd.n13905 185
R28293 vdd.n8672 vdd.n8658 185
R28294 vdd.n8658 vdd.n8656 185
R28295 vdd.n8666 vdd.n8665 185
R28296 vdd.n8665 vdd.n8664 185
R28297 vdd.n8660 vdd.n8659 185
R28298 vdd.n8663 vdd.n8659 185
R28299 vdd.n13966 vdd.n13965 185
R28300 vdd.n13967 vdd.n13966 185
R28301 vdd.n13964 vdd.n8623 185
R28302 vdd.n8623 vdd.n8621 185
R28303 vdd.n8625 vdd.n8612 185
R28304 vdd.n13974 vdd.n8612 185
R28305 vdd.n13980 vdd.n13979 185
R28306 vdd.n13979 vdd.n8593 185
R28307 vdd.n13978 vdd.n8611 185
R28308 vdd.n13978 vdd.n8594 185
R28309 vdd.n13989 vdd.n8603 185
R28310 vdd.n8603 vdd.n8600 185
R28311 vdd.n8568 vdd.n8566 185
R28312 vdd.n8566 vdd.n8564 185
R28313 vdd.n14061 vdd.n14060 185
R28314 vdd.n14062 vdd.n14061 185
R28315 vdd.n8573 vdd.n8572 185
R28316 vdd.n14051 vdd.n8573 185
R28317 vdd.n14041 vdd.n14039 185
R28318 vdd.n14039 vdd.n8560 185
R28319 vdd.n14040 vdd.n8558 185
R28320 vdd.n14068 vdd.n8558 185
R28321 vdd.n8554 vdd.n8553 185
R28322 vdd.n8553 vdd.n8552 185
R28323 vdd.n8515 vdd.n8513 185
R28324 vdd.n8513 vdd.n8512 185
R28325 vdd.n14117 vdd.n14116 185
R28326 vdd.n14118 vdd.n14117 185
R28327 vdd.n14128 vdd.n8507 185
R28328 vdd.n14128 vdd.n14127 185
R28329 vdd.n8521 vdd.n8506 185
R28330 vdd.n14125 vdd.n8506 185
R28331 vdd.n14131 vdd.n14130 185
R28332 vdd.n14130 vdd.n8490 185
R28333 vdd.n14132 vdd.n8499 185
R28334 vdd.n8499 vdd.n8498 185
R28335 vdd.n14138 vdd.n14137 185
R28336 vdd.n14137 vdd.n8484 185
R28337 vdd.n8503 vdd.n8501 185
R28338 vdd.n8501 vdd.n8500 185
R28339 vdd.n14187 vdd.n14186 185
R28340 vdd.n14188 vdd.n14187 185
R28341 vdd.n14185 vdd.n8460 185
R28342 vdd.n8460 vdd.n8458 185
R28343 vdd.n8467 vdd.n8452 185
R28344 vdd.n8471 vdd.n8452 185
R28345 vdd.n8469 vdd.n8468 185
R28346 vdd.n8472 vdd.n8469 185
R28347 vdd.n14196 vdd.n8451 185
R28348 vdd.n14196 vdd.n14195 185
R28349 vdd.n8448 vdd.n8437 185
R28350 vdd.n14194 vdd.n8437 185
R28351 vdd.n8443 vdd.n8442 185
R28352 vdd.n8442 vdd.n8420 185
R28353 vdd.n8440 vdd.n8439 185
R28354 vdd.n8439 vdd.n8438 185
R28355 vdd.n14256 vdd.n14255 185
R28356 vdd.n14257 vdd.n14256 185
R28357 vdd.n14254 vdd.n8401 185
R28358 vdd.n8401 vdd.n8399 185
R28359 vdd.n8403 vdd.n8390 185
R28360 vdd.n14264 vdd.n8390 185
R28361 vdd.n14270 vdd.n14269 185
R28362 vdd.n14269 vdd.n8371 185
R28363 vdd.n14268 vdd.n8389 185
R28364 vdd.n14268 vdd.n8372 185
R28365 vdd.n14280 vdd.n8381 185
R28366 vdd.n8381 vdd.n8378 185
R28367 vdd.n8350 vdd.n8348 185
R28368 vdd.n8348 vdd.n8346 185
R28369 vdd.n14336 vdd.n14335 185
R28370 vdd.n14337 vdd.n14336 185
R28371 vdd.n8356 vdd.n8355 185
R28372 vdd.n14326 vdd.n8356 185
R28373 vdd.n8341 vdd.n8340 185
R28374 vdd.n8341 vdd.n8318 185
R28375 vdd.n14347 vdd.n14346 185
R28376 vdd.n14346 vdd.n14345 185
R28377 vdd.n14357 vdd.n8335 185
R28378 vdd.n8335 vdd.n8333 185
R28379 vdd.n8302 vdd.n8301 185
R28380 vdd.n8303 vdd.n8302 185
R28381 vdd.n14398 vdd.n14397 185
R28382 vdd.n14397 vdd.n14396 185
R28383 vdd.n14427 vdd.n8276 185
R28384 vdd.n8276 vdd.n8274 185
R28385 vdd.n14429 vdd.n14428 185
R28386 vdd.n14430 vdd.n14429 185
R28387 vdd.n8284 vdd.n8283 185
R28388 vdd.n8287 vdd.n8284 185
R28389 vdd.n8282 vdd.n8242 185
R28390 vdd.n8286 vdd.n8242 185
R28391 vdd.n8251 vdd.n8248 185
R28392 vdd.n14438 vdd.n8251 185
R28393 vdd.n8245 vdd.n8243 185
R28394 vdd.n14437 vdd.n8243 185
R28395 vdd.n8252 vdd.n8249 185
R28396 vdd.n8262 vdd.n8252 185
R28397 vdd.n8260 vdd.n8259 185
R28398 vdd.n8261 vdd.n8260 185
R28399 vdd.n14490 vdd.n14489 185
R28400 vdd.n14489 vdd.n14488 185
R28401 vdd.n8221 vdd.n8220 185
R28402 vdd.n8222 vdd.n8221 185
R28403 vdd.n14499 vdd.n14498 185
R28404 vdd.n14500 vdd.n14499 185
R28405 vdd.n14497 vdd.n8211 185
R28406 vdd.n8216 vdd.n8211 185
R28407 vdd.n13179 vdd.n13178 185
R28408 vdd.n13178 vdd.n13177 185
R28409 vdd.n9216 vdd.n9214 185
R28410 vdd.n9214 vdd.n9212 185
R28411 vdd.n9272 vdd.n9271 185
R28412 vdd.n9272 vdd.n9245 185
R28413 vdd.n13120 vdd.n13119 185
R28414 vdd.n13119 vdd.n13118 185
R28415 vdd.n13131 vdd.n13130 185
R28416 vdd.n13132 vdd.n13131 185
R28417 vdd.n13129 vdd.n9266 185
R28418 vdd.n9266 vdd.n9264 185
R28419 vdd.n13197 vdd.n13196 185
R28420 vdd.n13198 vdd.n13197 185
R28421 vdd.n13190 vdd.n13189 185
R28422 vdd.n13189 vdd.n13188 185
R28423 vdd.n9221 vdd.n9220 185
R28424 vdd.n13187 vdd.n9221 185
R28425 vdd.n9208 vdd.n9206 185
R28426 vdd.n13204 vdd.n9208 185
R28427 vdd.n9204 vdd.n9203 185
R28428 vdd.n9203 vdd.n9191 185
R28429 vdd.n13215 vdd.n13214 185
R28430 vdd.n13216 vdd.n13215 185
R28431 vdd.n13144 vdd.n13143 185
R28432 vdd.n13145 vdd.n13144 185
R28433 vdd.n13142 vdd.n9247 185
R28434 vdd.n9247 vdd.n9245 185
R28435 vdd.n14613 vdd.n14612 185
R28436 vdd.n14614 vdd.n14613 185
R28437 vdd.n8180 vdd.n8179 185
R28438 vdd.n14566 vdd.n8180 185
R28439 vdd.n14539 vdd.n14538 185
R28440 vdd.n14548 vdd.n14539 185
R28441 vdd.n14558 vdd.n14557 185
R28442 vdd.n14559 vdd.n14558 185
R28443 vdd.n8196 vdd.n8194 185
R28444 vdd.n8197 vdd.n8196 185
R28445 vdd.n14484 vdd.n8226 185
R28446 vdd.n8226 vdd.n8224 185
R28447 vdd.n14470 vdd.n14469 185
R28448 vdd.n14469 vdd.n14468 185
R28449 vdd.n8264 vdd.n8263 185
R28450 vdd.n14439 vdd.n8263 185
R28451 vdd.n14413 vdd.n8240 185
R28452 vdd.n14461 vdd.n8240 185
R28453 vdd.n8296 vdd.n8294 185
R28454 vdd.n8296 vdd.n8273 185
R28455 vdd.n8308 vdd.n8306 185
R28456 vdd.n8306 vdd.n8297 185
R28457 vdd.n14383 vdd.n14382 185
R28458 vdd.n14382 vdd.n14381 185
R28459 vdd.n8326 vdd.n8325 185
R28460 vdd.n14361 vdd.n8326 185
R28461 vdd.n14371 vdd.n14370 185
R28462 vdd.n14372 vdd.n14371 185
R28463 vdd.n8359 vdd.n8358 185
R28464 vdd.n8358 vdd.n8357 185
R28465 vdd.n8364 vdd.n8363 185
R28466 vdd.n14301 vdd.n8363 185
R28467 vdd.n14286 vdd.n14285 185
R28468 vdd.n14285 vdd.n14284 185
R28469 vdd.n14242 vdd.n14241 185
R28470 vdd.n14241 vdd.n8392 185
R28471 vdd.n8412 vdd.n8409 185
R28472 vdd.n8409 vdd.n8407 185
R28473 vdd.n8419 vdd.n8415 185
R28474 vdd.n14224 vdd.n8419 185
R28475 vdd.n8435 vdd.n8434 185
R28476 vdd.n14206 vdd.n8435 185
R28477 vdd.n14216 vdd.n14215 185
R28478 vdd.n14217 vdd.n14216 185
R28479 vdd.n8474 vdd.n8473 185
R28480 vdd.n8473 vdd.n8470 185
R28481 vdd.n8480 vdd.n8479 185
R28482 vdd.n14159 vdd.n8479 185
R28483 vdd.n14147 vdd.n14146 185
R28484 vdd.n14146 vdd.n14145 185
R28485 vdd.n14104 vdd.n8527 185
R28486 vdd.n8527 vdd.n8525 185
R28487 vdd.n8534 vdd.n8532 185
R28488 vdd.n14096 vdd.n8534 185
R28489 vdd.n8551 vdd.n8550 185
R28490 vdd.n14079 vdd.n8551 185
R28491 vdd.n14089 vdd.n14088 185
R28492 vdd.n14090 vdd.n14089 185
R28493 vdd.n8579 vdd.n8577 185
R28494 vdd.n8577 vdd.n8576 185
R28495 vdd.n14024 vdd.n14023 185
R28496 vdd.n14023 vdd.n8574 185
R28497 vdd.n8583 vdd.n8582 185
R28498 vdd.n14011 vdd.n8582 185
R28499 vdd.n13995 vdd.n13994 185
R28500 vdd.n13994 vdd.n13993 185
R28501 vdd.n13952 vdd.n13951 185
R28502 vdd.n13951 vdd.n8614 185
R28503 vdd.n8634 vdd.n8630 185
R28504 vdd.n8630 vdd.n8629 185
R28505 vdd.n8641 vdd.n8637 185
R28506 vdd.n13934 vdd.n8641 185
R28507 vdd.n8655 vdd.n8654 185
R28508 vdd.n13916 vdd.n8655 185
R28509 vdd.n13926 vdd.n13925 185
R28510 vdd.n13927 vdd.n13926 185
R28511 vdd.n8697 vdd.n8696 185
R28512 vdd.n8696 vdd.n8693 185
R28513 vdd.n8703 vdd.n8702 185
R28514 vdd.n13870 vdd.n8702 185
R28515 vdd.n13858 vdd.n13857 185
R28516 vdd.n13857 vdd.n13856 185
R28517 vdd.n13819 vdd.n13818 185
R28518 vdd.n13820 vdd.n13819 185
R28519 vdd.n8748 vdd.n8744 185
R28520 vdd.n13809 vdd.n8748 185
R28521 vdd.n8764 vdd.n8763 185
R28522 vdd.n13792 vdd.n8764 185
R28523 vdd.n13802 vdd.n13801 185
R28524 vdd.n13803 vdd.n13802 185
R28525 vdd.n8787 vdd.n8786 185
R28526 vdd.n8786 vdd.n8785 185
R28527 vdd.n8792 vdd.n8791 185
R28528 vdd.n13736 vdd.n8791 185
R28529 vdd.n8811 vdd.n8810 185
R28530 vdd.n13719 vdd.n8811 185
R28531 vdd.n13729 vdd.n13728 185
R28532 vdd.n13730 vdd.n13729 185
R28533 vdd.n13673 vdd.n13672 185
R28534 vdd.n13672 vdd.n8824 185
R28535 vdd.n8866 vdd.n8857 185
R28536 vdd.n8857 vdd.n8842 185
R28537 vdd.n13654 vdd.n8853 185
R28538 vdd.n8853 vdd.n8851 185
R28539 vdd.n8899 vdd.n8890 185
R28540 vdd.n13619 vdd.n8890 185
R28541 vdd.n13624 vdd.n8886 185
R28542 vdd.n8886 vdd.n8884 185
R28543 vdd.n13607 vdd.n13606 185
R28544 vdd.n13608 vdd.n13607 185
R28545 vdd.n8917 vdd.n8915 185
R28546 vdd.n8930 vdd.n8917 185
R28547 vdd.n13570 vdd.n13569 185
R28548 vdd.n13569 vdd.n13568 185
R28549 vdd.n13533 vdd.n8959 185
R28550 vdd.n13529 vdd.n8959 185
R28551 vdd.n8980 vdd.n8979 185
R28552 vdd.n8980 vdd.n8949 185
R28553 vdd.n13520 vdd.n13519 185
R28554 vdd.n13521 vdd.n13520 185
R28555 vdd.n9007 vdd.n9005 185
R28556 vdd.n9005 vdd.n9004 185
R28557 vdd.n13458 vdd.n13457 185
R28558 vdd.n13457 vdd.n9002 185
R28559 vdd.n9011 vdd.n9010 185
R28560 vdd.n13445 vdd.n9010 185
R28561 vdd.n9031 vdd.n9030 185
R28562 vdd.n13427 vdd.n9031 185
R28563 vdd.n13437 vdd.n13436 185
R28564 vdd.n13438 vdd.n13437 185
R28565 vdd.n13381 vdd.n13380 185
R28566 vdd.n13380 vdd.n9045 185
R28567 vdd.n9086 vdd.n9077 185
R28568 vdd.n9077 vdd.n9062 185
R28569 vdd.n13362 vdd.n9073 185
R28570 vdd.n9073 vdd.n9071 185
R28571 vdd.n9120 vdd.n9111 185
R28572 vdd.n13327 vdd.n9111 185
R28573 vdd.n13332 vdd.n9107 185
R28574 vdd.n9107 vdd.n9105 185
R28575 vdd.n13315 vdd.n13314 185
R28576 vdd.n13316 vdd.n13315 185
R28577 vdd.n9139 vdd.n9137 185
R28578 vdd.n9151 vdd.n9139 185
R28579 vdd.n13278 vdd.n13277 185
R28580 vdd.n13277 vdd.n13276 185
R28581 vdd.n13241 vdd.n9180 185
R28582 vdd.n13237 vdd.n9180 185
R28583 vdd.n9202 vdd.n9201 185
R28584 vdd.n13218 vdd.n9202 185
R28585 vdd.n13228 vdd.n13227 185
R28586 vdd.n13229 vdd.n13228 185
R28587 vdd.n9227 vdd.n9226 185
R28588 vdd.n9226 vdd.n9225 185
R28589 vdd.n13161 vdd.n9233 185
R28590 vdd.n13161 vdd.n9222 185
R28591 vdd.n9235 vdd.n9234 185
R28592 vdd.n13152 vdd.n9234 185
R28593 vdd.n13135 vdd.n13134 185
R28594 vdd.n13134 vdd.n13133 185
R28595 vdd.n14611 vdd.n8168 185
R28596 vdd.n8174 vdd.n8168 185
R28597 vdd.n14541 vdd.n14540 185
R28598 vdd.n14540 vdd.n8183 185
R28599 vdd.n14551 vdd.n14550 185
R28600 vdd.n14550 vdd.n14549 185
R28601 vdd.n8191 vdd.n8189 185
R28602 vdd.n8189 vdd.n8187 185
R28603 vdd.n14481 vdd.n14479 185
R28604 vdd.n14481 vdd.n14480 185
R28605 vdd.n14486 vdd.n14485 185
R28606 vdd.n14487 vdd.n14486 185
R28607 vdd.n8231 vdd.n8230 185
R28608 vdd.n8232 vdd.n8231 185
R28609 vdd.n14442 vdd.n14441 185
R28610 vdd.n14441 vdd.n14440 185
R28611 vdd.n8291 vdd.n8289 185
R28612 vdd.n8289 vdd.n8239 185
R28613 vdd.n8290 vdd.n8288 185
R28614 vdd.n8288 vdd.n8285 185
R28615 vdd.n14388 vdd.n8295 185
R28616 vdd.n14407 vdd.n8295 185
R28617 vdd.n14384 vdd.n8305 185
R28618 vdd.n8305 vdd.n8303 185
R28619 vdd.n8332 vdd.n8331 185
R28620 vdd.n14360 vdd.n8332 185
R28621 vdd.n14369 vdd.n8320 185
R28622 vdd.n8320 vdd.n8318 185
R28623 vdd.n14318 vdd.n14317 185
R28624 vdd.n14327 vdd.n14318 185
R28625 vdd.n14309 vdd.n14308 185
R28626 vdd.n14309 vdd.n8346 185
R28627 vdd.n14287 vdd.n8367 185
R28628 vdd.n14283 vdd.n8367 185
R28629 vdd.n14243 vdd.n8411 185
R28630 vdd.n8411 vdd.n8410 185
R28631 vdd.n14235 vdd.n14234 185
R28632 vdd.n14234 vdd.n14233 185
R28633 vdd.n14227 vdd.n14226 185
R28634 vdd.n14226 vdd.n14225 185
R28635 vdd.n14209 vdd.n14208 185
R28636 vdd.n14208 vdd.n14207 185
R28637 vdd.n8429 vdd.n8427 185
R28638 vdd.n8427 vdd.n8425 185
R28639 vdd.n14170 vdd.n14169 185
R28640 vdd.n14169 vdd.n14168 185
R28641 vdd.n14162 vdd.n14161 185
R28642 vdd.n14161 vdd.n14160 185
R28643 vdd.n8494 vdd.n8492 185
R28644 vdd.n8496 vdd.n8492 185
R28645 vdd.n8493 vdd.n8491 185
R28646 vdd.n14126 vdd.n8491 185
R28647 vdd.n8531 vdd.n8526 185
R28648 vdd.n8526 vdd.n8524 185
R28649 vdd.n8549 vdd.n8533 185
R28650 vdd.n8533 vdd.n8512 185
R28651 vdd.n14087 vdd.n8543 185
R28652 vdd.n8543 vdd.n8541 185
R28653 vdd.n14031 vdd.n14030 185
R28654 vdd.n14030 vdd.n8560 185
R28655 vdd.n14025 vdd.n8575 185
R28656 vdd.n14052 vdd.n8575 185
R28657 vdd.n14020 vdd.n14019 185
R28658 vdd.n14020 vdd.n8564 185
R28659 vdd.n13996 vdd.n8587 185
R28660 vdd.n13992 vdd.n8587 185
R28661 vdd.n13953 vdd.n8633 185
R28662 vdd.n8633 vdd.n8632 185
R28663 vdd.n13945 vdd.n13944 185
R28664 vdd.n13944 vdd.n13943 185
R28665 vdd.n13937 vdd.n13936 185
R28666 vdd.n13936 vdd.n13935 185
R28667 vdd.n13919 vdd.n13918 185
R28668 vdd.n13918 vdd.n13917 185
R28669 vdd.n8649 vdd.n8647 185
R28670 vdd.n8647 vdd.t110 185
R28671 vdd.n13881 vdd.n13880 185
R28672 vdd.n13880 vdd.n13879 185
R28673 vdd.n13873 vdd.n13872 185
R28674 vdd.n13872 vdd.n13871 185
R28675 vdd.n8716 vdd.n8714 185
R28676 vdd.n8718 vdd.n8714 185
R28677 vdd.n8715 vdd.n8713 185
R28678 vdd.n13822 vdd.n8713 185
R28679 vdd.n8747 vdd.n8746 185
R28680 vdd.n8747 vdd.n8731 185
R28681 vdd.n8762 vdd.n8745 185
R28682 vdd.n13791 vdd.n8745 185
R28683 vdd.n13800 vdd.n8756 185
R28684 vdd.n8756 vdd.n8754 185
R28685 vdd.n13754 vdd.n13753 185
R28686 vdd.n13762 vdd.n13754 185
R28687 vdd.n13744 vdd.n13743 185
R28688 vdd.n13744 vdd.n8776 185
R28689 vdd.n8809 vdd.n8795 185
R28690 vdd.n13718 vdd.n8795 185
R28691 vdd.n13727 vdd.n8803 185
R28692 vdd.n8803 vdd.n8801 185
R28693 vdd.n13671 vdd.n8840 185
R28694 vdd.n13671 vdd.n13670 185
R28695 vdd.n8868 vdd.n8867 185
R28696 vdd.n13646 vdd.n8868 185
R28697 vdd.n13656 vdd.n13655 185
R28698 vdd.n13657 vdd.n13656 185
R28699 vdd.n13621 vdd.n8900 185
R28700 vdd.n13621 vdd.n13620 185
R28701 vdd.n13626 vdd.n13625 185
R28702 vdd.n13627 vdd.n13626 185
R28703 vdd.n8912 vdd.n8911 185
R28704 vdd.n8920 vdd.n8911 185
R28705 vdd.n13577 vdd.n13576 185
R28706 vdd.n13578 vdd.n13577 185
R28707 vdd.n8935 vdd.n8934 185
R28708 vdd.n13556 vdd.n8935 185
R28709 vdd.n13536 vdd.n13535 185
R28710 vdd.n13537 vdd.n13536 185
R28711 vdd.n8978 vdd.n8963 185
R28712 vdd.n8963 vdd.n8950 185
R28713 vdd.n13518 vdd.n8971 185
R28714 vdd.n8981 vdd.n8971 185
R28715 vdd.n13465 vdd.n13464 185
R28716 vdd.n13464 vdd.n8988 185
R28717 vdd.n13459 vdd.n9003 185
R28718 vdd.n13482 vdd.n9003 185
R28719 vdd.n13454 vdd.n13453 185
R28720 vdd.n13454 vdd.n8992 185
R28721 vdd.n9029 vdd.n9015 185
R28722 vdd.n13426 vdd.n9015 185
R28723 vdd.n13435 vdd.n9023 185
R28724 vdd.n9023 vdd.n9021 185
R28725 vdd.n13379 vdd.n9060 185
R28726 vdd.n13379 vdd.n13378 185
R28727 vdd.n9088 vdd.n9087 185
R28728 vdd.n13354 vdd.n9088 185
R28729 vdd.n13364 vdd.n13363 185
R28730 vdd.n13365 vdd.n13364 185
R28731 vdd.n13329 vdd.n9121 185
R28732 vdd.n13329 vdd.n13328 185
R28733 vdd.n13334 vdd.n13333 185
R28734 vdd.n13335 vdd.n13334 185
R28735 vdd.n9134 vdd.n9133 185
R28736 vdd.n9133 vdd.n9130 185
R28737 vdd.n13285 vdd.n13284 185
R28738 vdd.n13286 vdd.n13285 185
R28739 vdd.n9156 vdd.n9155 185
R28740 vdd.n9157 vdd.n9156 185
R28741 vdd.n13244 vdd.n13243 185
R28742 vdd.n13245 vdd.n13244 185
R28743 vdd.n9200 vdd.n9184 185
R28744 vdd.n9184 vdd.n9170 185
R28745 vdd.n13226 vdd.n9193 185
R28746 vdd.n9193 vdd.n9191 185
R28747 vdd.n13176 vdd.n13175 185
R28748 vdd.n13177 vdd.n13176 185
R28749 vdd.n9230 vdd.n9223 185
R28750 vdd.n13188 vdd.n9223 185
R28751 vdd.n13160 vdd.n13159 185
R28752 vdd.n13160 vdd.n9212 185
R28753 vdd.n9261 vdd.n9238 185
R28754 vdd.n13132 vdd.n9238 185
R28755 vdd.n11627 vdd.n11626 185
R28756 vdd.n11628 vdd.n11627 185
R28757 vdd.n11579 vdd.n11575 185
R28758 vdd.n11575 vdd.n11567 185
R28759 vdd.n10336 vdd.n10333 185
R28760 vdd.n10392 vdd.n10336 185
R28761 vdd.n10325 vdd.n10324 185
R28762 vdd.n10404 vdd.n10325 185
R28763 vdd.n10414 vdd.n10413 185
R28764 vdd.n10415 vdd.n10414 185
R28765 vdd.n10314 vdd.n10311 185
R28766 vdd.n10319 vdd.n10314 185
R28767 vdd.n10428 vdd.n10427 185
R28768 vdd.n10429 vdd.n10428 185
R28769 vdd.n10438 vdd.n10298 185
R28770 vdd.n10298 vdd.n10297 185
R28771 vdd.n10457 vdd.n10456 185
R28772 vdd.n10456 vdd.n10455 185
R28773 vdd.n10281 vdd.n10278 185
R28774 vdd.n10466 vdd.n10278 185
R28775 vdd.n10471 vdd.n10273 185
R28776 vdd.n10276 vdd.n10273 185
R28777 vdd.n10478 vdd.n10477 185
R28778 vdd.n10151 vdd.n10037 185
R28779 vdd.t299 vdd.n10037 185
R28780 vdd.n10033 vdd.n10030 185
R28781 vdd.n10038 vdd.n10030 185
R28782 vdd.n12647 vdd.n12646 185
R28783 vdd.n12646 vdd.n12645 185
R28784 vdd.n10020 vdd.n10017 185
R28785 vdd.n12656 vdd.n10017 185
R28786 vdd.n12663 vdd.n12662 185
R28787 vdd.n12664 vdd.n12663 185
R28788 vdd.n9989 vdd.n9988 185
R28789 vdd.n10008 vdd.n9989 185
R28790 vdd.n9997 vdd.n9996 185
R28791 vdd.n9996 vdd.n9975 185
R28792 vdd.n12676 vdd.n9971 185
R28793 vdd.n9974 vdd.n9971 185
R28794 vdd.n12678 vdd.n12677 185
R28795 vdd.n12679 vdd.n12678 185
R28796 vdd.n9966 vdd.n9964 185
R28797 vdd.n9968 vdd.n9966 185
R28798 vdd.n9959 vdd.n9931 185
R28799 vdd.n9931 vdd.n9929 185
R28800 vdd.n9952 vdd.n9951 185
R28801 vdd.n9953 vdd.n9952 185
R28802 vdd.n12699 vdd.n9919 185
R28803 vdd.n12699 vdd.n12698 185
R28804 vdd.n12708 vdd.n12707 185
R28805 vdd.n12709 vdd.n12708 185
R28806 vdd.n9912 vdd.n9909 185
R28807 vdd.n9914 vdd.n9912 185
R28808 vdd.n9904 vdd.n9887 185
R28809 vdd.n9887 vdd.n9885 185
R28810 vdd.n9870 vdd.n9867 185
R28811 vdd.n12739 vdd.n9867 185
R28812 vdd.n12746 vdd.n12745 185
R28813 vdd.n12747 vdd.n12746 185
R28814 vdd.n9842 vdd.n9841 185
R28815 vdd.n9858 vdd.n9842 185
R28816 vdd.n9847 vdd.n9823 185
R28817 vdd.n9826 vdd.n9823 185
R28818 vdd.n9819 vdd.n9816 185
R28819 vdd.n9824 vdd.n9816 185
R28820 vdd.n12768 vdd.n12767 185
R28821 vdd.n12767 vdd.n12766 185
R28822 vdd.n9783 vdd.n9781 185
R28823 vdd.n12777 vdd.n9781 185
R28824 vdd.n12784 vdd.n12783 185
R28825 vdd.n12785 vdd.n12784 185
R28826 vdd.n9779 vdd.n9777 185
R28827 vdd.n9777 vdd.n9775 185
R28828 vdd.n9803 vdd.n9802 185
R28829 vdd.n9802 vdd.n9801 185
R28830 vdd.n12794 vdd.n9765 185
R28831 vdd.n12794 vdd.n12793 185
R28832 vdd.n12803 vdd.n12802 185
R28833 vdd.n12804 vdd.n12803 185
R28834 vdd.n9757 vdd.n9754 185
R28835 vdd.n9759 vdd.n9757 185
R28836 vdd.n9749 vdd.n9721 185
R28837 vdd.n9721 vdd.n9719 185
R28838 vdd.n9742 vdd.n9741 185
R28839 vdd.n9743 vdd.n9742 185
R28840 vdd.n9713 vdd.n9712 185
R28841 vdd.n12823 vdd.n9713 185
R28842 vdd.n9696 vdd.n9677 185
R28843 vdd.n9680 vdd.n9677 185
R28844 vdd.n9673 vdd.n9670 185
R28845 vdd.n9678 vdd.n9670 185
R28846 vdd.n12855 vdd.n12854 185
R28847 vdd.n12854 vdd.n12853 185
R28848 vdd.n9660 vdd.n9657 185
R28849 vdd.n12864 vdd.n9657 185
R28850 vdd.n12871 vdd.n12870 185
R28851 vdd.n12872 vdd.n12871 185
R28852 vdd.n9629 vdd.n9628 185
R28853 vdd.n9648 vdd.n9629 185
R28854 vdd.n9637 vdd.n9636 185
R28855 vdd.n9636 vdd.n9615 185
R28856 vdd.n12884 vdd.n9611 185
R28857 vdd.n9614 vdd.n9611 185
R28858 vdd.n12886 vdd.n12885 185
R28859 vdd.n12887 vdd.n12886 185
R28860 vdd.n9606 vdd.n9604 185
R28861 vdd.n9608 vdd.n9606 185
R28862 vdd.n9599 vdd.n9572 185
R28863 vdd.n9572 vdd.n9570 185
R28864 vdd.n9592 vdd.n9591 185
R28865 vdd.n9593 vdd.n9592 185
R28866 vdd.n12907 vdd.n9560 185
R28867 vdd.n12907 vdd.n12906 185
R28868 vdd.n12916 vdd.n12915 185
R28869 vdd.n12917 vdd.n12916 185
R28870 vdd.n9552 vdd.n9549 185
R28871 vdd.n9554 vdd.n9552 185
R28872 vdd.n9544 vdd.n9526 185
R28873 vdd.n9540 vdd.n9526 185
R28874 vdd.n9510 vdd.n9507 185
R28875 vdd.n12947 vdd.n9507 185
R28876 vdd.n12954 vdd.n12953 185
R28877 vdd.n12955 vdd.n12954 185
R28878 vdd.n9482 vdd.n9481 185
R28879 vdd.n9498 vdd.n9482 185
R28880 vdd.n9487 vdd.n9463 185
R28881 vdd.n9466 vdd.n9463 185
R28882 vdd.n9459 vdd.n9456 185
R28883 vdd.n9464 vdd.n9456 185
R28884 vdd.n12976 vdd.n12975 185
R28885 vdd.n12975 vdd.n12974 185
R28886 vdd.n9423 vdd.n9420 185
R28887 vdd.n12985 vdd.n9420 185
R28888 vdd.n12992 vdd.n12991 185
R28889 vdd.n12993 vdd.n12992 185
R28890 vdd.n9418 vdd.n9416 185
R28891 vdd.n9416 vdd.n9414 185
R28892 vdd.n9444 vdd.n9443 185
R28893 vdd.n9443 vdd.n9442 185
R28894 vdd.n13002 vdd.n9405 185
R28895 vdd.n13002 vdd.n13001 185
R28896 vdd.n13011 vdd.n13010 185
R28897 vdd.n13012 vdd.n13011 185
R28898 vdd.n9397 vdd.n9394 185
R28899 vdd.n9399 vdd.n9397 185
R28900 vdd.n9389 vdd.n9361 185
R28901 vdd.n9361 vdd.n9359 185
R28902 vdd.n9382 vdd.n9381 185
R28903 vdd.n9383 vdd.n9382 185
R28904 vdd.n9353 vdd.n9352 185
R28905 vdd.n13031 vdd.n9353 185
R28906 vdd.n9336 vdd.n9316 185
R28907 vdd.n9318 vdd.n9316 185
R28908 vdd.n9312 vdd.n9309 185
R28909 vdd.n9319 vdd.n9309 185
R28910 vdd.n13063 vdd.n13062 185
R28911 vdd.n13062 vdd.n13061 185
R28912 vdd.n9300 vdd.n9296 185
R28913 vdd.n13072 vdd.n9296 185
R28914 vdd.n13079 vdd.n13078 185
R28915 vdd.n13080 vdd.n13079 185
R28916 vdd.n10358 vdd.n10356 185
R28917 vdd.n10369 vdd.n10356 185
R28918 vdd.n10351 vdd.n10345 185
R28919 vdd.n10345 vdd.n10344 185
R28920 vdd.n10383 vdd.n10382 185
R28921 vdd.n10382 vdd.n10381 185
R28922 vdd.n10384 vdd.n10340 185
R28923 vdd.n10340 vdd.n10339 185
R28924 vdd.n10390 vdd.n10338 185
R28925 vdd.n10055 vdd.n10054 185
R28926 vdd.n12614 vdd.n10055 185
R28927 vdd.n10187 vdd.n10186 185
R28928 vdd.n10188 vdd.n10187 185
R28929 vdd.n10137 vdd.n10063 185
R28930 vdd.n10063 vdd.n10061 185
R28931 vdd.n12602 vdd.n10064 185
R28932 vdd.n10105 vdd.n10064 185
R28933 vdd.n10110 vdd.n10097 185
R28934 vdd.n10111 vdd.n10110 185
R28935 vdd.n10101 vdd.n10100 185
R28936 vdd.t83 vdd.n10101 185
R28937 vdd.n10246 vdd.n10245 185
R28938 vdd.n10245 vdd.n10244 185
R28939 vdd.n10122 vdd.n10120 185
R28940 vdd.n10120 vdd.n10118 185
R28941 vdd.n10481 vdd.n10123 185
R28942 vdd.n10486 vdd.n10481 185
R28943 vdd.n10492 vdd.n10491 185
R28944 vdd.n10493 vdd.n10492 185
R28945 vdd.n12586 vdd.n12585 185
R28946 vdd.n12587 vdd.n12586 185
R28947 vdd.n10109 vdd.n10066 185
R28948 vdd.n11936 vdd.n11550 185
R28949 vdd.n11550 vdd.n11549 185
R28950 vdd.n11948 vdd.n11947 185
R28951 vdd.n11947 vdd.n11946 185
R28952 vdd.n11448 vdd.n11446 185
R28953 vdd.n11446 vdd.n11444 185
R28954 vdd.n11524 vdd.n11457 185
R28955 vdd.n11526 vdd.n11524 185
R28956 vdd.n11505 vdd.n11436 185
R28957 vdd.n11964 vdd.n11436 185
R28958 vdd.n11970 vdd.n11969 185
R28959 vdd.n11971 vdd.n11970 185
R28960 vdd.n11976 vdd.n11427 185
R28961 vdd.n11427 vdd.n11426 185
R28962 vdd.n11978 vdd.n11977 185
R28963 vdd.n11979 vdd.n11978 185
R28964 vdd.n11485 vdd.n11484 185
R28965 vdd.n11484 vdd.n11424 185
R28966 vdd.n11474 vdd.n11472 185
R28967 vdd.n11472 vdd.n11414 185
R28968 vdd.n11412 vdd.n11409 185
R28969 vdd.n11415 vdd.n11412 185
R28970 vdd.n11998 vdd.n11997 185
R28971 vdd.n11999 vdd.n11998 185
R28972 vdd.n12008 vdd.n11378 185
R28973 vdd.n11378 vdd.n11376 185
R28974 vdd.n11397 vdd.n11396 185
R28975 vdd.n11396 vdd.n11395 185
R28976 vdd.n11386 vdd.n11384 185
R28977 vdd.n11384 vdd.n11371 185
R28978 vdd.n11365 vdd.n11362 185
R28979 vdd.n11370 vdd.n11365 185
R28980 vdd.n11352 vdd.n11340 185
R28981 vdd.n11353 vdd.n11352 185
R28982 vdd.n11343 vdd.n11324 185
R28983 vdd.n12036 vdd.n11324 185
R28984 vdd.n11320 vdd.n11317 185
R28985 vdd.n11317 vdd.n11316 185
R28986 vdd.n12050 vdd.n12049 185
R28987 vdd.n12049 vdd.n12048 185
R28988 vdd.n11285 vdd.n11283 185
R28989 vdd.n11283 vdd.n11281 185
R28990 vdd.n11304 vdd.n11303 185
R28991 vdd.n11305 vdd.n11304 185
R28992 vdd.n11296 vdd.n11272 185
R28993 vdd.n12065 vdd.n11272 185
R28994 vdd.n12071 vdd.n12070 185
R28995 vdd.n12072 vdd.n12071 185
R28996 vdd.n11269 vdd.n11268 185
R28997 vdd.n12073 vdd.n11269 185
R28998 vdd.n12081 vdd.n11243 185
R28999 vdd.n11243 vdd.n11241 185
R29000 vdd.n11262 vdd.n11261 185
R29001 vdd.n11261 vdd.n11260 185
R29002 vdd.n11251 vdd.n11249 185
R29003 vdd.n11249 vdd.n11231 185
R29004 vdd.n11228 vdd.n11225 185
R29005 vdd.n11230 vdd.n11228 185
R29006 vdd.n12102 vdd.n12101 185
R29007 vdd.n12103 vdd.n12102 185
R29008 vdd.n12112 vdd.n11194 185
R29009 vdd.n11194 vdd.n11192 185
R29010 vdd.n11213 vdd.n11212 185
R29011 vdd.n11212 vdd.n11211 185
R29012 vdd.n11202 vdd.n11200 185
R29013 vdd.n11200 vdd.n11185 185
R29014 vdd.n12136 vdd.n12135 185
R29015 vdd.n12135 vdd.n12134 185
R29016 vdd.n11149 vdd.n11147 185
R29017 vdd.n11147 vdd.n11145 185
R29018 vdd.n11167 vdd.n11166 185
R29019 vdd.n11168 vdd.n11167 185
R29020 vdd.n11159 vdd.n11136 185
R29021 vdd.n12151 vdd.n11136 185
R29022 vdd.n11132 vdd.n11129 185
R29023 vdd.n11129 vdd.n11128 185
R29024 vdd.n12165 vdd.n12164 185
R29025 vdd.n12164 vdd.n12163 185
R29026 vdd.n11109 vdd.n11107 185
R29027 vdd.n11107 vdd.n11105 185
R29028 vdd.n11116 vdd.n11115 185
R29029 vdd.n11117 vdd.n11116 185
R29030 vdd.n11094 vdd.n11092 185
R29031 vdd.n11096 vdd.n11094 185
R29032 vdd.n11093 vdd.n11090 185
R29033 vdd.n11095 vdd.n11093 185
R29034 vdd.n12190 vdd.n12189 185
R29035 vdd.n12191 vdd.n12190 185
R29036 vdd.n12200 vdd.n11059 185
R29037 vdd.n11059 vdd.n11057 185
R29038 vdd.n11078 vdd.n11077 185
R29039 vdd.n11077 vdd.n11076 185
R29040 vdd.n11067 vdd.n11065 185
R29041 vdd.n11065 vdd.n11046 185
R29042 vdd.n11043 vdd.n11040 185
R29043 vdd.n11045 vdd.n11043 185
R29044 vdd.n12221 vdd.n12220 185
R29045 vdd.n12222 vdd.n12221 185
R29046 vdd.n12231 vdd.n11014 185
R29047 vdd.n11014 vdd.n11012 185
R29048 vdd.n11021 vdd.n11002 185
R29049 vdd.n12241 vdd.n11002 185
R29050 vdd.n10998 vdd.n10995 185
R29051 vdd.n10995 vdd.n10994 185
R29052 vdd.n12255 vdd.n12254 185
R29053 vdd.n12254 vdd.n12253 185
R29054 vdd.n10963 vdd.n10961 185
R29055 vdd.n10961 vdd.n10959 185
R29056 vdd.n10982 vdd.n10981 185
R29057 vdd.n10983 vdd.n10982 185
R29058 vdd.n10974 vdd.n10951 185
R29059 vdd.n12270 vdd.n10951 185
R29060 vdd.n12276 vdd.n12275 185
R29061 vdd.n12277 vdd.n12276 185
R29062 vdd.n12282 vdd.n10918 185
R29063 vdd.n10918 vdd.n10917 185
R29064 vdd.n12284 vdd.n12283 185
R29065 vdd.n12285 vdd.n12284 185
R29066 vdd.n10941 vdd.n10940 185
R29067 vdd.n10940 vdd.n10915 185
R29068 vdd.n10930 vdd.n10928 185
R29069 vdd.n10928 vdd.n10906 185
R29070 vdd.n10903 vdd.n10900 185
R29071 vdd.n10905 vdd.n10903 185
R29072 vdd.n12304 vdd.n12303 185
R29073 vdd.n12305 vdd.n12304 185
R29074 vdd.n12314 vdd.n10869 185
R29075 vdd.n10869 vdd.n10867 185
R29076 vdd.n10888 vdd.n10887 185
R29077 vdd.n10887 vdd.n10886 185
R29078 vdd.n10877 vdd.n10875 185
R29079 vdd.n10875 vdd.n10862 185
R29080 vdd.n10856 vdd.n10853 185
R29081 vdd.n10861 vdd.n10856 185
R29082 vdd.n10843 vdd.n10831 185
R29083 vdd.n10844 vdd.n10843 185
R29084 vdd.n10834 vdd.n10815 185
R29085 vdd.n12342 vdd.n10815 185
R29086 vdd.n10811 vdd.n10808 185
R29087 vdd.n10808 vdd.n10807 185
R29088 vdd.n12356 vdd.n12355 185
R29089 vdd.n12355 vdd.n12354 185
R29090 vdd.n10777 vdd.n10775 185
R29091 vdd.n10775 vdd.n10773 185
R29092 vdd.n10795 vdd.n10794 185
R29093 vdd.n10796 vdd.n10795 185
R29094 vdd.n10787 vdd.n10756 185
R29095 vdd.n12371 vdd.n10756 185
R29096 vdd.n10761 vdd.n10760 185
R29097 vdd.n10762 vdd.n10761 185
R29098 vdd.n10759 vdd.n10758 185
R29099 vdd.n10758 vdd.n10757 185
R29100 vdd.n12381 vdd.n12380 185
R29101 vdd.n12382 vdd.n12381 185
R29102 vdd.n12391 vdd.n10722 185
R29103 vdd.n10722 vdd.n10720 185
R29104 vdd.n10741 vdd.n10740 185
R29105 vdd.n10740 vdd.n10739 185
R29106 vdd.n10730 vdd.n10728 185
R29107 vdd.n10728 vdd.n10709 185
R29108 vdd.n10706 vdd.n10703 185
R29109 vdd.n10708 vdd.n10706 185
R29110 vdd.n12412 vdd.n12411 185
R29111 vdd.n12413 vdd.n12412 185
R29112 vdd.n12422 vdd.n10674 185
R29113 vdd.n10674 vdd.n10672 185
R29114 vdd.n10692 vdd.n10691 185
R29115 vdd.n10691 vdd.n10690 185
R29116 vdd.n10660 vdd.n10657 185
R29117 vdd.n10657 vdd.n10656 185
R29118 vdd.n12445 vdd.n12444 185
R29119 vdd.n12444 vdd.n12443 185
R29120 vdd.n10626 vdd.n10624 185
R29121 vdd.n10624 vdd.n10622 185
R29122 vdd.n10644 vdd.n10643 185
R29123 vdd.n10645 vdd.n10644 185
R29124 vdd.n10636 vdd.n10613 185
R29125 vdd.n12460 vdd.n10613 185
R29126 vdd.n10609 vdd.n10606 185
R29127 vdd.n10606 vdd.n10605 185
R29128 vdd.n12474 vdd.n12473 185
R29129 vdd.n12473 vdd.n12472 185
R29130 vdd.n10587 vdd.n10585 185
R29131 vdd.n10585 vdd.n10583 185
R29132 vdd.n10596 vdd.n10591 185
R29133 vdd.n10597 vdd.n10596 185
R29134 vdd.n10595 vdd.n10594 185
R29135 vdd.n10595 vdd.n10574 185
R29136 vdd.n10571 vdd.n10568 185
R29137 vdd.n10573 vdd.n10571 185
R29138 vdd.n12500 vdd.n12499 185
R29139 vdd.n12501 vdd.n12500 185
R29140 vdd.n12510 vdd.n10531 185
R29141 vdd.n10531 vdd.n10529 185
R29142 vdd.n10556 vdd.n10555 185
R29143 vdd.n10555 vdd.n10554 185
R29144 vdd.n10545 vdd.n10537 185
R29145 vdd.n10537 vdd.n10523 185
R29146 vdd.n12523 vdd.n12522 185
R29147 vdd.n12522 vdd.n12521 185
R29148 vdd.n11922 vdd.n11566 185
R29149 vdd.n11566 vdd.n11565 185
R29150 vdd.n22139 vdd.n22138 185
R29151 vdd.n22197 vdd.n22196 185
R29152 vdd.n22201 vdd.n22200 185
R29153 vdd.n22206 vdd.n22205 185
R29154 vdd.n22211 vdd.n22210 185
R29155 vdd.n22237 vdd.n22236 185
R29156 vdd.n22337 vdd.n22336 185
R29157 vdd.n22055 vdd.n22054 185
R29158 vdd.n22059 vdd.n22058 185
R29159 vdd.n22070 vdd.n22069 185
R29160 vdd.n22075 vdd.n22074 185
R29161 vdd.n22113 vdd.n22112 185
R29162 vdd.n11824 vdd.n11817 183.59
R29163 vdd.n21915 vdd.n21908 183.59
R29164 vdd.n11740 vdd.n11729 183.477
R29165 vdd.n11738 vdd.n11730 174.534
R29166 vdd.n11822 vdd.n11813 174.534
R29167 vdd.n21818 vdd.n21817 174.534
R29168 vdd.n21913 vdd.n21904 174.534
R29169 vdd.n14504 vdd.n8198 133.655
R29170 vdd.n13116 vdd.n9211 133.655
R29171 vdd.n13199 vdd.n9211 133.655
R29172 vdd.n13199 vdd.n9209 133.655
R29173 vdd.n13203 vdd.n9209 133.655
R29174 vdd.n13203 vdd.n9169 133.655
R29175 vdd.n13258 vdd.n9169 133.655
R29176 vdd.n13258 vdd.n9166 133.655
R29177 vdd.n13264 vdd.n9166 133.655
R29178 vdd.n13264 vdd.n9167 133.655
R29179 vdd.n9167 vdd.n9141 133.655
R29180 vdd.n9141 vdd.n9092 133.655
R29181 vdd.n13349 vdd.n9092 133.655
R29182 vdd.n13349 vdd.n9090 133.655
R29183 vdd.n13353 vdd.n9090 133.655
R29184 vdd.n13353 vdd.n9044 133.655
R29185 vdd.n13405 vdd.n9044 133.655
R29186 vdd.n13405 vdd.n9042 133.655
R29187 vdd.n13409 vdd.n9042 133.655
R29188 vdd.n13409 vdd.n8991 133.655
R29189 vdd.n13493 vdd.n8991 133.655
R29190 vdd.n13493 vdd.n8989 133.655
R29191 vdd.n13497 vdd.n8989 133.655
R29192 vdd.n13497 vdd.n8948 133.655
R29193 vdd.n13549 vdd.n8948 133.655
R29194 vdd.n13549 vdd.n8945 133.655
R29195 vdd.n13555 vdd.n8945 133.655
R29196 vdd.n13555 vdd.n8946 133.655
R29197 vdd.n8946 vdd.n8919 133.655
R29198 vdd.n8919 vdd.n8872 133.655
R29199 vdd.n13641 vdd.n8872 133.655
R29200 vdd.n13641 vdd.n8870 133.655
R29201 vdd.n13645 vdd.n8870 133.655
R29202 vdd.n13645 vdd.n8823 133.655
R29203 vdd.n13698 vdd.n8823 133.655
R29204 vdd.n13698 vdd.n8821 133.655
R29205 vdd.n13702 vdd.n8821 133.655
R29206 vdd.n13702 vdd.n8775 133.655
R29207 vdd.n13773 vdd.n8775 133.655
R29208 vdd.n13773 vdd.n8773 133.655
R29209 vdd.n13777 vdd.n8773 133.655
R29210 vdd.n13777 vdd.n8730 133.655
R29211 vdd.n13834 vdd.n8730 133.655
R29212 vdd.n13834 vdd.n8728 133.655
R29213 vdd.n13838 vdd.n8728 133.655
R29214 vdd.n13838 vdd.n8680 133.655
R29215 vdd.n13900 vdd.n8680 133.655
R29216 vdd.n13900 vdd.n8678 133.655
R29217 vdd.n13904 vdd.n8678 133.655
R29218 vdd.n13904 vdd.n8618 133.655
R29219 vdd.n13968 vdd.n8618 133.655
R29220 vdd.n13968 vdd.n8615 133.655
R29221 vdd.n13973 vdd.n8615 133.655
R29222 vdd.n13973 vdd.n8616 133.655
R29223 vdd.n8616 vdd.n8563 133.655
R29224 vdd.n14063 vdd.n8563 133.655
R29225 vdd.n14063 vdd.n8561 133.655
R29226 vdd.n14067 vdd.n8561 133.655
R29227 vdd.n14067 vdd.n8511 133.655
R29228 vdd.n14119 vdd.n8511 133.655
R29229 vdd.n14119 vdd.n8508 133.655
R29230 vdd.n14124 vdd.n8508 133.655
R29231 vdd.n14124 vdd.n8509 133.655
R29232 vdd.n8509 vdd.n8456 133.655
R29233 vdd.n14189 vdd.n8456 133.655
R29234 vdd.n14189 vdd.n8454 133.655
R29235 vdd.n14193 vdd.n8454 133.655
R29236 vdd.n14193 vdd.n8396 133.655
R29237 vdd.n14258 vdd.n8396 133.655
R29238 vdd.n14258 vdd.n8393 133.655
R29239 vdd.n14263 vdd.n8393 133.655
R29240 vdd.n14263 vdd.n8394 133.655
R29241 vdd.n8394 vdd.n8345 133.655
R29242 vdd.n14338 vdd.n8345 133.655
R29243 vdd.n14338 vdd.n8342 133.655
R29244 vdd.n14344 vdd.n8342 133.655
R29245 vdd.n14344 vdd.n8343 133.655
R29246 vdd.n8343 vdd.n8304 133.655
R29247 vdd.n8304 vdd.n8272 133.655
R29248 vdd.n14431 vdd.n8272 133.655
R29249 vdd.n14431 vdd.n8269 133.655
R29250 vdd.n14436 vdd.n8269 133.655
R29251 vdd.n14436 vdd.n8270 133.655
R29252 vdd.n8270 vdd.n8214 133.655
R29253 vdd.n14501 vdd.n8214 133.655
R29254 vdd.n13104 vdd.n9283 133.655
R29255 vdd.n13102 vdd.n13101 133.655
R29256 vdd.n13098 vdd.n13097 133.655
R29257 vdd.n13094 vdd.n13093 133.655
R29258 vdd.n13090 vdd.n13089 133.655
R29259 vdd.n13112 vdd.n9275 133.655
R29260 vdd.n14596 vdd.n14574 133.655
R29261 vdd.n14594 vdd.n14593 133.655
R29262 vdd.n14590 vdd.n14589 133.655
R29263 vdd.n14586 vdd.n14585 133.655
R29264 vdd.n14582 vdd.n14581 133.655
R29265 vdd.n14578 vdd.n14577 133.655
R29266 vdd.n14703 vdd.n8114 133.655
R29267 vdd.n14877 vdd.n8029 133.655
R29268 vdd.n14946 vdd.n7988 133.655
R29269 vdd.n14657 vdd.n8142 133.655
R29270 vdd.n14661 vdd.n8142 133.655
R29271 vdd.n14661 vdd.n8123 133.655
R29272 vdd.n14696 vdd.n8123 133.655
R29273 vdd.n14696 vdd.n8120 133.655
R29274 vdd.n14701 vdd.n8120 133.655
R29275 vdd.n14701 vdd.n8121 133.655
R29276 vdd.n8121 vdd.n8103 133.655
R29277 vdd.n14742 vdd.n8103 133.655
R29278 vdd.n14742 vdd.n8101 133.655
R29279 vdd.n14747 vdd.n8101 133.655
R29280 vdd.n14747 vdd.n8081 133.655
R29281 vdd.n14774 vdd.n8081 133.655
R29282 vdd.n14775 vdd.n14774 133.655
R29283 vdd.n14775 vdd.n8074 133.655
R29284 vdd.n14779 vdd.n8074 133.655
R29285 vdd.n14779 vdd.n8053 133.655
R29286 vdd.n14829 vdd.n8053 133.655
R29287 vdd.n14829 vdd.n8051 133.655
R29288 vdd.n14833 vdd.n8051 133.655
R29289 vdd.n14833 vdd.n8033 133.655
R29290 vdd.n14870 vdd.n8033 133.655
R29291 vdd.n14870 vdd.n8031 133.655
R29292 vdd.n14874 vdd.n8031 133.655
R29293 vdd.n14874 vdd.n8019 133.655
R29294 vdd.n14907 vdd.n8019 133.655
R29295 vdd.n14907 vdd.n8017 133.655
R29296 vdd.n14912 vdd.n8017 133.655
R29297 vdd.n14912 vdd.n8010 133.655
R29298 vdd.n8010 vdd.n8000 133.655
R29299 vdd.n14943 vdd.n8000 133.655
R29300 vdd.n14638 vdd.n8167 133.655
R29301 vdd.n14636 vdd.n14635 133.655
R29302 vdd.n14632 vdd.n14631 133.655
R29303 vdd.n14628 vdd.n14627 133.655
R29304 vdd.n14624 vdd.n14623 133.655
R29305 vdd.n14620 vdd.n14619 133.655
R29306 vdd.n11629 vdd.n9243 133.655
R29307 vdd.n13146 vdd.n9243 133.655
R29308 vdd.n13146 vdd.n9240 133.655
R29309 vdd.n13151 vdd.n9240 133.655
R29310 vdd.n13151 vdd.n9241 133.655
R29311 vdd.n9241 vdd.n9189 133.655
R29312 vdd.n13230 vdd.n9189 133.655
R29313 vdd.n13230 vdd.n9186 133.655
R29314 vdd.n13236 vdd.n9186 133.655
R29315 vdd.n13236 vdd.n9187 133.655
R29316 vdd.n9187 vdd.n9159 133.655
R29317 vdd.n9159 vdd.n9129 133.655
R29318 vdd.n13317 vdd.n9129 133.655
R29319 vdd.n13317 vdd.n9126 133.655
R29320 vdd.n13326 vdd.n9126 133.655
R29321 vdd.n13326 vdd.n9127 133.655
R29322 vdd.n13322 vdd.n9127 133.655
R29323 vdd.n13322 vdd.n13321 133.655
R29324 vdd.n13321 vdd.n9019 133.655
R29325 vdd.n13439 vdd.n9019 133.655
R29326 vdd.n13439 vdd.n9016 133.655
R29327 vdd.n13444 vdd.n9016 133.655
R29328 vdd.n13444 vdd.n9017 133.655
R29329 vdd.n9017 vdd.n8968 133.655
R29330 vdd.n13522 vdd.n8968 133.655
R29331 vdd.n13522 vdd.n8965 133.655
R29332 vdd.n13528 vdd.n8965 133.655
R29333 vdd.n13528 vdd.n8966 133.655
R29334 vdd.n8966 vdd.n8937 133.655
R29335 vdd.n8937 vdd.n8908 133.655
R29336 vdd.n13609 vdd.n8908 133.655
R29337 vdd.n13609 vdd.n8905 133.655
R29338 vdd.n13618 vdd.n8905 133.655
R29339 vdd.n13618 vdd.n8906 133.655
R29340 vdd.n13614 vdd.n8906 133.655
R29341 vdd.n13614 vdd.n13613 133.655
R29342 vdd.n13613 vdd.n8799 133.655
R29343 vdd.n13731 vdd.n8799 133.655
R29344 vdd.n13731 vdd.n8797 133.655
R29345 vdd.n13735 vdd.n8797 133.655
R29346 vdd.n13735 vdd.n8752 133.655
R29347 vdd.n13804 vdd.n8752 133.655
R29348 vdd.n13804 vdd.n8750 133.655
R29349 vdd.n13808 vdd.n8750 133.655
R29350 vdd.n13808 vdd.n8711 133.655
R29351 vdd.n13865 vdd.n8711 133.655
R29352 vdd.n13865 vdd.n8709 133.655
R29353 vdd.n13869 vdd.n8709 133.655
R29354 vdd.n13869 vdd.n8645 133.655
R29355 vdd.n13928 vdd.n8645 133.655
R29356 vdd.n13928 vdd.n8642 133.655
R29357 vdd.n13933 vdd.n8642 133.655
R29358 vdd.n13933 vdd.n8643 133.655
R29359 vdd.n8643 vdd.n8592 133.655
R29360 vdd.n14005 vdd.n8592 133.655
R29361 vdd.n14005 vdd.n8589 133.655
R29362 vdd.n14010 vdd.n8589 133.655
R29363 vdd.n14010 vdd.n8590 133.655
R29364 vdd.n8590 vdd.n8539 133.655
R29365 vdd.n14091 vdd.n8539 133.655
R29366 vdd.n14091 vdd.n8537 133.655
R29367 vdd.n14095 vdd.n8537 133.655
R29368 vdd.n14095 vdd.n8488 133.655
R29369 vdd.n14154 vdd.n8488 133.655
R29370 vdd.n14154 vdd.n8486 133.655
R29371 vdd.n14158 vdd.n8486 133.655
R29372 vdd.n14158 vdd.n8424 133.655
R29373 vdd.n14218 vdd.n8424 133.655
R29374 vdd.n14218 vdd.n8421 133.655
R29375 vdd.n14223 vdd.n8421 133.655
R29376 vdd.n14223 vdd.n8422 133.655
R29377 vdd.n8422 vdd.n8370 133.655
R29378 vdd.n14296 vdd.n8370 133.655
R29379 vdd.n14296 vdd.n8368 133.655
R29380 vdd.n14300 vdd.n8368 133.655
R29381 vdd.n14300 vdd.n8316 133.655
R29382 vdd.n14373 vdd.n8316 133.655
R29383 vdd.n14373 vdd.n8313 133.655
R29384 vdd.n14380 vdd.n8313 133.655
R29385 vdd.n14380 vdd.n8314 133.655
R29386 vdd.n14376 vdd.n8314 133.655
R29387 vdd.n14376 vdd.n8238 133.655
R29388 vdd.n14462 vdd.n8238 133.655
R29389 vdd.n14462 vdd.n8235 133.655
R29390 vdd.n14467 vdd.n8235 133.655
R29391 vdd.n14467 vdd.n8236 133.655
R29392 vdd.n8236 vdd.n8186 133.655
R29393 vdd.n14560 vdd.n8186 133.655
R29394 vdd.n14560 vdd.n8184 133.655
R29395 vdd.n14565 vdd.n8184 133.655
R29396 vdd.n14565 vdd.n8171 133.655
R29397 vdd.n14615 vdd.n8171 133.655
R29398 vdd.n11652 vdd.n11574 133.655
R29399 vdd.n11650 vdd.n11649 133.655
R29400 vdd.n11646 vdd.n11645 133.655
R29401 vdd.n11642 vdd.n11641 133.655
R29402 vdd.n11638 vdd.n11637 133.655
R29403 vdd.n11634 vdd.n11633 133.655
R29404 vdd.n20539 vdd.n20511 117.283
R29405 vdd.n21740 vdd.n21739 114.647
R29406 vdd.n24871 vdd.n24870 112.187
R29407 vdd.n24874 vdd.n24873 112.187
R29408 vdd.n24858 vdd.n24857 112.187
R29409 vdd.n24852 vdd.n24851 112.187
R29410 vdd.t188 vdd.n11730 111.965
R29411 vdd.n11834 vdd.n11813 111.965
R29412 vdd.n21925 vdd.n21904 111.965
R29413 vdd.t296 vdd.n9297 111.65
R29414 vdd.n24568 vdd.t199 110.607
R29415 vdd.n24992 vdd.t205 110.602
R29416 vdd.n24568 vdd.t238 110.599
R29417 vdd.n24992 vdd.t235 110.586
R29418 vdd.n13131 vdd.n9265 104.172
R29419 vdd.n13127 vdd.n9214 104.172
R29420 vdd.n13189 vdd.n9215 104.172
R29421 vdd.n13185 vdd.n13178 104.172
R29422 vdd.n13206 vdd.n9203 104.172
R29423 vdd.n13247 vdd.n9164 104.172
R29424 vdd.n13275 vdd.n9160 104.172
R29425 vdd.n13288 vdd.n9143 104.172
R29426 vdd.n13294 vdd.n9144 104.172
R29427 vdd.n13337 vdd.n9095 104.172
R29428 vdd.n9124 vdd.n9096 104.172
R29429 vdd.n13367 vdd.n9069 104.172
R29430 vdd.n13374 vdd.n9063 104.172
R29431 vdd.n13374 vdd.n9047 104.172
R29432 vdd.n9054 vdd.n9048 104.172
R29433 vdd.n13392 vdd.n9041 104.172
R29434 vdd.n13425 vdd.n9034 104.172
R29435 vdd.n13421 vdd.n8994 104.172
R29436 vdd.n13483 vdd.n8995 104.172
R29437 vdd.n13479 vdd.n13473 104.172
R29438 vdd.n13500 vdd.n8982 104.172
R29439 vdd.n13539 vdd.n8943 104.172
R29440 vdd.n13567 vdd.n8938 104.172
R29441 vdd.n13580 vdd.n8922 104.172
R29442 vdd.n13586 vdd.n8923 104.172
R29443 vdd.n13629 vdd.n8875 104.172
R29444 vdd.n8903 vdd.n8876 104.172
R29445 vdd.n13659 vdd.n8849 104.172
R29446 vdd.n13666 vdd.n8843 104.172
R29447 vdd.n13666 vdd.n8826 104.172
R29448 vdd.n8834 vdd.n8827 104.172
R29449 vdd.n13684 vdd.n8820 104.172
R29450 vdd.n13717 vdd.n8813 104.172
R29451 vdd.n13713 vdd.n8777 104.172
R29452 vdd.n13763 vdd.n8778 104.172
R29453 vdd.n13759 vdd.n8772 104.172
R29454 vdd.n13790 vdd.n8767 104.172
R29455 vdd.n13824 vdd.n8727 104.172
R29456 vdd.n13855 vdd.n8720 104.172
R29457 vdd.n13848 vdd.n8683 104.172
R29458 vdd.n13890 vdd.n8684 104.172
R29459 vdd.n13907 vdd.n8676 104.172
R29460 vdd.n13914 vdd.n8658 104.172
R29461 vdd.n8665 vdd.n8622 104.172
R29462 vdd.n13962 vdd.n8623 104.172
R29463 vdd.n13962 vdd.n8628 104.172
R29464 vdd.n13979 vdd.n13977 104.172
R29465 vdd.n13991 vdd.n8602 104.172
R29466 vdd.n13987 vdd.n8566 104.172
R29467 vdd.n14053 vdd.n8567 104.172
R29468 vdd.n14049 vdd.n14039 104.172
R29469 vdd.n14071 vdd.n14070 104.172
R29470 vdd.n14077 vdd.n8513 104.172
R29471 vdd.n14129 vdd.n14128 104.172
R29472 vdd.n14144 vdd.n8499 104.172
R29473 vdd.n14137 vdd.n8459 104.172
R29474 vdd.n14179 vdd.n8460 104.172
R29475 vdd.n14197 vdd.n8452 104.172
R29476 vdd.n14204 vdd.n8437 104.172
R29477 vdd.n8442 vdd.n8400 104.172
R29478 vdd.n14252 vdd.n8401 104.172
R29479 vdd.n14252 vdd.n8406 104.172
R29480 vdd.n14269 vdd.n14267 104.172
R29481 vdd.n14282 vdd.n8380 104.172
R29482 vdd.n14278 vdd.n8348 104.172
R29483 vdd.n14328 vdd.n8349 104.172
R29484 vdd.n14324 vdd.n8341 104.172
R29485 vdd.n14359 vdd.n8334 104.172
R29486 vdd.n14355 vdd.n8302 104.172
R29487 vdd.n14421 vdd.n8276 104.172
R29488 vdd.n14460 vdd.n8242 104.172
R29489 vdd.n14453 vdd.n8251 104.172
R29490 vdd.n8260 vdd.n8253 104.172
R29491 vdd.n14489 vdd.n8217 104.172
R29492 vdd.n14647 vdd.n8148 104.172
R29493 vdd.n8159 vdd.n8139 104.172
R29494 vdd.n14671 vdd.n8135 104.172
R29495 vdd.n14675 vdd.n8126 104.172
R29496 vdd.n14686 vdd.n8127 104.172
R29497 vdd.n14703 vdd.n8118 104.172
R29498 vdd.n14711 vdd.n8114 104.172
R29499 vdd.n14715 vdd.n8106 104.172
R29500 vdd.n14732 vdd.n8107 104.172
R29501 vdd.n14728 vdd.n8099 104.172
R29502 vdd.n14757 vdd.n8095 104.172
R29503 vdd.n14761 vdd.n8084 104.172
R29504 vdd.n8088 vdd.n8085 104.172
R29505 vdd.n14790 vdd.n8071 104.172
R29506 vdd.n14799 vdd.n8065 104.172
R29507 vdd.n14803 vdd.n8056 104.172
R29508 vdd.n14819 vdd.n8057 104.172
R29509 vdd.n14815 vdd.n8049 104.172
R29510 vdd.n14843 vdd.n8045 104.172
R29511 vdd.n14847 vdd.n8036 104.172
R29512 vdd.n14860 vdd.n8037 104.172
R29513 vdd.n14856 vdd.n8029 104.172
R29514 vdd.n14877 vdd.n8022 104.172
R29515 vdd.n14897 vdd.n8023 104.172
R29516 vdd.n14893 vdd.n14886 104.172
R29517 vdd.n14915 vdd.n8011 104.172
R29518 vdd.n14933 vdd.n8007 104.172
R29519 vdd.n14929 vdd.n8002 104.172
R29520 vdd.n9262 vdd.n9247 104.172
R29521 vdd.n13154 vdd.n9238 104.172
R29522 vdd.n13163 vdd.n13160 104.172
R29523 vdd.n13169 vdd.n9223 104.172
R29524 vdd.n13176 vdd.n9192 104.172
R29525 vdd.n13220 vdd.n9193 104.172
R29526 vdd.n13239 vdd.n9184 104.172
R29527 vdd.n13244 vdd.n9181 104.172
R29528 vdd.n9181 vdd.n9156 104.172
R29529 vdd.n13285 vdd.n9152 104.172
R29530 vdd.n13305 vdd.n9133 104.172
R29531 vdd.n13334 vdd.n9106 104.172
R29532 vdd.n13330 vdd.n13329 104.172
R29533 vdd.n13364 vdd.n9072 104.172
R29534 vdd.n13360 vdd.n9088 104.172
R29535 vdd.n13379 vdd.n9061 104.172
R29536 vdd.n13429 vdd.n9023 104.172
R29537 vdd.n13447 vdd.n9015 104.172
R29538 vdd.n13456 vdd.n13454 104.172
R29539 vdd.n13471 vdd.n9003 104.172
R29540 vdd.n13464 vdd.n8970 104.172
R29541 vdd.n13512 vdd.n8971 104.172
R29542 vdd.n13531 vdd.n8963 104.172
R29543 vdd.n13536 vdd.n8960 104.172
R29544 vdd.n8960 vdd.n8935 104.172
R29545 vdd.n13577 vdd.n8931 104.172
R29546 vdd.n13597 vdd.n8911 104.172
R29547 vdd.n13626 vdd.n8885 104.172
R29548 vdd.n13622 vdd.n13621 104.172
R29549 vdd.n13656 vdd.n8852 104.172
R29550 vdd.n13652 vdd.n8868 104.172
R29551 vdd.n13671 vdd.n8841 104.172
R29552 vdd.n13721 vdd.n8803 104.172
R29553 vdd.n13738 vdd.n8795 104.172
R29554 vdd.n13747 vdd.n13744 104.172
R29555 vdd.n13754 vdd.n8755 104.172
R29556 vdd.n13794 vdd.n8756 104.172
R29557 vdd.n13811 vdd.n8745 104.172
R29558 vdd.n8747 vdd.n8740 104.172
R29559 vdd.n13863 vdd.n8713 104.172
R29560 vdd.n13863 vdd.n8714 104.172
R29561 vdd.n13872 vdd.n8706 104.172
R29562 vdd.n13880 vdd.n13878 104.172
R29563 vdd.n13887 vdd.n8647 104.172
R29564 vdd.n13918 vdd.n8648 104.172
R29565 vdd.n13936 vdd.n8640 104.172
R29566 vdd.n13944 vdd.n8620 104.172
R29567 vdd.n13959 vdd.n8633 104.172
R29568 vdd.n14013 vdd.n8587 104.172
R29569 vdd.n14022 vdd.n14020 104.172
R29570 vdd.n14037 vdd.n8575 104.172
R29571 vdd.n14030 vdd.n8542 104.172
R29572 vdd.n14081 vdd.n8543 104.172
R29573 vdd.n14098 vdd.n8533 104.172
R29574 vdd.n14106 vdd.n8526 104.172
R29575 vdd.n14152 vdd.n8491 104.172
R29576 vdd.n14152 vdd.n8492 104.172
R29577 vdd.n14161 vdd.n8483 104.172
R29578 vdd.n14169 vdd.n14167 104.172
R29579 vdd.n14176 vdd.n8427 104.172
R29580 vdd.n14208 vdd.n8428 104.172
R29581 vdd.n14226 vdd.n8418 104.172
R29582 vdd.n14234 vdd.n8398 104.172
R29583 vdd.n14249 vdd.n8411 104.172
R29584 vdd.n14303 vdd.n8367 104.172
R29585 vdd.n14311 vdd.n14309 104.172
R29586 vdd.n14318 vdd.n8319 104.172
R29587 vdd.n14363 vdd.n8320 104.172
R29588 vdd.n8332 vdd.n8311 104.172
R29589 vdd.n14393 vdd.n8305 104.172
R29590 vdd.n14410 vdd.n8295 104.172
R29591 vdd.n14418 vdd.n8288 104.172
R29592 vdd.n14418 vdd.n8289 104.172
R29593 vdd.n14441 vdd.n8268 104.172
R29594 vdd.n14450 vdd.n8231 104.172
R29595 vdd.n14486 vdd.n8225 104.172
R29596 vdd.n14482 vdd.n14481 104.172
R29597 vdd.n14532 vdd.n8189 104.172
R29598 vdd.n14550 vdd.n8190 104.172
R29599 vdd.n14546 vdd.n14540 104.172
R29600 vdd.n13256 vdd.n9171 102.206
R29601 vdd.n13256 vdd.n9172 102.206
R29602 vdd.n13547 vdd.n8951 102.206
R29603 vdd.n13547 vdd.n8952 102.206
R29604 vdd.n13832 vdd.n8732 102.206
R29605 vdd.n13832 vdd.n8733 102.206
R29606 vdd.n8523 vdd.n8514 102.206
R29607 vdd.n14109 vdd.n8523 102.206
R29608 vdd.n14405 vdd.n8298 102.206
R29609 vdd.n14405 vdd.n8275 102.206
R29610 vdd.n11581 vdd.n11578 102.206
R29611 vdd.n11581 vdd.n9246 102.206
R29612 vdd.n13388 vdd.n9057 102.206
R29613 vdd.n13388 vdd.n9022 102.206
R29614 vdd.n13680 vdd.n8837 102.206
R29615 vdd.n13680 vdd.n8802 102.206
R29616 vdd.n14003 vdd.n8595 102.206
R29617 vdd.n14003 vdd.n8596 102.206
R29618 vdd.n14294 vdd.n8373 102.206
R29619 vdd.n14294 vdd.n8374 102.206
R29620 vdd.n14604 vdd.n8182 102.206
R29621 vdd.n8182 vdd.n8175 102.206
R29622 vdd.n10520 vdd.n10517 97.78
R29623 vdd.n24834 vdd.t138 97.742
R29624 vdd.t204 vdd.n24846 97.742
R29625 vdd.n35841 vdd.n35840 92.5
R29626 vdd.n35834 vdd.n35833 92.5
R29627 vdd.n35831 vdd.n35830 92.5
R29628 vdd.n35829 vdd.n35828 92.5
R29629 vdd.n35826 vdd.n35825 92.5
R29630 vdd.n35824 vdd.n35823 92.5
R29631 vdd.n35821 vdd.n35820 92.5
R29632 vdd.n35819 vdd.n35818 92.5
R29633 vdd.n35816 vdd.n35815 92.5
R29634 vdd.n35814 vdd.n35813 92.5
R29635 vdd.n35811 vdd.n35810 92.5
R29636 vdd.n35809 vdd.n35808 92.5
R29637 vdd.n35806 vdd.n35805 92.5
R29638 vdd.n35804 vdd.n35803 92.5
R29639 vdd.n35801 vdd.n35800 92.5
R29640 vdd.n35799 vdd.n35798 92.5
R29641 vdd.n35796 vdd.n35795 92.5
R29642 vdd.n35794 vdd.n35793 92.5
R29643 vdd.n35791 vdd.n35790 92.5
R29644 vdd.n35789 vdd.n35788 92.5
R29645 vdd.n35786 vdd.n35785 92.5
R29646 vdd.n35784 vdd.n35783 92.5
R29647 vdd.n35781 vdd.n35780 92.5
R29648 vdd.n35779 vdd.n35778 92.5
R29649 vdd.n35776 vdd.n35775 92.5
R29650 vdd.n35774 vdd.n35773 92.5
R29651 vdd.n35771 vdd.n35770 92.5
R29652 vdd.n35769 vdd.n35768 92.5
R29653 vdd.n35766 vdd.n35765 92.5
R29654 vdd.n35764 vdd.n35763 92.5
R29655 vdd.n35761 vdd.n35760 92.5
R29656 vdd.n35759 vdd.n35758 92.5
R29657 vdd.n35756 vdd.n35755 92.5
R29658 vdd.n35754 vdd.n35753 92.5
R29659 vdd.n35751 vdd.n35750 92.5
R29660 vdd.n35749 vdd.n35748 92.5
R29661 vdd.n35746 vdd.n35745 92.5
R29662 vdd.n35744 vdd.n35743 92.5
R29663 vdd.n35741 vdd.n35740 92.5
R29664 vdd.n35739 vdd.n35738 92.5
R29665 vdd.n35736 vdd.n35735 92.5
R29666 vdd.n35734 vdd.n35733 92.5
R29667 vdd.n35731 vdd.n35730 92.5
R29668 vdd.n35729 vdd.n35728 92.5
R29669 vdd.n35726 vdd.n35725 92.5
R29670 vdd.n35724 vdd.n35723 92.5
R29671 vdd.n29682 vdd.n29681 92.5
R29672 vdd.n28155 vdd.n28154 92.5
R29673 vdd.n28341 vdd.n28340 92.5
R29674 vdd.n37899 vdd.n37898 92.5
R29675 vdd.n32896 vdd.n32895 92.5
R29676 vdd.n33227 vdd.n33226 92.5
R29677 vdd.n36613 vdd.n36612 92.5
R29678 vdd.n36151 vdd.n36150 92.5
R29679 vdd.n35920 vdd.n35919 92.5
R29680 vdd.n36382 vdd.n36381 92.5
R29681 vdd.n36844 vdd.n36843 92.5
R29682 vdd.n37241 vdd.n37240 92.5
R29683 vdd.n38116 vdd.n38115 92.5
R29684 vdd.n37668 vdd.n37667 92.5
R29685 vdd.n28572 vdd.n28571 92.5
R29686 vdd.n27758 vdd.n27757 92.5
R29687 vdd.n30573 vdd.n30572 92.5
R29688 vdd.n30361 vdd.n30360 92.5
R29689 vdd.n30365 vdd.n30364 92.5
R29690 vdd.n30371 vdd.n30370 92.5
R29691 vdd.n30369 vdd.n30368 92.5
R29692 vdd.n30374 vdd.n30373 92.5
R29693 vdd.n30377 vdd.n30376 92.5
R29694 vdd.n30380 vdd.n30379 92.5
R29695 vdd.n30383 vdd.n30382 92.5
R29696 vdd.n30386 vdd.n30385 92.5
R29697 vdd.n30390 vdd.n30389 92.5
R29698 vdd.n30395 vdd.n30394 92.5
R29699 vdd.n30393 vdd.n30392 92.5
R29700 vdd.n30399 vdd.n30398 92.5
R29701 vdd.n30404 vdd.n30403 92.5
R29702 vdd.n30402 vdd.n30401 92.5
R29703 vdd.n30410 vdd.n30409 92.5
R29704 vdd.n30408 vdd.n30407 92.5
R29705 vdd.n30414 vdd.n30413 92.5
R29706 vdd.n30419 vdd.n30418 92.5
R29707 vdd.n30417 vdd.n30416 92.5
R29708 vdd.n30422 vdd.n30421 92.5
R29709 vdd.n30428 vdd.n30427 92.5
R29710 vdd.n30426 vdd.n30425 92.5
R29711 vdd.n30431 vdd.n30430 92.5
R29712 vdd.n30437 vdd.n30436 92.5
R29713 vdd.n30435 vdd.n30434 92.5
R29714 vdd.n30441 vdd.n30440 92.5
R29715 vdd.n30446 vdd.n30445 92.5
R29716 vdd.n30444 vdd.n30443 92.5
R29717 vdd.n30449 vdd.n30448 92.5
R29718 vdd.n30455 vdd.n30454 92.5
R29719 vdd.n30453 vdd.n30452 92.5
R29720 vdd.n30461 vdd.n30460 92.5
R29721 vdd.n30459 vdd.n30458 92.5
R29722 vdd.n30464 vdd.n30463 92.5
R29723 vdd.n30468 vdd.n30467 92.5
R29724 vdd.n30473 vdd.n30472 92.5
R29725 vdd.n30471 vdd.n30470 92.5
R29726 vdd.n30476 vdd.n30475 92.5
R29727 vdd.n30479 vdd.n30478 92.5
R29728 vdd.n30482 vdd.n30481 92.5
R29729 vdd.n30500 vdd.n30347 92.5
R29730 vdd.n31020 vdd.n31019 92.5
R29731 vdd.n32238 vdd.n32237 92.5
R29732 vdd.n2022 vdd.n2021 92.5
R29733 vdd.n2800 vdd.n2799 92.5
R29734 vdd.n2981 vdd.n2980 92.5
R29735 vdd.n3162 vdd.n3161 92.5
R29736 vdd.n3343 vdd.n3342 92.5
R29737 vdd.n3524 vdd.n3523 92.5
R29738 vdd.n2681 vdd.n2680 92.5
R29739 vdd.n2002 vdd.n2001 92.5
R29740 vdd.n1733 vdd.n1732 92.5
R29741 vdd.n1562 vdd.n1561 92.5
R29742 vdd.n1381 vdd.n1380 92.5
R29743 vdd.n26847 vdd.n26846 92.5
R29744 vdd.n27028 vdd.n27027 92.5
R29745 vdd.n26747 vdd.n26746 92.5
R29746 vdd.n31688 vdd.n31687 92.5
R29747 vdd.n14944 vdd.n14943 92.5
R29748 vdd.n14943 vdd.n14942 92.5
R29749 vdd.n14931 vdd.n8000 92.5
R29750 vdd.n14926 vdd.n8010 92.5
R29751 vdd.n14913 vdd.n14912 92.5
R29752 vdd.n14895 vdd.n8017 92.5
R29753 vdd.n14907 vdd.n14906 92.5
R29754 vdd.n14858 vdd.n8031 92.5
R29755 vdd.n14870 vdd.n14869 92.5
R29756 vdd.n14845 vdd.n8033 92.5
R29757 vdd.n14834 vdd.n14833 92.5
R29758 vdd.n14817 vdd.n8051 92.5
R29759 vdd.n14829 vdd.n14828 92.5
R29760 vdd.n14801 vdd.n8053 92.5
R29761 vdd.n14780 vdd.n14779 92.5
R29762 vdd.n14787 vdd.n8074 92.5
R29763 vdd.n14775 vdd.n8072 92.5
R29764 vdd.n14774 vdd.n14773 92.5
R29765 vdd.n14759 vdd.n8081 92.5
R29766 vdd.n14748 vdd.n14747 92.5
R29767 vdd.n14730 vdd.n8101 92.5
R29768 vdd.n14742 vdd.n14741 92.5
R29769 vdd.n14713 vdd.n8103 92.5
R29770 vdd.n14684 vdd.n8120 92.5
R29771 vdd.n14696 vdd.n14695 92.5
R29772 vdd.n14673 vdd.n8123 92.5
R29773 vdd.n14947 vdd.n14946 92.5
R29774 vdd.n14949 vdd.n14948 92.5
R29775 vdd.n14951 vdd.n14950 92.5
R29776 vdd.n14953 vdd.n14952 92.5
R29777 vdd.n14955 vdd.n14954 92.5
R29778 vdd.n14957 vdd.n14956 92.5
R29779 vdd.n14959 vdd.n14958 92.5
R29780 vdd.n14961 vdd.n14960 92.5
R29781 vdd.n14963 vdd.n14962 92.5
R29782 vdd.n14965 vdd.n14964 92.5
R29783 vdd.n14967 vdd.n14966 92.5
R29784 vdd.n7986 vdd.n7984 92.5
R29785 vdd.n14972 vdd.n14971 92.5
R29786 vdd.n8029 vdd.n8028 92.5
R29787 vdd.n14875 vdd.n8029 92.5
R29788 vdd.n14705 vdd.n8114 92.5
R29789 vdd.n8114 vdd.n8113 92.5
R29790 vdd.n14704 vdd.n14703 92.5
R29791 vdd.n14703 vdd.n14702 92.5
R29792 vdd.n14878 vdd.n14877 92.5
R29793 vdd.n14877 vdd.n14876 92.5
R29794 vdd.n14945 vdd.n7988 92.5
R29795 vdd.n14969 vdd.n7988 92.5
R29796 vdd.n8000 vdd.n7999 92.5
R29797 vdd.n14910 vdd.n8010 92.5
R29798 vdd.n14912 vdd.n14911 92.5
R29799 vdd.n14909 vdd.n8017 92.5
R29800 vdd.n14908 vdd.n14907 92.5
R29801 vdd.n8019 vdd.n8018 92.5
R29802 vdd.n14876 vdd.n8019 92.5
R29803 vdd.n14874 vdd.n14873 92.5
R29804 vdd.n14875 vdd.n14874 92.5
R29805 vdd.n14872 vdd.n8031 92.5
R29806 vdd.n14871 vdd.n14870 92.5
R29807 vdd.n8033 vdd.n8032 92.5
R29808 vdd.n14833 vdd.n14832 92.5
R29809 vdd.n14831 vdd.n8051 92.5
R29810 vdd.n14830 vdd.n14829 92.5
R29811 vdd.n8053 vdd.n8052 92.5
R29812 vdd.n14779 vdd.n14778 92.5
R29813 vdd.n14777 vdd.n8074 92.5
R29814 vdd.n14776 vdd.n14775 92.5
R29815 vdd.n14774 vdd.n8080 92.5
R29816 vdd.n14745 vdd.n8081 92.5
R29817 vdd.n14747 vdd.n14746 92.5
R29818 vdd.n14744 vdd.n8101 92.5
R29819 vdd.n14743 vdd.n14742 92.5
R29820 vdd.n8103 vdd.n8102 92.5
R29821 vdd.n14699 vdd.n8121 92.5
R29822 vdd.n8121 vdd.n8113 92.5
R29823 vdd.n14701 vdd.n14700 92.5
R29824 vdd.n14702 vdd.n14701 92.5
R29825 vdd.n14698 vdd.n8120 92.5
R29826 vdd.n14697 vdd.n14696 92.5
R29827 vdd.n8123 vdd.n8122 92.5
R29828 vdd.n14662 vdd.n14661 92.5
R29829 vdd.n14645 vdd.n8142 92.5
R29830 vdd.n14661 vdd.n14660 92.5
R29831 vdd.n14659 vdd.n8142 92.5
R29832 vdd.n14598 vdd.n14574 92.5
R29833 vdd.n14597 vdd.n14596 92.5
R29834 vdd.n14595 vdd.n14594 92.5
R29835 vdd.n14593 vdd.n14592 92.5
R29836 vdd.n14591 vdd.n14590 92.5
R29837 vdd.n14589 vdd.n14588 92.5
R29838 vdd.n14587 vdd.n14586 92.5
R29839 vdd.n14585 vdd.n14584 92.5
R29840 vdd.n14583 vdd.n14582 92.5
R29841 vdd.n14581 vdd.n14580 92.5
R29842 vdd.n14579 vdd.n14578 92.5
R29843 vdd.n14577 vdd.n14576 92.5
R29844 vdd.n8144 vdd.n8143 92.5
R29845 vdd.n14657 vdd.n14656 92.5
R29846 vdd.n14658 vdd.n14657 92.5
R29847 vdd.n14600 vdd.n14599 92.5
R29848 vdd.n14505 vdd.n14504 92.5
R29849 vdd.n14507 vdd.n14506 92.5
R29850 vdd.n14509 vdd.n14508 92.5
R29851 vdd.n14511 vdd.n14510 92.5
R29852 vdd.n14513 vdd.n14512 92.5
R29853 vdd.n14515 vdd.n14514 92.5
R29854 vdd.n14517 vdd.n14516 92.5
R29855 vdd.n14519 vdd.n14518 92.5
R29856 vdd.n14521 vdd.n14520 92.5
R29857 vdd.n14523 vdd.n14522 92.5
R29858 vdd.n14525 vdd.n14524 92.5
R29859 vdd.n14526 vdd.n8210 92.5
R29860 vdd.n14528 vdd.n14527 92.5
R29861 vdd.n14503 vdd.n8198 92.5
R29862 vdd.n14530 vdd.n8198 92.5
R29863 vdd.n14502 vdd.n14501 92.5
R29864 vdd.n14501 vdd.n14500 92.5
R29865 vdd.n8214 vdd.n8213 92.5
R29866 vdd.n8222 vdd.n8214 92.5
R29867 vdd.n14434 vdd.n8270 92.5
R29868 vdd.n8270 vdd.n8262 92.5
R29869 vdd.n14436 vdd.n14435 92.5
R29870 vdd.n14437 vdd.n14436 92.5
R29871 vdd.n14433 vdd.n8269 92.5
R29872 vdd.n8287 vdd.n8269 92.5
R29873 vdd.n14432 vdd.n14431 92.5
R29874 vdd.n14431 vdd.n14430 92.5
R29875 vdd.n8272 vdd.n8271 92.5
R29876 vdd.n14406 vdd.n8272 92.5
R29877 vdd.n14341 vdd.n8304 92.5
R29878 vdd.n14396 vdd.n8304 92.5
R29879 vdd.n14342 vdd.n8343 92.5
R29880 vdd.n8343 vdd.n8333 92.5
R29881 vdd.n14344 vdd.n14343 92.5
R29882 vdd.n14345 vdd.n14344 92.5
R29883 vdd.n14340 vdd.n8342 92.5
R29884 vdd.n14326 vdd.n8342 92.5
R29885 vdd.n14339 vdd.n14338 92.5
R29886 vdd.n14338 vdd.n14337 92.5
R29887 vdd.n8345 vdd.n8344 92.5
R29888 vdd.n8378 vdd.n8345 92.5
R29889 vdd.n14261 vdd.n8394 92.5
R29890 vdd.n8394 vdd.n8372 92.5
R29891 vdd.n14263 vdd.n14262 92.5
R29892 vdd.n14264 vdd.n14263 92.5
R29893 vdd.n14260 vdd.n8393 92.5
R29894 vdd.n14251 vdd.n8393 92.5
R29895 vdd.n14259 vdd.n14258 92.5
R29896 vdd.n14258 vdd.n14257 92.5
R29897 vdd.n8396 vdd.n8395 92.5
R29898 vdd.n8438 vdd.n8396 92.5
R29899 vdd.n14193 vdd.n14192 92.5
R29900 vdd.n14195 vdd.n14193 92.5
R29901 vdd.n14191 vdd.n8454 92.5
R29902 vdd.n8472 vdd.n8454 92.5
R29903 vdd.n14190 vdd.n14189 92.5
R29904 vdd.n14189 vdd.n14188 92.5
R29905 vdd.n8456 vdd.n8455 92.5
R29906 vdd.n8500 vdd.n8456 92.5
R29907 vdd.n14122 vdd.n8509 92.5
R29908 vdd.n8509 vdd.n8490 92.5
R29909 vdd.n14124 vdd.n14123 92.5
R29910 vdd.n14125 vdd.n14124 92.5
R29911 vdd.n14121 vdd.n8508 92.5
R29912 vdd.n8536 vdd.n8508 92.5
R29913 vdd.n14120 vdd.n14119 92.5
R29914 vdd.n14119 vdd.n14118 92.5
R29915 vdd.n8511 vdd.n8510 92.5
R29916 vdd.n8552 vdd.n8511 92.5
R29917 vdd.n14067 vdd.n14066 92.5
R29918 vdd.n14068 vdd.n14067 92.5
R29919 vdd.n14065 vdd.n8561 92.5
R29920 vdd.n14051 vdd.n8561 92.5
R29921 vdd.n14064 vdd.n14063 92.5
R29922 vdd.n14063 vdd.n14062 92.5
R29923 vdd.n8563 vdd.n8562 92.5
R29924 vdd.n8600 vdd.n8563 92.5
R29925 vdd.n13971 vdd.n8616 92.5
R29926 vdd.n8616 vdd.n8594 92.5
R29927 vdd.n13973 vdd.n13972 92.5
R29928 vdd.n13974 vdd.n13973 92.5
R29929 vdd.n13970 vdd.n8615 92.5
R29930 vdd.n13961 vdd.n8615 92.5
R29931 vdd.n13969 vdd.n13968 92.5
R29932 vdd.n13968 vdd.n13967 92.5
R29933 vdd.n8618 vdd.n8617 92.5
R29934 vdd.n8663 vdd.n8618 92.5
R29935 vdd.n13904 vdd.n13903 92.5
R29936 vdd.n13905 vdd.n13904 92.5
R29937 vdd.n13902 vdd.n8678 92.5
R29938 vdd.n8695 vdd.n8678 92.5
R29939 vdd.n13901 vdd.n13900 92.5
R29940 vdd.n13900 vdd.n13899 92.5
R29941 vdd.n8680 vdd.n8679 92.5
R29942 vdd.n8721 vdd.n8680 92.5
R29943 vdd.n13838 vdd.n13837 92.5
R29944 vdd.n13840 vdd.n13838 92.5
R29945 vdd.n13836 vdd.n8728 92.5
R29946 vdd.n13821 vdd.n8728 92.5
R29947 vdd.n13835 vdd.n13834 92.5
R29948 vdd.n13834 vdd.n13833 92.5
R29949 vdd.n8730 vdd.n8729 92.5
R29950 vdd.n8766 vdd.n8730 92.5
R29951 vdd.n13777 vdd.n13776 92.5
R29952 vdd.n13778 vdd.n13777 92.5
R29953 vdd.n13775 vdd.n8773 92.5
R29954 vdd.n13761 vdd.n8773 92.5
R29955 vdd.n13774 vdd.n13773 92.5
R29956 vdd.n13773 vdd.n13772 92.5
R29957 vdd.n8775 vdd.n8774 92.5
R29958 vdd.n8812 vdd.n8775 92.5
R29959 vdd.n13702 vdd.n13701 92.5
R29960 vdd.n13704 vdd.n13702 92.5
R29961 vdd.n13700 vdd.n8821 92.5
R29962 vdd.n13682 vdd.n8821 92.5
R29963 vdd.n13699 vdd.n13698 92.5
R29964 vdd.n13698 vdd.n13697 92.5
R29965 vdd.n8823 vdd.n8822 92.5
R29966 vdd.n13667 vdd.n8823 92.5
R29967 vdd.n13645 vdd.n13644 92.5
R29968 vdd.n13651 vdd.n13645 92.5
R29969 vdd.n13643 vdd.n8870 92.5
R29970 vdd.n8870 vdd.n8850 92.5
R29971 vdd.n13642 vdd.n13641 92.5
R29972 vdd.n13641 vdd.n13640 92.5
R29973 vdd.n8872 vdd.n8871 92.5
R29974 vdd.n8882 vdd.n8872 92.5
R29975 vdd.n13552 vdd.n8919 92.5
R29976 vdd.n13595 vdd.n8919 92.5
R29977 vdd.n13553 vdd.n8946 92.5
R29978 vdd.n8946 vdd.n8929 92.5
R29979 vdd.n13555 vdd.n13554 92.5
R29980 vdd.n13558 vdd.n13555 92.5
R29981 vdd.n13551 vdd.n8945 92.5
R29982 vdd.n8957 vdd.n8945 92.5
R29983 vdd.n13550 vdd.n13549 92.5
R29984 vdd.n13549 vdd.n13548 92.5
R29985 vdd.n8948 vdd.n8947 92.5
R29986 vdd.n13509 vdd.n8948 92.5
R29987 vdd.n13497 vdd.n13496 92.5
R29988 vdd.n13498 vdd.n13497 92.5
R29989 vdd.n13495 vdd.n8989 92.5
R29990 vdd.n13481 vdd.n8989 92.5
R29991 vdd.n13494 vdd.n13493 92.5
R29992 vdd.n13493 vdd.n13492 92.5
R29993 vdd.n8991 vdd.n8990 92.5
R29994 vdd.n9033 vdd.n8991 92.5
R29995 vdd.n13409 vdd.n13408 92.5
R29996 vdd.n13410 vdd.n13409 92.5
R29997 vdd.n13407 vdd.n9042 92.5
R29998 vdd.n13390 vdd.n9042 92.5
R29999 vdd.n13406 vdd.n13405 92.5
R30000 vdd.n13405 vdd.n13404 92.5
R30001 vdd.n9044 vdd.n9043 92.5
R30002 vdd.n13375 vdd.n9044 92.5
R30003 vdd.n13353 vdd.n13352 92.5
R30004 vdd.n13359 vdd.n13353 92.5
R30005 vdd.n13351 vdd.n9090 92.5
R30006 vdd.n9090 vdd.n9070 92.5
R30007 vdd.n13350 vdd.n13349 92.5
R30008 vdd.n13349 vdd.n13348 92.5
R30009 vdd.n9092 vdd.n9091 92.5
R30010 vdd.n9103 vdd.n9092 92.5
R30011 vdd.n13261 vdd.n9141 92.5
R30012 vdd.n13303 vdd.n9141 92.5
R30013 vdd.n13262 vdd.n9167 92.5
R30014 vdd.n9167 vdd.n9150 92.5
R30015 vdd.n13264 vdd.n13263 92.5
R30016 vdd.n13266 vdd.n13264 92.5
R30017 vdd.n13260 vdd.n9166 92.5
R30018 vdd.n9178 vdd.n9166 92.5
R30019 vdd.n13259 vdd.n13258 92.5
R30020 vdd.n13258 vdd.n13257 92.5
R30021 vdd.n13256 vdd.n13255 92.5
R30022 vdd.n13257 vdd.n13256 92.5
R30023 vdd.n13547 vdd.n13546 92.5
R30024 vdd.n13548 vdd.n13547 92.5
R30025 vdd.n13832 vdd.n13831 92.5
R30026 vdd.n13833 vdd.n13832 92.5
R30027 vdd.n8523 vdd.n8522 92.5
R30028 vdd.n8536 vdd.n8523 92.5
R30029 vdd.n14405 vdd.n14404 92.5
R30030 vdd.n14406 vdd.n14405 92.5
R30031 vdd.n9169 vdd.n9168 92.5
R30032 vdd.n13216 vdd.n9169 92.5
R30033 vdd.n13203 vdd.n13202 92.5
R30034 vdd.n13204 vdd.n13203 92.5
R30035 vdd.n13201 vdd.n9209 92.5
R30036 vdd.n13187 vdd.n9209 92.5
R30037 vdd.n13200 vdd.n13199 92.5
R30038 vdd.n13199 vdd.n13198 92.5
R30039 vdd.n9211 vdd.n9210 92.5
R30040 vdd.n9264 vdd.n9211 92.5
R30041 vdd.n13106 vdd.n9283 92.5
R30042 vdd.n13105 vdd.n13104 92.5
R30043 vdd.n13103 vdd.n13102 92.5
R30044 vdd.n13101 vdd.n13100 92.5
R30045 vdd.n13099 vdd.n13098 92.5
R30046 vdd.n13097 vdd.n13096 92.5
R30047 vdd.n13095 vdd.n13094 92.5
R30048 vdd.n13093 vdd.n13092 92.5
R30049 vdd.n13091 vdd.n13090 92.5
R30050 vdd.n13089 vdd.n13088 92.5
R30051 vdd.n9275 vdd.n9274 92.5
R30052 vdd.n13113 vdd.n13112 92.5
R30053 vdd.n13114 vdd.n9273 92.5
R30054 vdd.n13116 vdd.n13115 92.5
R30055 vdd.n13118 vdd.n13116 92.5
R30056 vdd.n13108 vdd.n13107 92.5
R30057 vdd.n11582 vdd.n11581 92.5
R30058 vdd.n11581 vdd.n9277 92.5
R30059 vdd.n8182 vdd.n8181 92.5
R30060 vdd.n14567 vdd.n8182 92.5
R30061 vdd.n14294 vdd.n14293 92.5
R30062 vdd.n14295 vdd.n14294 92.5
R30063 vdd.n14003 vdd.n14002 92.5
R30064 vdd.n14004 vdd.n14003 92.5
R30065 vdd.n13680 vdd.n13679 92.5
R30066 vdd.n13681 vdd.n13680 92.5
R30067 vdd.n13388 vdd.n13387 92.5
R30068 vdd.n13389 vdd.n13388 92.5
R30069 vdd.n14640 vdd.n8167 92.5
R30070 vdd.n14639 vdd.n14638 92.5
R30071 vdd.n14637 vdd.n14636 92.5
R30072 vdd.n14635 vdd.n14634 92.5
R30073 vdd.n14633 vdd.n14632 92.5
R30074 vdd.n14631 vdd.n14630 92.5
R30075 vdd.n14629 vdd.n14628 92.5
R30076 vdd.n14627 vdd.n14626 92.5
R30077 vdd.n14625 vdd.n14624 92.5
R30078 vdd.n14623 vdd.n14622 92.5
R30079 vdd.n14621 vdd.n14620 92.5
R30080 vdd.n14619 vdd.n14618 92.5
R30081 vdd.n14617 vdd.n14616 92.5
R30082 vdd.n14642 vdd.n14641 92.5
R30083 vdd.n14615 vdd.n14614 92.5
R30084 vdd.n14566 vdd.n14565 92.5
R30085 vdd.n14548 vdd.n8184 92.5
R30086 vdd.n14560 vdd.n14559 92.5
R30087 vdd.n8197 vdd.n8186 92.5
R30088 vdd.n8236 vdd.n8224 92.5
R30089 vdd.n14468 vdd.n14467 92.5
R30090 vdd.n14439 vdd.n8235 92.5
R30091 vdd.n14376 vdd.n8273 92.5
R30092 vdd.n8314 vdd.n8297 92.5
R30093 vdd.n14381 vdd.n14380 92.5
R30094 vdd.n14361 vdd.n8313 92.5
R30095 vdd.n14373 vdd.n14372 92.5
R30096 vdd.n8357 vdd.n8316 92.5
R30097 vdd.n14301 vdd.n14300 92.5
R30098 vdd.n14284 vdd.n8368 92.5
R30099 vdd.n8392 vdd.n8370 92.5
R30100 vdd.n8422 vdd.n8407 92.5
R30101 vdd.n14224 vdd.n14223 92.5
R30102 vdd.n14206 vdd.n8421 92.5
R30103 vdd.n14218 vdd.n14217 92.5
R30104 vdd.n8470 vdd.n8424 92.5
R30105 vdd.n14159 vdd.n14158 92.5
R30106 vdd.n8525 vdd.n8488 92.5
R30107 vdd.n14096 vdd.n14095 92.5
R30108 vdd.n14079 vdd.n8537 92.5
R30109 vdd.n14091 vdd.n14090 92.5
R30110 vdd.n8576 vdd.n8539 92.5
R30111 vdd.n8590 vdd.n8574 92.5
R30112 vdd.n14011 vdd.n14010 92.5
R30113 vdd.n13993 vdd.n8589 92.5
R30114 vdd.n8614 vdd.n8592 92.5
R30115 vdd.n8643 vdd.n8629 92.5
R30116 vdd.n13934 vdd.n13933 92.5
R30117 vdd.n13916 vdd.n8642 92.5
R30118 vdd.n13928 vdd.n13927 92.5
R30119 vdd.n8693 vdd.n8645 92.5
R30120 vdd.n13870 vdd.n13869 92.5
R30121 vdd.n13820 vdd.n8711 92.5
R30122 vdd.n13809 vdd.n13808 92.5
R30123 vdd.n13792 vdd.n8750 92.5
R30124 vdd.n13804 vdd.n13803 92.5
R30125 vdd.n8785 vdd.n8752 92.5
R30126 vdd.n13736 vdd.n13735 92.5
R30127 vdd.n13719 vdd.n8797 92.5
R30128 vdd.n13731 vdd.n13730 92.5
R30129 vdd.n13613 vdd.n8824 92.5
R30130 vdd.n13614 vdd.n8842 92.5
R30131 vdd.n8906 vdd.n8851 92.5
R30132 vdd.n13619 vdd.n13618 92.5
R30133 vdd.n8905 vdd.n8884 92.5
R30134 vdd.n13609 vdd.n13608 92.5
R30135 vdd.n8930 vdd.n8908 92.5
R30136 vdd.n13529 vdd.n13528 92.5
R30137 vdd.n8965 vdd.n8949 92.5
R30138 vdd.n13522 vdd.n13521 92.5
R30139 vdd.n9004 vdd.n8968 92.5
R30140 vdd.n9017 vdd.n9002 92.5
R30141 vdd.n13445 vdd.n13444 92.5
R30142 vdd.n13427 vdd.n9016 92.5
R30143 vdd.n13439 vdd.n13438 92.5
R30144 vdd.n13321 vdd.n9045 92.5
R30145 vdd.n13322 vdd.n9062 92.5
R30146 vdd.n9127 vdd.n9071 92.5
R30147 vdd.n13327 vdd.n13326 92.5
R30148 vdd.n9126 vdd.n9105 92.5
R30149 vdd.n13317 vdd.n13316 92.5
R30150 vdd.n9151 vdd.n9129 92.5
R30151 vdd.n13237 vdd.n13236 92.5
R30152 vdd.n13218 vdd.n9186 92.5
R30153 vdd.n13230 vdd.n13229 92.5
R30154 vdd.n9225 vdd.n9189 92.5
R30155 vdd.n9241 vdd.n9222 92.5
R30156 vdd.n13152 vdd.n13151 92.5
R30157 vdd.n13133 vdd.n9240 92.5
R30158 vdd.n13146 vdd.n13145 92.5
R30159 vdd.n9243 vdd.n9242 92.5
R30160 vdd.n9277 vdd.n9243 92.5
R30161 vdd.n13147 vdd.n13146 92.5
R30162 vdd.n13148 vdd.n9240 92.5
R30163 vdd.n13151 vdd.n13150 92.5
R30164 vdd.n13149 vdd.n9241 92.5
R30165 vdd.n9189 vdd.n9188 92.5
R30166 vdd.n13231 vdd.n13230 92.5
R30167 vdd.n13232 vdd.n9186 92.5
R30168 vdd.n13236 vdd.n13235 92.5
R30169 vdd.n13234 vdd.n9187 92.5
R30170 vdd.n9187 vdd.n9165 92.5
R30171 vdd.n13233 vdd.n9159 92.5
R30172 vdd.n13276 vdd.n9159 92.5
R30173 vdd.n9129 vdd.n9128 92.5
R30174 vdd.n13318 vdd.n13317 92.5
R30175 vdd.n13319 vdd.n9126 92.5
R30176 vdd.n13326 vdd.n13325 92.5
R30177 vdd.n13324 vdd.n9127 92.5
R30178 vdd.n13323 vdd.n13322 92.5
R30179 vdd.n13321 vdd.n13320 92.5
R30180 vdd.n9019 vdd.n9018 92.5
R30181 vdd.n13389 vdd.n9019 92.5
R30182 vdd.n13440 vdd.n13439 92.5
R30183 vdd.n13441 vdd.n9016 92.5
R30184 vdd.n13444 vdd.n13443 92.5
R30185 vdd.n13442 vdd.n9017 92.5
R30186 vdd.n8968 vdd.n8967 92.5
R30187 vdd.n13523 vdd.n13522 92.5
R30188 vdd.n13524 vdd.n8965 92.5
R30189 vdd.n13528 vdd.n13527 92.5
R30190 vdd.n13526 vdd.n8966 92.5
R30191 vdd.n8966 vdd.n8944 92.5
R30192 vdd.n13525 vdd.n8937 92.5
R30193 vdd.n13568 vdd.n8937 92.5
R30194 vdd.n8908 vdd.n8907 92.5
R30195 vdd.n13610 vdd.n13609 92.5
R30196 vdd.n13611 vdd.n8905 92.5
R30197 vdd.n13618 vdd.n13617 92.5
R30198 vdd.n13616 vdd.n8906 92.5
R30199 vdd.n13615 vdd.n13614 92.5
R30200 vdd.n13613 vdd.n13612 92.5
R30201 vdd.n8799 vdd.n8798 92.5
R30202 vdd.n13681 vdd.n8799 92.5
R30203 vdd.n13732 vdd.n13731 92.5
R30204 vdd.n13733 vdd.n8797 92.5
R30205 vdd.n13735 vdd.n13734 92.5
R30206 vdd.n8752 vdd.n8751 92.5
R30207 vdd.n13805 vdd.n13804 92.5
R30208 vdd.n13806 vdd.n8750 92.5
R30209 vdd.n13808 vdd.n13807 92.5
R30210 vdd.n8711 vdd.n8710 92.5
R30211 vdd.n13866 vdd.n13865 92.5
R30212 vdd.n13865 vdd.n13864 92.5
R30213 vdd.n13867 vdd.n8709 92.5
R30214 vdd.n13856 vdd.n8709 92.5
R30215 vdd.n13869 vdd.n13868 92.5
R30216 vdd.n8645 vdd.n8644 92.5
R30217 vdd.n13929 vdd.n13928 92.5
R30218 vdd.n13930 vdd.n8642 92.5
R30219 vdd.n13933 vdd.n13932 92.5
R30220 vdd.n13931 vdd.n8643 92.5
R30221 vdd.n8592 vdd.n8591 92.5
R30222 vdd.n14006 vdd.n14005 92.5
R30223 vdd.n14005 vdd.n14004 92.5
R30224 vdd.n14007 vdd.n8589 92.5
R30225 vdd.n14010 vdd.n14009 92.5
R30226 vdd.n14008 vdd.n8590 92.5
R30227 vdd.n8539 vdd.n8538 92.5
R30228 vdd.n14092 vdd.n14091 92.5
R30229 vdd.n14093 vdd.n8537 92.5
R30230 vdd.n14095 vdd.n14094 92.5
R30231 vdd.n8488 vdd.n8487 92.5
R30232 vdd.n14155 vdd.n14154 92.5
R30233 vdd.n14154 vdd.n14153 92.5
R30234 vdd.n14156 vdd.n8486 92.5
R30235 vdd.n14145 vdd.n8486 92.5
R30236 vdd.n14158 vdd.n14157 92.5
R30237 vdd.n8424 vdd.n8423 92.5
R30238 vdd.n14219 vdd.n14218 92.5
R30239 vdd.n14220 vdd.n8421 92.5
R30240 vdd.n14223 vdd.n14222 92.5
R30241 vdd.n14221 vdd.n8422 92.5
R30242 vdd.n8370 vdd.n8369 92.5
R30243 vdd.n14297 vdd.n14296 92.5
R30244 vdd.n14296 vdd.n14295 92.5
R30245 vdd.n14298 vdd.n8368 92.5
R30246 vdd.n14300 vdd.n14299 92.5
R30247 vdd.n8316 vdd.n8315 92.5
R30248 vdd.n14374 vdd.n14373 92.5
R30249 vdd.n14375 vdd.n8313 92.5
R30250 vdd.n14380 vdd.n14379 92.5
R30251 vdd.n14378 vdd.n8314 92.5
R30252 vdd.n14377 vdd.n14376 92.5
R30253 vdd.n8238 vdd.n8237 92.5
R30254 vdd.n14419 vdd.n8238 92.5
R30255 vdd.n14463 vdd.n14462 92.5
R30256 vdd.n14462 vdd.n14461 92.5
R30257 vdd.n14464 vdd.n8235 92.5
R30258 vdd.n14467 vdd.n14466 92.5
R30259 vdd.n14465 vdd.n8236 92.5
R30260 vdd.n8186 vdd.n8185 92.5
R30261 vdd.n14561 vdd.n14560 92.5
R30262 vdd.n14562 vdd.n8184 92.5
R30263 vdd.n14565 vdd.n14564 92.5
R30264 vdd.n14563 vdd.n8171 92.5
R30265 vdd.n14567 vdd.n8171 92.5
R30266 vdd.n14615 vdd.n8170 92.5
R30267 vdd.n11629 vdd.n11577 92.5
R30268 vdd.n11629 vdd.n11628 92.5
R30269 vdd.n11656 vdd.n11655 92.5
R30270 vdd.n11654 vdd.n11574 92.5
R30271 vdd.n11653 vdd.n11652 92.5
R30272 vdd.n11651 vdd.n11650 92.5
R30273 vdd.n11649 vdd.n11648 92.5
R30274 vdd.n11647 vdd.n11646 92.5
R30275 vdd.n11645 vdd.n11644 92.5
R30276 vdd.n11643 vdd.n11642 92.5
R30277 vdd.n11641 vdd.n11640 92.5
R30278 vdd.n11639 vdd.n11638 92.5
R30279 vdd.n11637 vdd.n11636 92.5
R30280 vdd.n11635 vdd.n11634 92.5
R30281 vdd.n11633 vdd.n11632 92.5
R30282 vdd.n11631 vdd.n11630 92.5
R30283 vdd.n10476 vdd.n10475 92.5
R30284 vdd.n10469 vdd.n10277 92.5
R30285 vdd.n10470 vdd.n10469 92.5
R30286 vdd.n10464 vdd.n10463 92.5
R30287 vdd.n10465 vdd.n10464 92.5
R30288 vdd.n10454 vdd.n10289 92.5
R30289 vdd.n10289 vdd.n10288 92.5
R30290 vdd.n10294 vdd.n10291 92.5
R30291 vdd.n10291 vdd.n10290 92.5
R30292 vdd.n10445 vdd.n10444 92.5
R30293 vdd.n10444 vdd.n10443 92.5
R30294 vdd.n10440 vdd.n10439 92.5
R30295 vdd.n10441 vdd.n10440 92.5
R30296 vdd.n10430 vdd.n10306 92.5
R30297 vdd.n10306 vdd.n10305 92.5
R30298 vdd.n10317 vdd.n10316 92.5
R30299 vdd.n10318 vdd.n10317 92.5
R30300 vdd.n10416 vdd.n10315 92.5
R30301 vdd.n10315 vdd.n10312 92.5
R30302 vdd.n10407 vdd.n10406 92.5
R30303 vdd.n10406 vdd.n10405 92.5
R30304 vdd.n10327 vdd.n10326 92.5
R30305 vdd.n10330 vdd.n10327 92.5
R30306 vdd.n10391 vdd.n10334 92.5
R30307 vdd.n10393 vdd.n10391 92.5
R30308 vdd.n10479 vdd.n10270 92.5
R30309 vdd.n10270 vdd.n10269 92.5
R30310 vdd.n10488 vdd.n10487 92.5
R30311 vdd.n10121 vdd.n10119 92.5
R30312 vdd.n10241 vdd.n10240 92.5
R30313 vdd.n10239 vdd.n10237 92.5
R30314 vdd.n12597 vdd.n12596 92.5
R30315 vdd.n12596 vdd.n12595 92.5
R30316 vdd.n10109 vdd.n10104 92.5
R30317 vdd.n12604 vdd.n12603 92.5
R30318 vdd.n12604 vdd.n10062 92.5
R30319 vdd.n10192 vdd.n10191 92.5
R30320 vdd.n10193 vdd.n10192 92.5
R30321 vdd.n10185 vdd.n10141 92.5
R30322 vdd.n10141 vdd.n10139 92.5
R30323 vdd.n12617 vdd.n12616 92.5
R30324 vdd.n12616 vdd.n12615 92.5
R30325 vdd.n12625 vdd.n12624 92.5
R30326 vdd.n12626 vdd.n12625 92.5
R30327 vdd.n10146 vdd.n10048 92.5
R30328 vdd.n10155 vdd.n10048 92.5
R30329 vdd.n10387 vdd.n10386 92.5
R30330 vdd.n10386 vdd.n10385 92.5
R30331 vdd.n10343 vdd.n10342 92.5
R30332 vdd.n10380 vdd.n10343 92.5
R30333 vdd.n10357 vdd.n10355 92.5
R30334 vdd.n10355 vdd.n10353 92.5
R30335 vdd.n10367 vdd.n10366 92.5
R30336 vdd.n10368 vdd.n10367 92.5
R30337 vdd.n9292 vdd.n9290 92.5
R30338 vdd.n13077 vdd.n9292 92.5
R30339 vdd.n13070 vdd.n13069 92.5
R30340 vdd.n13071 vdd.n13070 92.5
R30341 vdd.n13060 vdd.n9307 92.5
R30342 vdd.n9307 vdd.n9306 92.5
R30343 vdd.n9315 vdd.n9313 92.5
R30344 vdd.n9317 vdd.n9315 92.5
R30345 vdd.n9341 vdd.n9340 92.5
R30346 vdd.n9340 vdd.n9335 92.5
R30347 vdd.n9347 vdd.n9330 92.5
R30348 vdd.n9330 vdd.n9328 92.5
R30349 vdd.n13041 vdd.n13040 92.5
R30350 vdd.n13042 vdd.n13041 92.5
R30351 vdd.n13034 vdd.n13033 92.5
R30352 vdd.n13033 vdd.n13032 92.5
R30353 vdd.n9369 vdd.n9368 92.5
R30354 vdd.n9370 vdd.n9369 92.5
R30355 vdd.n9388 vdd.n9387 92.5
R30356 vdd.n9387 vdd.n9386 92.5
R30357 vdd.n9362 vdd.n9360 92.5
R30358 vdd.n9364 vdd.n9362 92.5
R30359 vdd.n9398 vdd.n9395 92.5
R30360 vdd.n13013 vdd.n9398 92.5
R30361 vdd.n13003 vdd.n9407 92.5
R30362 vdd.n13004 vdd.n13003 92.5
R30363 vdd.n9432 vdd.n9431 92.5
R30364 vdd.n9435 vdd.n9432 92.5
R30365 vdd.n9439 vdd.n9438 92.5
R30366 vdd.n9438 vdd.n9437 92.5
R30367 vdd.n12990 vdd.n9417 92.5
R30368 vdd.n9417 vdd.n9415 92.5
R30369 vdd.n12984 vdd.n12983 92.5
R30370 vdd.n12983 vdd.n12982 92.5
R30371 vdd.n9453 vdd.n9452 92.5
R30372 vdd.n12973 vdd.n9453 92.5
R30373 vdd.n9465 vdd.n9462 92.5
R30374 vdd.n9462 vdd.n9460 92.5
R30375 vdd.n9485 vdd.n9484 92.5
R30376 vdd.n9484 vdd.n9483 92.5
R30377 vdd.n9500 vdd.n9499 92.5
R30378 vdd.n9501 vdd.n9500 92.5
R30379 vdd.n12952 vdd.n9477 92.5
R30380 vdd.n9477 vdd.n9475 92.5
R30381 vdd.n12946 vdd.n12945 92.5
R30382 vdd.n12945 vdd.n12944 92.5
R30383 vdd.n12938 vdd.n12937 92.5
R30384 vdd.n12937 vdd.n12936 92.5
R30385 vdd.n9531 vdd.n9517 92.5
R30386 vdd.n9519 vdd.n9517 92.5
R30387 vdd.n9543 vdd.n9542 92.5
R30388 vdd.n9542 vdd.n9541 92.5
R30389 vdd.n9527 vdd.n9525 92.5
R30390 vdd.n9529 vdd.n9527 92.5
R30391 vdd.n9553 vdd.n9550 92.5
R30392 vdd.n12918 vdd.n9553 92.5
R30393 vdd.n12908 vdd.n9562 92.5
R30394 vdd.n12909 vdd.n12908 92.5
R30395 vdd.n9581 vdd.n9580 92.5
R30396 vdd.n9580 vdd.n9579 92.5
R30397 vdd.n9597 vdd.n9596 92.5
R30398 vdd.n9598 vdd.n9597 92.5
R30399 vdd.n9575 vdd.n9573 92.5
R30400 vdd.n9573 vdd.n9571 92.5
R30401 vdd.n12888 vdd.n9607 92.5
R30402 vdd.n9607 vdd.n9605 92.5
R30403 vdd.n12883 vdd.n12882 92.5
R30404 vdd.n12882 vdd.n12881 92.5
R30405 vdd.n9631 vdd.n9630 92.5
R30406 vdd.n9632 vdd.n9631 92.5
R30407 vdd.n9651 vdd.n9650 92.5
R30408 vdd.n9650 vdd.n9649 92.5
R30409 vdd.n9624 vdd.n9622 92.5
R30410 vdd.n12869 vdd.n9624 92.5
R30411 vdd.n12862 vdd.n12861 92.5
R30412 vdd.n12863 vdd.n12862 92.5
R30413 vdd.n12852 vdd.n9667 92.5
R30414 vdd.n9667 vdd.n9666 92.5
R30415 vdd.n9676 vdd.n9674 92.5
R30416 vdd.n9679 vdd.n9676 92.5
R30417 vdd.n9701 vdd.n9700 92.5
R30418 vdd.n9700 vdd.n9695 92.5
R30419 vdd.n9707 vdd.n9690 92.5
R30420 vdd.n9690 vdd.n9688 92.5
R30421 vdd.n12833 vdd.n12832 92.5
R30422 vdd.n12834 vdd.n12833 92.5
R30423 vdd.n12826 vdd.n12825 92.5
R30424 vdd.n12825 vdd.n12824 92.5
R30425 vdd.n9729 vdd.n9728 92.5
R30426 vdd.n9730 vdd.n9729 92.5
R30427 vdd.n9748 vdd.n9747 92.5
R30428 vdd.n9747 vdd.n9746 92.5
R30429 vdd.n9722 vdd.n9720 92.5
R30430 vdd.n9724 vdd.n9722 92.5
R30431 vdd.n9758 vdd.n9755 92.5
R30432 vdd.n12805 vdd.n9758 92.5
R30433 vdd.n12795 vdd.n9767 92.5
R30434 vdd.n12796 vdd.n12795 92.5
R30435 vdd.n9792 vdd.n9791 92.5
R30436 vdd.n9794 vdd.n9792 92.5
R30437 vdd.n9798 vdd.n9797 92.5
R30438 vdd.n9797 vdd.n9796 92.5
R30439 vdd.n12782 vdd.n9778 92.5
R30440 vdd.n9778 vdd.n9776 92.5
R30441 vdd.n12776 vdd.n12775 92.5
R30442 vdd.n12775 vdd.n12774 92.5
R30443 vdd.n9812 vdd.n9811 92.5
R30444 vdd.n12765 vdd.n9812 92.5
R30445 vdd.n9825 vdd.n9822 92.5
R30446 vdd.n9822 vdd.n9820 92.5
R30447 vdd.n9845 vdd.n9844 92.5
R30448 vdd.n9844 vdd.n9843 92.5
R30449 vdd.n9860 vdd.n9859 92.5
R30450 vdd.n9861 vdd.n9860 92.5
R30451 vdd.n12744 vdd.n9837 92.5
R30452 vdd.n9837 vdd.n9835 92.5
R30453 vdd.n12738 vdd.n12737 92.5
R30454 vdd.n12737 vdd.n12736 92.5
R30455 vdd.n12730 vdd.n12729 92.5
R30456 vdd.n12729 vdd.n12728 92.5
R30457 vdd.n9892 vdd.n9877 92.5
R30458 vdd.n9879 vdd.n9877 92.5
R30459 vdd.n9903 vdd.n9902 92.5
R30460 vdd.n9902 vdd.n9901 92.5
R30461 vdd.n9888 vdd.n9886 92.5
R30462 vdd.n9890 vdd.n9888 92.5
R30463 vdd.n9913 vdd.n9910 92.5
R30464 vdd.n12710 vdd.n9913 92.5
R30465 vdd.n12700 vdd.n9920 92.5
R30466 vdd.n12701 vdd.n12700 92.5
R30467 vdd.n9941 vdd.n9940 92.5
R30468 vdd.n9940 vdd.n9939 92.5
R30469 vdd.n9957 vdd.n9956 92.5
R30470 vdd.n9958 vdd.n9957 92.5
R30471 vdd.n9934 vdd.n9932 92.5
R30472 vdd.n9932 vdd.n9930 92.5
R30473 vdd.n12680 vdd.n9967 92.5
R30474 vdd.n9967 vdd.n9965 92.5
R30475 vdd.n12675 vdd.n12674 92.5
R30476 vdd.n12674 vdd.n12673 92.5
R30477 vdd.n9991 vdd.n9990 92.5
R30478 vdd.n9992 vdd.n9991 92.5
R30479 vdd.n10011 vdd.n10010 92.5
R30480 vdd.n10010 vdd.n10009 92.5
R30481 vdd.n9984 vdd.n9982 92.5
R30482 vdd.n12661 vdd.n9984 92.5
R30483 vdd.n12654 vdd.n12653 92.5
R30484 vdd.n12655 vdd.n12654 92.5
R30485 vdd.n12644 vdd.n10027 92.5
R30486 vdd.n10027 vdd.n10026 92.5
R30487 vdd.n10036 vdd.n10034 92.5
R30488 vdd.n10039 vdd.n10036 92.5
R30489 vdd.n10153 vdd.n10152 92.5
R30490 vdd.n10154 vdd.n10153 92.5
R30491 vdd.n12528 vdd.n10517 92.5
R30492 vdd.n10544 vdd.n10524 92.5
R30493 vdd.n12519 vdd.n10524 92.5
R30494 vdd.n10536 vdd.n10535 92.5
R30495 vdd.n10553 vdd.n10536 92.5
R30496 vdd.n12512 vdd.n12511 92.5
R30497 vdd.n12513 vdd.n12512 92.5
R30498 vdd.n10563 vdd.n10562 92.5
R30499 vdd.n12502 vdd.n10563 92.5
R30500 vdd.n10576 vdd.n10575 92.5
R30501 vdd.n10577 vdd.n10576 92.5
R30502 vdd.n10572 vdd.n10569 92.5
R30503 vdd.n12488 vdd.n10572 92.5
R30504 vdd.n12481 vdd.n12480 92.5
R30505 vdd.n12482 vdd.n12481 92.5
R30506 vdd.n10604 vdd.n10603 92.5
R30507 vdd.n12471 vdd.n10604 92.5
R30508 vdd.n10612 vdd.n10610 92.5
R30509 vdd.n10614 vdd.n10612 92.5
R30510 vdd.n10637 vdd.n10616 92.5
R30511 vdd.n12459 vdd.n10616 92.5
R30512 vdd.n10631 vdd.n10629 92.5
R30513 vdd.n10646 vdd.n10631 92.5
R30514 vdd.n12452 vdd.n12451 92.5
R30515 vdd.n12453 vdd.n12452 92.5
R30516 vdd.n10655 vdd.n10654 92.5
R30517 vdd.n12442 vdd.n10655 92.5
R30518 vdd.n10663 vdd.n10661 92.5
R30519 vdd.n10665 vdd.n10663 92.5
R30520 vdd.n10681 vdd.n10664 92.5
R30521 vdd.n12431 vdd.n10664 92.5
R30522 vdd.n10679 vdd.n10678 92.5
R30523 vdd.n10689 vdd.n10679 92.5
R30524 vdd.n12424 vdd.n12423 92.5
R30525 vdd.n12425 vdd.n12424 92.5
R30526 vdd.n10699 vdd.n10698 92.5
R30527 vdd.n12414 vdd.n10699 92.5
R30528 vdd.n10712 vdd.n10711 92.5
R30529 vdd.n10713 vdd.n10712 92.5
R30530 vdd.n10707 vdd.n10704 92.5
R30531 vdd.n12400 vdd.n10707 92.5
R30532 vdd.n10727 vdd.n10726 92.5
R30533 vdd.n10738 vdd.n10727 92.5
R30534 vdd.n12393 vdd.n12392 92.5
R30535 vdd.n12394 vdd.n12393 92.5
R30536 vdd.n10748 vdd.n10747 92.5
R30537 vdd.n12383 vdd.n10748 92.5
R30538 vdd.n10755 vdd.n10753 92.5
R30539 vdd.n10763 vdd.n10755 92.5
R30540 vdd.n10788 vdd.n10765 92.5
R30541 vdd.n12370 vdd.n10765 92.5
R30542 vdd.n10782 vdd.n10780 92.5
R30543 vdd.n10797 vdd.n10782 92.5
R30544 vdd.n12363 vdd.n12362 92.5
R30545 vdd.n12364 vdd.n12363 92.5
R30546 vdd.n10806 vdd.n10805 92.5
R30547 vdd.n12353 vdd.n10806 92.5
R30548 vdd.n10814 vdd.n10812 92.5
R30549 vdd.n10816 vdd.n10814 92.5
R30550 vdd.n10832 vdd.n10818 92.5
R30551 vdd.n12341 vdd.n10818 92.5
R30552 vdd.n10847 vdd.n10846 92.5
R30553 vdd.n10846 vdd.n10845 92.5
R30554 vdd.n12334 vdd.n12333 92.5
R30555 vdd.n12335 vdd.n12334 92.5
R30556 vdd.n10859 vdd.n10858 92.5
R30557 vdd.n10860 vdd.n10859 92.5
R30558 vdd.n10857 vdd.n10854 92.5
R30559 vdd.n12323 vdd.n10857 92.5
R30560 vdd.n10874 vdd.n10873 92.5
R30561 vdd.n10885 vdd.n10874 92.5
R30562 vdd.n12316 vdd.n12315 92.5
R30563 vdd.n12317 vdd.n12316 92.5
R30564 vdd.n10895 vdd.n10894 92.5
R30565 vdd.n12306 vdd.n10895 92.5
R30566 vdd.n10908 vdd.n10907 92.5
R30567 vdd.n10909 vdd.n10908 92.5
R30568 vdd.n10904 vdd.n10901 92.5
R30569 vdd.n12292 vdd.n10904 92.5
R30570 vdd.n10939 vdd.n10927 92.5
R30571 vdd.n10939 vdd.n10938 92.5
R30572 vdd.n12281 vdd.n12280 92.5
R30573 vdd.n12280 vdd.n12279 92.5
R30574 vdd.n12274 vdd.n10923 92.5
R30575 vdd.n10923 vdd.n10922 92.5
R30576 vdd.n10975 vdd.n10953 92.5
R30577 vdd.n12269 vdd.n10953 92.5
R30578 vdd.n10968 vdd.n10966 92.5
R30579 vdd.n10984 vdd.n10968 92.5
R30580 vdd.n12262 vdd.n12261 92.5
R30581 vdd.n12263 vdd.n12262 92.5
R30582 vdd.n10993 vdd.n10992 92.5
R30583 vdd.n12252 vdd.n10993 92.5
R30584 vdd.n11001 vdd.n10999 92.5
R30585 vdd.n11003 vdd.n11001 92.5
R30586 vdd.n11019 vdd.n11005 92.5
R30587 vdd.n12240 vdd.n11005 92.5
R30588 vdd.n11030 vdd.n11029 92.5
R30589 vdd.n11029 vdd.n11028 92.5
R30590 vdd.n12233 vdd.n12232 92.5
R30591 vdd.n12234 vdd.n12233 92.5
R30592 vdd.n11036 vdd.n11035 92.5
R30593 vdd.n12223 vdd.n11036 92.5
R30594 vdd.n11049 vdd.n11048 92.5
R30595 vdd.n11050 vdd.n11049 92.5
R30596 vdd.n11044 vdd.n11041 92.5
R30597 vdd.n12209 vdd.n11044 92.5
R30598 vdd.n11064 vdd.n11063 92.5
R30599 vdd.n11075 vdd.n11064 92.5
R30600 vdd.n12202 vdd.n12201 92.5
R30601 vdd.n12203 vdd.n12202 92.5
R30602 vdd.n11085 vdd.n11084 92.5
R30603 vdd.n12192 vdd.n11085 92.5
R30604 vdd.n11098 vdd.n11097 92.5
R30605 vdd.n11099 vdd.n11098 92.5
R30606 vdd.n11114 vdd.n11112 92.5
R30607 vdd.n11118 vdd.n11114 92.5
R30608 vdd.n12172 vdd.n12171 92.5
R30609 vdd.n12173 vdd.n12172 92.5
R30610 vdd.n11127 vdd.n11126 92.5
R30611 vdd.n12162 vdd.n11127 92.5
R30612 vdd.n11135 vdd.n11133 92.5
R30613 vdd.n11137 vdd.n11135 92.5
R30614 vdd.n11160 vdd.n11139 92.5
R30615 vdd.n12150 vdd.n11139 92.5
R30616 vdd.n11154 vdd.n11152 92.5
R30617 vdd.n11169 vdd.n11154 92.5
R30618 vdd.n12143 vdd.n12142 92.5
R30619 vdd.n12144 vdd.n12143 92.5
R30620 vdd.n11177 vdd.n11176 92.5
R30621 vdd.n12133 vdd.n11177 92.5
R30622 vdd.n11181 vdd.n11178 92.5
R30623 vdd.n11184 vdd.n11178 92.5
R30624 vdd.n11183 vdd.n11182 92.5
R30625 vdd.n12121 vdd.n11183 92.5
R30626 vdd.n11199 vdd.n11198 92.5
R30627 vdd.n11210 vdd.n11199 92.5
R30628 vdd.n12114 vdd.n12113 92.5
R30629 vdd.n12115 vdd.n12114 92.5
R30630 vdd.n11220 vdd.n11219 92.5
R30631 vdd.n12104 vdd.n11220 92.5
R30632 vdd.n11233 vdd.n11232 92.5
R30633 vdd.n11234 vdd.n11233 92.5
R30634 vdd.n11229 vdd.n11226 92.5
R30635 vdd.n12090 vdd.n11229 92.5
R30636 vdd.n11248 vdd.n11247 92.5
R30637 vdd.n11259 vdd.n11248 92.5
R30638 vdd.n12083 vdd.n12082 92.5
R30639 vdd.n12084 vdd.n12083 92.5
R30640 vdd.n12069 vdd.n11270 92.5
R30641 vdd.n11273 vdd.n11270 92.5
R30642 vdd.n11297 vdd.n11275 92.5
R30643 vdd.n12064 vdd.n11275 92.5
R30644 vdd.n11290 vdd.n11288 92.5
R30645 vdd.n11306 vdd.n11290 92.5
R30646 vdd.n12057 vdd.n12056 92.5
R30647 vdd.n12058 vdd.n12057 92.5
R30648 vdd.n11315 vdd.n11314 92.5
R30649 vdd.n12047 vdd.n11315 92.5
R30650 vdd.n11323 vdd.n11321 92.5
R30651 vdd.n11325 vdd.n11323 92.5
R30652 vdd.n11341 vdd.n11327 92.5
R30653 vdd.n12035 vdd.n11327 92.5
R30654 vdd.n11356 vdd.n11355 92.5
R30655 vdd.n11355 vdd.n11354 92.5
R30656 vdd.n12028 vdd.n12027 92.5
R30657 vdd.n12029 vdd.n12028 92.5
R30658 vdd.n11368 vdd.n11367 92.5
R30659 vdd.n11369 vdd.n11368 92.5
R30660 vdd.n11366 vdd.n11363 92.5
R30661 vdd.n12017 vdd.n11366 92.5
R30662 vdd.n11383 vdd.n11382 92.5
R30663 vdd.n11394 vdd.n11383 92.5
R30664 vdd.n12010 vdd.n12009 92.5
R30665 vdd.n12011 vdd.n12010 92.5
R30666 vdd.n11404 vdd.n11403 92.5
R30667 vdd.n12000 vdd.n11404 92.5
R30668 vdd.n11417 vdd.n11416 92.5
R30669 vdd.n11418 vdd.n11417 92.5
R30670 vdd.n11413 vdd.n11410 92.5
R30671 vdd.n11986 vdd.n11413 92.5
R30672 vdd.n11483 vdd.n11471 92.5
R30673 vdd.n11483 vdd.n11482 92.5
R30674 vdd.n11975 vdd.n11974 92.5
R30675 vdd.n11974 vdd.n11973 92.5
R30676 vdd.n11968 vdd.n11432 92.5
R30677 vdd.n11432 vdd.n11431 92.5
R30678 vdd.n11504 vdd.n11438 92.5
R30679 vdd.n11963 vdd.n11438 92.5
R30680 vdd.n11530 vdd.n11529 92.5
R30681 vdd.n11529 vdd.n11528 92.5
R30682 vdd.n11956 vdd.n11955 92.5
R30683 vdd.n11957 vdd.n11956 92.5
R30684 vdd.n11548 vdd.n11547 92.5
R30685 vdd.n11945 vdd.n11548 92.5
R30686 vdd.n11935 vdd.n11934 92.5
R30687 vdd.n11934 vdd.n11933 92.5
R30688 vdd.n12524 vdd.n10519 92.5
R30689 vdd.n10519 vdd.n10518 92.5
R30690 vdd.n11921 vdd.n11661 92.5
R30691 vdd.n11661 vdd.n11660 92.5
R30692 vdd.n13083 vdd.n13082 92.5
R30693 vdd.n13082 vdd.n13081 92.5
R30694 vdd.n9288 vdd.n9286 92.5
R30695 vdd.n13073 vdd.n9288 92.5
R30696 vdd.n9324 vdd.n9323 92.5
R30697 vdd.n9323 vdd.n9308 92.5
R30698 vdd.n9325 vdd.n9321 92.5
R30699 vdd.n9321 vdd.n9320 92.5
R30700 vdd.n13048 vdd.n13047 92.5
R30701 vdd.n13049 vdd.n13048 92.5
R30702 vdd.n13046 vdd.n9322 92.5
R30703 vdd.n9342 vdd.n9322 92.5
R30704 vdd.n13045 vdd.n13044 92.5
R30705 vdd.n13044 vdd.n13043 92.5
R30706 vdd.n9327 vdd.n9326 92.5
R30707 vdd.n9329 vdd.n9327 92.5
R30708 vdd.n13029 vdd.n13028 92.5
R30709 vdd.n13030 vdd.n13029 92.5
R30710 vdd.n13027 vdd.n9356 92.5
R30711 vdd.n9384 vdd.n9356 92.5
R30712 vdd.n13026 vdd.n13025 92.5
R30713 vdd.n13025 vdd.n13024 92.5
R30714 vdd.n9358 vdd.n9357 92.5
R30715 vdd.n9400 vdd.n9358 92.5
R30716 vdd.n9411 vdd.n9409 92.5
R30717 vdd.n9409 vdd.n9401 92.5
R30718 vdd.n12999 vdd.n12998 92.5
R30719 vdd.n13000 vdd.n12999 92.5
R30720 vdd.n12997 vdd.n9410 92.5
R30721 vdd.n9441 vdd.n9410 92.5
R30722 vdd.n12996 vdd.n12995 92.5
R30723 vdd.n12995 vdd.n12994 92.5
R30724 vdd.n9413 vdd.n9412 92.5
R30725 vdd.n12986 vdd.n9413 92.5
R30726 vdd.n9470 vdd.n9469 92.5
R30727 vdd.n9469 vdd.n9454 92.5
R30728 vdd.n9471 vdd.n9467 92.5
R30729 vdd.n9467 vdd.n9455 92.5
R30730 vdd.n12961 vdd.n12960 92.5
R30731 vdd.n12962 vdd.n12961 92.5
R30732 vdd.n12959 vdd.n9468 92.5
R30733 vdd.n9497 vdd.n9468 92.5
R30734 vdd.n12958 vdd.n12957 92.5
R30735 vdd.n12957 vdd.n12956 92.5
R30736 vdd.n9473 vdd.n9472 92.5
R30737 vdd.n12948 vdd.n9473 92.5
R30738 vdd.n9522 vdd.n9520 92.5
R30739 vdd.n9520 vdd.n9518 92.5
R30740 vdd.n12934 vdd.n12933 92.5
R30741 vdd.n12935 vdd.n12934 92.5
R30742 vdd.n12932 vdd.n9521 92.5
R30743 vdd.n9538 vdd.n9521 92.5
R30744 vdd.n12931 vdd.n12930 92.5
R30745 vdd.n12930 vdd.n12929 92.5
R30746 vdd.n9524 vdd.n9523 92.5
R30747 vdd.n9555 vdd.n9524 92.5
R30748 vdd.n9567 vdd.n9565 92.5
R30749 vdd.n9565 vdd.n9556 92.5
R30750 vdd.n12904 vdd.n12903 92.5
R30751 vdd.n12905 vdd.n12904 92.5
R30752 vdd.n12902 vdd.n9566 92.5
R30753 vdd.n9594 vdd.n9566 92.5
R30754 vdd.n12901 vdd.n12900 92.5
R30755 vdd.n12900 vdd.n12899 92.5
R30756 vdd.n9569 vdd.n9568 92.5
R30757 vdd.n9609 vdd.n9569 92.5
R30758 vdd.n9618 vdd.n9616 92.5
R30759 vdd.n9616 vdd.n9610 92.5
R30760 vdd.n12878 vdd.n12877 92.5
R30761 vdd.n12879 vdd.n12878 92.5
R30762 vdd.n12876 vdd.n9617 92.5
R30763 vdd.n9647 vdd.n9617 92.5
R30764 vdd.n12875 vdd.n12874 92.5
R30765 vdd.n12874 vdd.n12873 92.5
R30766 vdd.n9620 vdd.n9619 92.5
R30767 vdd.n12865 vdd.n9620 92.5
R30768 vdd.n9684 vdd.n9683 92.5
R30769 vdd.n9683 vdd.n9668 92.5
R30770 vdd.n9685 vdd.n9681 92.5
R30771 vdd.n9681 vdd.n9669 92.5
R30772 vdd.n12840 vdd.n12839 92.5
R30773 vdd.n12841 vdd.n12840 92.5
R30774 vdd.n12838 vdd.n9682 92.5
R30775 vdd.n9702 vdd.n9682 92.5
R30776 vdd.n12837 vdd.n12836 92.5
R30777 vdd.n12836 vdd.n12835 92.5
R30778 vdd.n9687 vdd.n9686 92.5
R30779 vdd.n9689 vdd.n9687 92.5
R30780 vdd.n12821 vdd.n12820 92.5
R30781 vdd.n12822 vdd.n12821 92.5
R30782 vdd.n12819 vdd.n9716 92.5
R30783 vdd.n9744 vdd.n9716 92.5
R30784 vdd.n12818 vdd.n12817 92.5
R30785 vdd.n12817 vdd.n12816 92.5
R30786 vdd.n9718 vdd.n9717 92.5
R30787 vdd.n9760 vdd.n9718 92.5
R30788 vdd.n9772 vdd.n9770 92.5
R30789 vdd.n9770 vdd.n9761 92.5
R30790 vdd.n12791 vdd.n12790 92.5
R30791 vdd.n12792 vdd.n12791 92.5
R30792 vdd.n12789 vdd.n9771 92.5
R30793 vdd.n9800 vdd.n9771 92.5
R30794 vdd.n12788 vdd.n12787 92.5
R30795 vdd.n12787 vdd.n12786 92.5
R30796 vdd.n9774 vdd.n9773 92.5
R30797 vdd.n12778 vdd.n9774 92.5
R30798 vdd.n9830 vdd.n9829 92.5
R30799 vdd.n9829 vdd.n9814 92.5
R30800 vdd.n9831 vdd.n9827 92.5
R30801 vdd.n9827 vdd.n9815 92.5
R30802 vdd.n12753 vdd.n12752 92.5
R30803 vdd.n12754 vdd.n12753 92.5
R30804 vdd.n12751 vdd.n9828 92.5
R30805 vdd.n9857 vdd.n9828 92.5
R30806 vdd.n12750 vdd.n12749 92.5
R30807 vdd.n12749 vdd.n12748 92.5
R30808 vdd.n9833 vdd.n9832 92.5
R30809 vdd.n12740 vdd.n9833 92.5
R30810 vdd.n9882 vdd.n9880 92.5
R30811 vdd.n9880 vdd.n9878 92.5
R30812 vdd.n12726 vdd.n12725 92.5
R30813 vdd.n12727 vdd.n12726 92.5
R30814 vdd.n12724 vdd.n9881 92.5
R30815 vdd.n9899 vdd.n9881 92.5
R30816 vdd.n12723 vdd.n12722 92.5
R30817 vdd.n12722 vdd.n12721 92.5
R30818 vdd.n9884 vdd.n9883 92.5
R30819 vdd.n9915 vdd.n9884 92.5
R30820 vdd.n9926 vdd.n9924 92.5
R30821 vdd.n9924 vdd.n9923 92.5
R30822 vdd.n12696 vdd.n12695 92.5
R30823 vdd.n12697 vdd.n12696 92.5
R30824 vdd.n12694 vdd.n9925 92.5
R30825 vdd.n9954 vdd.n9925 92.5
R30826 vdd.n12693 vdd.n12692 92.5
R30827 vdd.n12692 vdd.n12691 92.5
R30828 vdd.n9928 vdd.n9927 92.5
R30829 vdd.n9969 vdd.n9928 92.5
R30830 vdd.n9978 vdd.n9976 92.5
R30831 vdd.n9976 vdd.n9970 92.5
R30832 vdd.n12670 vdd.n12669 92.5
R30833 vdd.n12671 vdd.n12670 92.5
R30834 vdd.n12668 vdd.n9977 92.5
R30835 vdd.n10007 vdd.n9977 92.5
R30836 vdd.n12667 vdd.n12666 92.5
R30837 vdd.n12666 vdd.n12665 92.5
R30838 vdd.n9980 vdd.n9979 92.5
R30839 vdd.n12657 vdd.n9980 92.5
R30840 vdd.n10043 vdd.n10042 92.5
R30841 vdd.n10042 vdd.n10028 92.5
R30842 vdd.n10044 vdd.n10040 92.5
R30843 vdd.n10040 vdd.n10029 92.5
R30844 vdd.n12632 vdd.n12631 92.5
R30845 vdd.n12633 vdd.n12632 92.5
R30846 vdd.n12630 vdd.n10041 92.5
R30847 vdd.n10156 vdd.n10041 92.5
R30848 vdd.n12629 vdd.n12628 92.5
R30849 vdd.n12628 vdd.n12627 92.5
R30850 vdd.n10046 vdd.n10045 92.5
R30851 vdd.n10047 vdd.n10046 92.5
R30852 vdd.n12612 vdd.n12611 92.5
R30853 vdd.n12613 vdd.n12612 92.5
R30854 vdd.n12610 vdd.n10058 92.5
R30855 vdd.n10189 vdd.n10058 92.5
R30856 vdd.n12609 vdd.n12608 92.5
R30857 vdd.n12608 vdd.n12607 92.5
R30858 vdd.n10060 vdd.n10059 92.5
R30859 vdd.n10106 vdd.n10060 92.5
R30860 vdd.n10115 vdd.n10113 92.5
R30861 vdd.n10113 vdd.n10112 92.5
R30862 vdd.n12593 vdd.n12592 92.5
R30863 vdd.n12594 vdd.n12593 92.5
R30864 vdd.n12591 vdd.n10114 92.5
R30865 vdd.n10243 vdd.n10114 92.5
R30866 vdd.n12590 vdd.n12589 92.5
R30867 vdd.n12589 vdd.n12588 92.5
R30868 vdd.n10117 vdd.n10116 92.5
R30869 vdd.n10485 vdd.n10117 92.5
R30870 vdd.n10497 vdd.n10495 92.5
R30871 vdd.n10495 vdd.n10494 92.5
R30872 vdd.n12565 vdd.n12564 92.5
R30873 vdd.n12566 vdd.n12565 92.5
R30874 vdd.n12563 vdd.n10496 92.5
R30875 vdd.n10500 vdd.n10496 92.5
R30876 vdd.n12562 vdd.n12561 92.5
R30877 vdd.n12561 vdd.n12560 92.5
R30878 vdd.n10499 vdd.n10498 92.5
R30879 vdd.n12559 vdd.n10499 92.5
R30880 vdd.n12557 vdd.n12556 92.5
R30881 vdd.n12558 vdd.n12557 92.5
R30882 vdd.n12555 vdd.n10502 92.5
R30883 vdd.n10502 vdd.n10501 92.5
R30884 vdd.n12554 vdd.n12553 92.5
R30885 vdd.n12553 vdd.n12552 92.5
R30886 vdd.n10504 vdd.n10503 92.5
R30887 vdd.n12551 vdd.n10504 92.5
R30888 vdd.n12549 vdd.n12548 92.5
R30889 vdd.n12550 vdd.n12549 92.5
R30890 vdd.n12547 vdd.n10506 92.5
R30891 vdd.n10506 vdd.n10505 92.5
R30892 vdd.n12546 vdd.n12545 92.5
R30893 vdd.n12545 vdd.n12544 92.5
R30894 vdd.n10508 vdd.n10507 92.5
R30895 vdd.n12543 vdd.n10508 92.5
R30896 vdd.n12541 vdd.n12540 92.5
R30897 vdd.n12542 vdd.n12541 92.5
R30898 vdd.n12539 vdd.n10509 92.5
R30899 vdd.n10512 vdd.n10509 92.5
R30900 vdd.n12538 vdd.n12537 92.5
R30901 vdd.n12537 vdd.n12536 92.5
R30902 vdd.n10511 vdd.n10510 92.5
R30903 vdd.n12535 vdd.n10511 92.5
R30904 vdd.n12533 vdd.n12532 92.5
R30905 vdd.n12534 vdd.n12533 92.5
R30906 vdd.n12531 vdd.n10514 92.5
R30907 vdd.n10514 vdd.n10513 92.5
R30908 vdd.n12530 vdd.n12529 92.5
R30909 vdd.n12529 vdd.n12528 92.5
R30910 vdd.n10516 vdd.n10515 92.5
R30911 vdd.n10518 vdd.n10516 92.5
R30912 vdd.n12518 vdd.n12517 92.5
R30913 vdd.n12519 vdd.n12518 92.5
R30914 vdd.n12516 vdd.n10525 92.5
R30915 vdd.n10553 vdd.n10525 92.5
R30916 vdd.n12515 vdd.n12514 92.5
R30917 vdd.n12514 vdd.n12513 92.5
R30918 vdd.n10527 vdd.n10526 92.5
R30919 vdd.n12502 vdd.n10527 92.5
R30920 vdd.n10580 vdd.n10578 92.5
R30921 vdd.n10578 vdd.n10577 92.5
R30922 vdd.n12487 vdd.n12486 92.5
R30923 vdd.n12488 vdd.n12487 92.5
R30924 vdd.n12485 vdd.n10579 92.5
R30925 vdd.n10598 vdd.n10579 92.5
R30926 vdd.n12484 vdd.n12483 92.5
R30927 vdd.n12483 vdd.n12482 92.5
R30928 vdd.n10582 vdd.n10581 92.5
R30929 vdd.n12471 vdd.n10582 92.5
R30930 vdd.n10619 vdd.n10617 92.5
R30931 vdd.n10617 vdd.n10614 92.5
R30932 vdd.n12458 vdd.n12457 92.5
R30933 vdd.n12459 vdd.n12458 92.5
R30934 vdd.n12456 vdd.n10618 92.5
R30935 vdd.n10646 vdd.n10618 92.5
R30936 vdd.n12455 vdd.n12454 92.5
R30937 vdd.n12454 vdd.n12453 92.5
R30938 vdd.n10621 vdd.n10620 92.5
R30939 vdd.n12442 vdd.n10621 92.5
R30940 vdd.n10668 vdd.n10666 92.5
R30941 vdd.n10666 vdd.n10665 92.5
R30942 vdd.n12430 vdd.n12429 92.5
R30943 vdd.n12431 vdd.n12430 92.5
R30944 vdd.n12428 vdd.n10667 92.5
R30945 vdd.n10689 vdd.n10667 92.5
R30946 vdd.n12427 vdd.n12426 92.5
R30947 vdd.n12426 vdd.n12425 92.5
R30948 vdd.n10670 vdd.n10669 92.5
R30949 vdd.n12414 vdd.n10670 92.5
R30950 vdd.n10716 vdd.n10714 92.5
R30951 vdd.n10714 vdd.n10713 92.5
R30952 vdd.n12399 vdd.n12398 92.5
R30953 vdd.n12400 vdd.n12399 92.5
R30954 vdd.n12397 vdd.n10715 92.5
R30955 vdd.n10738 vdd.n10715 92.5
R30956 vdd.n12396 vdd.n12395 92.5
R30957 vdd.n12395 vdd.n12394 92.5
R30958 vdd.n10718 vdd.n10717 92.5
R30959 vdd.n12383 vdd.n10718 92.5
R30960 vdd.n10769 vdd.n10768 92.5
R30961 vdd.n10768 vdd.n10749 92.5
R30962 vdd.n10770 vdd.n10766 92.5
R30963 vdd.n10766 vdd.n10763 92.5
R30964 vdd.n12369 vdd.n12368 92.5
R30965 vdd.n12370 vdd.n12369 92.5
R30966 vdd.n12367 vdd.n10767 92.5
R30967 vdd.n10797 vdd.n10767 92.5
R30968 vdd.n12366 vdd.n12365 92.5
R30969 vdd.n12365 vdd.n12364 92.5
R30970 vdd.n10772 vdd.n10771 92.5
R30971 vdd.n12353 vdd.n10772 92.5
R30972 vdd.n10821 vdd.n10819 92.5
R30973 vdd.n10819 vdd.n10816 92.5
R30974 vdd.n12340 vdd.n12339 92.5
R30975 vdd.n12341 vdd.n12340 92.5
R30976 vdd.n12338 vdd.n10820 92.5
R30977 vdd.n10845 vdd.n10820 92.5
R30978 vdd.n12337 vdd.n12336 92.5
R30979 vdd.n12336 vdd.n12335 92.5
R30980 vdd.n10823 vdd.n10822 92.5
R30981 vdd.n10860 vdd.n10823 92.5
R30982 vdd.n12322 vdd.n12321 92.5
R30983 vdd.n12323 vdd.n12322 92.5
R30984 vdd.n12320 vdd.n10863 92.5
R30985 vdd.n10885 vdd.n10863 92.5
R30986 vdd.n12319 vdd.n12318 92.5
R30987 vdd.n12318 vdd.n12317 92.5
R30988 vdd.n10865 vdd.n10864 92.5
R30989 vdd.n12306 vdd.n10865 92.5
R30990 vdd.n10912 vdd.n10910 92.5
R30991 vdd.n10910 vdd.n10909 92.5
R30992 vdd.n12291 vdd.n12290 92.5
R30993 vdd.n12292 vdd.n12291 92.5
R30994 vdd.n12289 vdd.n10911 92.5
R30995 vdd.n10938 vdd.n10911 92.5
R30996 vdd.n12288 vdd.n12287 92.5
R30997 vdd.n12287 vdd.n12286 92.5
R30998 vdd.n10914 vdd.n10913 92.5
R30999 vdd.n12279 vdd.n10914 92.5
R31000 vdd.n10956 vdd.n10954 92.5
R31001 vdd.n10954 vdd.n10922 92.5
R31002 vdd.n12268 vdd.n12267 92.5
R31003 vdd.n12269 vdd.n12268 92.5
R31004 vdd.n12266 vdd.n10955 92.5
R31005 vdd.n10984 vdd.n10955 92.5
R31006 vdd.n12265 vdd.n12264 92.5
R31007 vdd.n12264 vdd.n12263 92.5
R31008 vdd.n10958 vdd.n10957 92.5
R31009 vdd.n12252 vdd.n10958 92.5
R31010 vdd.n11008 vdd.n11006 92.5
R31011 vdd.n11006 vdd.n11003 92.5
R31012 vdd.n12239 vdd.n12238 92.5
R31013 vdd.n12240 vdd.n12239 92.5
R31014 vdd.n12237 vdd.n11007 92.5
R31015 vdd.n11028 vdd.n11007 92.5
R31016 vdd.n12236 vdd.n12235 92.5
R31017 vdd.n12235 vdd.n12234 92.5
R31018 vdd.n11010 vdd.n11009 92.5
R31019 vdd.n12223 vdd.n11010 92.5
R31020 vdd.n11053 vdd.n11051 92.5
R31021 vdd.n11051 vdd.n11050 92.5
R31022 vdd.n12208 vdd.n12207 92.5
R31023 vdd.n12209 vdd.n12208 92.5
R31024 vdd.n12206 vdd.n11052 92.5
R31025 vdd.n11075 vdd.n11052 92.5
R31026 vdd.n12205 vdd.n12204 92.5
R31027 vdd.n12204 vdd.n12203 92.5
R31028 vdd.n11055 vdd.n11054 92.5
R31029 vdd.n12192 vdd.n11055 92.5
R31030 vdd.n11102 vdd.n11100 92.5
R31031 vdd.n11100 vdd.n11099 92.5
R31032 vdd.n12178 vdd.n12177 92.5
R31033 vdd.n12179 vdd.n12178 92.5
R31034 vdd.n12176 vdd.n11101 92.5
R31035 vdd.n11118 vdd.n11101 92.5
R31036 vdd.n12175 vdd.n12174 92.5
R31037 vdd.n12174 vdd.n12173 92.5
R31038 vdd.n11104 vdd.n11103 92.5
R31039 vdd.n12162 vdd.n11104 92.5
R31040 vdd.n11142 vdd.n11140 92.5
R31041 vdd.n11140 vdd.n11137 92.5
R31042 vdd.n12149 vdd.n12148 92.5
R31043 vdd.n12150 vdd.n12149 92.5
R31044 vdd.n12147 vdd.n11141 92.5
R31045 vdd.n11169 vdd.n11141 92.5
R31046 vdd.n12146 vdd.n12145 92.5
R31047 vdd.n12145 vdd.n12144 92.5
R31048 vdd.n11144 vdd.n11143 92.5
R31049 vdd.n12133 vdd.n11144 92.5
R31050 vdd.n11188 vdd.n11186 92.5
R31051 vdd.n11186 vdd.n11184 92.5
R31052 vdd.n12120 vdd.n12119 92.5
R31053 vdd.n12121 vdd.n12120 92.5
R31054 vdd.n12118 vdd.n11187 92.5
R31055 vdd.n11210 vdd.n11187 92.5
R31056 vdd.n12117 vdd.n12116 92.5
R31057 vdd.n12116 vdd.n12115 92.5
R31058 vdd.n11190 vdd.n11189 92.5
R31059 vdd.n12104 vdd.n11190 92.5
R31060 vdd.n11237 vdd.n11235 92.5
R31061 vdd.n11235 vdd.n11234 92.5
R31062 vdd.n12089 vdd.n12088 92.5
R31063 vdd.n12090 vdd.n12089 92.5
R31064 vdd.n12087 vdd.n11236 92.5
R31065 vdd.n11259 vdd.n11236 92.5
R31066 vdd.n12086 vdd.n12085 92.5
R31067 vdd.n12085 vdd.n12084 92.5
R31068 vdd.n11239 vdd.n11238 92.5
R31069 vdd.n12074 vdd.n11239 92.5
R31070 vdd.n11278 vdd.n11276 92.5
R31071 vdd.n11276 vdd.n11273 92.5
R31072 vdd.n12063 vdd.n12062 92.5
R31073 vdd.n12064 vdd.n12063 92.5
R31074 vdd.n12061 vdd.n11277 92.5
R31075 vdd.n11306 vdd.n11277 92.5
R31076 vdd.n12060 vdd.n12059 92.5
R31077 vdd.n12059 vdd.n12058 92.5
R31078 vdd.n11280 vdd.n11279 92.5
R31079 vdd.n12047 vdd.n11280 92.5
R31080 vdd.n11330 vdd.n11328 92.5
R31081 vdd.n11328 vdd.n11325 92.5
R31082 vdd.n12034 vdd.n12033 92.5
R31083 vdd.n12035 vdd.n12034 92.5
R31084 vdd.n12032 vdd.n11329 92.5
R31085 vdd.n11354 vdd.n11329 92.5
R31086 vdd.n12031 vdd.n12030 92.5
R31087 vdd.n12030 vdd.n12029 92.5
R31088 vdd.n11332 vdd.n11331 92.5
R31089 vdd.n11369 vdd.n11332 92.5
R31090 vdd.n12016 vdd.n12015 92.5
R31091 vdd.n12017 vdd.n12016 92.5
R31092 vdd.n12014 vdd.n11372 92.5
R31093 vdd.n11394 vdd.n11372 92.5
R31094 vdd.n12013 vdd.n12012 92.5
R31095 vdd.n12012 vdd.n12011 92.5
R31096 vdd.n11374 vdd.n11373 92.5
R31097 vdd.n12000 vdd.n11374 92.5
R31098 vdd.n11421 vdd.n11419 92.5
R31099 vdd.n11419 vdd.n11418 92.5
R31100 vdd.n11985 vdd.n11984 92.5
R31101 vdd.n11986 vdd.n11985 92.5
R31102 vdd.n11983 vdd.n11420 92.5
R31103 vdd.n11482 vdd.n11420 92.5
R31104 vdd.n11982 vdd.n11981 92.5
R31105 vdd.n11981 vdd.n11980 92.5
R31106 vdd.n11423 vdd.n11422 92.5
R31107 vdd.n11973 vdd.n11423 92.5
R31108 vdd.n11441 vdd.n11439 92.5
R31109 vdd.n11439 vdd.n11431 92.5
R31110 vdd.n11962 vdd.n11961 92.5
R31111 vdd.n11963 vdd.n11962 92.5
R31112 vdd.n11960 vdd.n11440 92.5
R31113 vdd.n11528 vdd.n11440 92.5
R31114 vdd.n11959 vdd.n11958 92.5
R31115 vdd.n11958 vdd.n11957 92.5
R31116 vdd.n11443 vdd.n11442 92.5
R31117 vdd.n11945 vdd.n11443 92.5
R31118 vdd.n11932 vdd.n11931 92.5
R31119 vdd.n11933 vdd.n11932 92.5
R31120 vdd.n11930 vdd.n11561 92.5
R31121 vdd.n11599 vdd.n11561 92.5
R31122 vdd.n11929 vdd.n11928 92.5
R31123 vdd.n11928 vdd.n11927 92.5
R31124 vdd.n11563 vdd.n11562 92.5
R31125 vdd.n11926 vdd.n11563 92.5
R31126 vdd.n11924 vdd.n11923 92.5
R31127 vdd.n11925 vdd.n11924 92.5
R31128 vdd.n24085 vdd.n24084 92.5
R31129 vdd.n24084 vdd.n24083 92.5
R31130 vdd.n24088 vdd.n24087 92.5
R31131 vdd.n24087 vdd.n24086 92.5
R31132 vdd.n23853 vdd.n23852 92.5
R31133 vdd.n23852 vdd.n23851 92.5
R31134 vdd.n23856 vdd.n23855 92.5
R31135 vdd.n23855 vdd.n23854 92.5
R31136 vdd.n23165 vdd.n23164 92.5
R31137 vdd.n23164 vdd.n23163 92.5
R31138 vdd.n23168 vdd.n23167 92.5
R31139 vdd.n23167 vdd.n23166 92.5
R31140 vdd.n23397 vdd.n23396 92.5
R31141 vdd.n23396 vdd.n23395 92.5
R31142 vdd.n23400 vdd.n23399 92.5
R31143 vdd.n23399 vdd.n23398 92.5
R31144 vdd.n22586 vdd.n22585 92.5
R31145 vdd.n22585 vdd.n22584 92.5
R31146 vdd.n22589 vdd.n22588 92.5
R31147 vdd.n22588 vdd.n22587 92.5
R31148 vdd.n22818 vdd.n22817 92.5
R31149 vdd.n22817 vdd.n22816 92.5
R31150 vdd.n22821 vdd.n22820 92.5
R31151 vdd.n22820 vdd.n22819 92.5
R31152 vdd.n23048 vdd.n23047 92.5
R31153 vdd.n23047 vdd.n23046 92.5
R31154 vdd.n22372 vdd.n22371 92.5
R31155 vdd.n22371 vdd.n22370 92.5
R31156 vdd.n22369 vdd.n22368 92.5
R31157 vdd.n22368 vdd.n22367 92.5
R31158 vdd.n24317 vdd.n24316 92.5
R31159 vdd.n24316 vdd.n24315 92.5
R31160 vdd.n24314 vdd.n24313 92.5
R31161 vdd.n24313 vdd.n24312 92.5
R31162 vdd.n16700 vdd.n16699 92.5
R31163 vdd.n16728 vdd.n16727 92.5
R31164 vdd.n16715 vdd.n16714 92.5
R31165 vdd.n16750 vdd.n16749 92.5
R31166 vdd.n16760 vdd.n16759 92.5
R31167 vdd.n15454 vdd.n15453 92.5
R31168 vdd.n15455 vdd.n15454 92.5
R31169 vdd.n15459 vdd.n15458 92.5
R31170 vdd.n15460 vdd.n15459 92.5
R31171 vdd.n15476 vdd.n15475 92.5
R31172 vdd.n15477 vdd.n15476 92.5
R31173 vdd.n15493 vdd.n15492 92.5
R31174 vdd.n15494 vdd.n15493 92.5
R31175 vdd.n15510 vdd.n15509 92.5
R31176 vdd.n15511 vdd.n15510 92.5
R31177 vdd.n15529 vdd.n15528 92.5
R31178 vdd.n15530 vdd.n15529 92.5
R31179 vdd.n15550 vdd.n15549 92.5
R31180 vdd.n15554 vdd.n15553 92.5
R31181 vdd.n15555 vdd.n15554 92.5
R31182 vdd.n15571 vdd.n15570 92.5
R31183 vdd.n15572 vdd.n15571 92.5
R31184 vdd.n15588 vdd.n15587 92.5
R31185 vdd.n15589 vdd.n15588 92.5
R31186 vdd.n15605 vdd.n15604 92.5
R31187 vdd.n15606 vdd.n15605 92.5
R31188 vdd.n15622 vdd.n15621 92.5
R31189 vdd.n15623 vdd.n15622 92.5
R31190 vdd.n15639 vdd.n15638 92.5
R31191 vdd.n15640 vdd.n15639 92.5
R31192 vdd.n15656 vdd.n15655 92.5
R31193 vdd.n15657 vdd.n15656 92.5
R31194 vdd.n15226 vdd.n15225 92.5
R31195 vdd.n15227 vdd.n15226 92.5
R31196 vdd.n15212 vdd.n15211 92.5
R31197 vdd.n15213 vdd.n15212 92.5
R31198 vdd.n15676 vdd.n15675 92.5
R31199 vdd.n15677 vdd.n15676 92.5
R31200 vdd.n15693 vdd.n15692 92.5
R31201 vdd.n15694 vdd.n15693 92.5
R31202 vdd.n15710 vdd.n15709 92.5
R31203 vdd.n15711 vdd.n15710 92.5
R31204 vdd.n15715 vdd.n15714 92.5
R31205 vdd.n15716 vdd.n15715 92.5
R31206 vdd.n15732 vdd.n15731 92.5
R31207 vdd.n15733 vdd.n15732 92.5
R31208 vdd.n15749 vdd.n15748 92.5
R31209 vdd.n15750 vdd.n15749 92.5
R31210 vdd.n15766 vdd.n15765 92.5
R31211 vdd.n15767 vdd.n15766 92.5
R31212 vdd.n15785 vdd.n15784 92.5
R31213 vdd.n15786 vdd.n15785 92.5
R31214 vdd.n15806 vdd.n15805 92.5
R31215 vdd.n15810 vdd.n15809 92.5
R31216 vdd.n15811 vdd.n15810 92.5
R31217 vdd.n15827 vdd.n15826 92.5
R31218 vdd.n15828 vdd.n15827 92.5
R31219 vdd.n15844 vdd.n15843 92.5
R31220 vdd.n15845 vdd.n15844 92.5
R31221 vdd.n15861 vdd.n15860 92.5
R31222 vdd.n15862 vdd.n15861 92.5
R31223 vdd.n15878 vdd.n15877 92.5
R31224 vdd.n15879 vdd.n15878 92.5
R31225 vdd.n15895 vdd.n15894 92.5
R31226 vdd.n15896 vdd.n15895 92.5
R31227 vdd.n15912 vdd.n15911 92.5
R31228 vdd.n15913 vdd.n15912 92.5
R31229 vdd.n15186 vdd.n15185 92.5
R31230 vdd.n15187 vdd.n15186 92.5
R31231 vdd.n15198 vdd.n15197 92.5
R31232 vdd.n15199 vdd.n15198 92.5
R31233 vdd.n15932 vdd.n15931 92.5
R31234 vdd.n15933 vdd.n15932 92.5
R31235 vdd.n15949 vdd.n15948 92.5
R31236 vdd.n15950 vdd.n15949 92.5
R31237 vdd.n15966 vdd.n15965 92.5
R31238 vdd.n15967 vdd.n15966 92.5
R31239 vdd.n15971 vdd.n15970 92.5
R31240 vdd.n15972 vdd.n15971 92.5
R31241 vdd.n15988 vdd.n15987 92.5
R31242 vdd.n15989 vdd.n15988 92.5
R31243 vdd.n16005 vdd.n16004 92.5
R31244 vdd.n16006 vdd.n16005 92.5
R31245 vdd.n16022 vdd.n16021 92.5
R31246 vdd.n16023 vdd.n16022 92.5
R31247 vdd.n16041 vdd.n16040 92.5
R31248 vdd.n16042 vdd.n16041 92.5
R31249 vdd.n16062 vdd.n16061 92.5
R31250 vdd.n16066 vdd.n16065 92.5
R31251 vdd.n16067 vdd.n16066 92.5
R31252 vdd.n16083 vdd.n16082 92.5
R31253 vdd.n16084 vdd.n16083 92.5
R31254 vdd.n16100 vdd.n16099 92.5
R31255 vdd.n16101 vdd.n16100 92.5
R31256 vdd.n16117 vdd.n16116 92.5
R31257 vdd.n16118 vdd.n16117 92.5
R31258 vdd.n16134 vdd.n16133 92.5
R31259 vdd.n16135 vdd.n16134 92.5
R31260 vdd.n16151 vdd.n16150 92.5
R31261 vdd.n16152 vdd.n16151 92.5
R31262 vdd.n16168 vdd.n16167 92.5
R31263 vdd.n16169 vdd.n16168 92.5
R31264 vdd.n15170 vdd.n15169 92.5
R31265 vdd.n15171 vdd.n15170 92.5
R31266 vdd.n15156 vdd.n15155 92.5
R31267 vdd.n15157 vdd.n15156 92.5
R31268 vdd.n16188 vdd.n16187 92.5
R31269 vdd.n16189 vdd.n16188 92.5
R31270 vdd.n16205 vdd.n16204 92.5
R31271 vdd.n16206 vdd.n16205 92.5
R31272 vdd.n16222 vdd.n16221 92.5
R31273 vdd.n16223 vdd.n16222 92.5
R31274 vdd.n16227 vdd.n16226 92.5
R31275 vdd.n16228 vdd.n16227 92.5
R31276 vdd.n16244 vdd.n16243 92.5
R31277 vdd.n16245 vdd.n16244 92.5
R31278 vdd.n16261 vdd.n16260 92.5
R31279 vdd.n16262 vdd.n16261 92.5
R31280 vdd.n16278 vdd.n16277 92.5
R31281 vdd.n16279 vdd.n16278 92.5
R31282 vdd.n16297 vdd.n16296 92.5
R31283 vdd.n16298 vdd.n16297 92.5
R31284 vdd.n16318 vdd.n16317 92.5
R31285 vdd.n16322 vdd.n16321 92.5
R31286 vdd.n16323 vdd.n16322 92.5
R31287 vdd.n16339 vdd.n16338 92.5
R31288 vdd.n16340 vdd.n16339 92.5
R31289 vdd.n16356 vdd.n16355 92.5
R31290 vdd.n16357 vdd.n16356 92.5
R31291 vdd.n16373 vdd.n16372 92.5
R31292 vdd.n16374 vdd.n16373 92.5
R31293 vdd.n16390 vdd.n16389 92.5
R31294 vdd.n16391 vdd.n16390 92.5
R31295 vdd.n16407 vdd.n16406 92.5
R31296 vdd.n16408 vdd.n16407 92.5
R31297 vdd.n16424 vdd.n16423 92.5
R31298 vdd.n16425 vdd.n16424 92.5
R31299 vdd.n15142 vdd.n15141 92.5
R31300 vdd.n15143 vdd.n15142 92.5
R31301 vdd.n15128 vdd.n15127 92.5
R31302 vdd.n15129 vdd.n15128 92.5
R31303 vdd.n16444 vdd.n16443 92.5
R31304 vdd.n16445 vdd.n16444 92.5
R31305 vdd.n16461 vdd.n16460 92.5
R31306 vdd.n16462 vdd.n16461 92.5
R31307 vdd.n16478 vdd.n16477 92.5
R31308 vdd.n16479 vdd.n16478 92.5
R31309 vdd.n16483 vdd.n16482 92.5
R31310 vdd.n16484 vdd.n16483 92.5
R31311 vdd.n16500 vdd.n16499 92.5
R31312 vdd.n16501 vdd.n16500 92.5
R31313 vdd.n16517 vdd.n16516 92.5
R31314 vdd.n16518 vdd.n16517 92.5
R31315 vdd.n16534 vdd.n16533 92.5
R31316 vdd.n16535 vdd.n16534 92.5
R31317 vdd.n16569 vdd.n16568 92.5
R31318 vdd.n16570 vdd.n16569 92.5
R31319 vdd.n16563 vdd.n16562 92.5
R31320 vdd.n16560 vdd.n16559 92.5
R31321 vdd.n16554 vdd.n16553 92.5
R31322 vdd.n16609 vdd.n16608 92.5
R31323 vdd.n16614 vdd.n16613 92.5
R31324 vdd.n16620 vdd.n16619 92.5
R31325 vdd.n16628 vdd.n16627 92.5
R31326 vdd.n16639 vdd.n16638 92.5
R31327 vdd.n16640 vdd.n16639 92.5
R31328 vdd.n16651 vdd.n16650 92.5
R31329 vdd.n16652 vdd.n16651 92.5
R31330 vdd.n16660 vdd.n16659 92.5
R31331 vdd.n16661 vdd.n16660 92.5
R31332 vdd.n15073 vdd.n15072 92.5
R31333 vdd.n15082 vdd.n15081 92.5
R31334 vdd.n15083 vdd.n15082 92.5
R31335 vdd.n15114 vdd.n15113 92.5
R31336 vdd.n15115 vdd.n15114 92.5
R31337 vdd.n15103 vdd.n15102 92.5
R31338 vdd.n15101 vdd.n15100 92.5
R31339 vdd.n15099 vdd.n15098 92.5
R31340 vdd.n15097 vdd.n15096 92.5
R31341 vdd.n15095 vdd.n15094 92.5
R31342 vdd.n15093 vdd.n15092 92.5
R31343 vdd.n15091 vdd.n15090 92.5
R31344 vdd.n15089 vdd.n15088 92.5
R31345 vdd.n15087 vdd.n15086 92.5
R31346 vdd.n16839 vdd.n16838 92.5
R31347 vdd.n16841 vdd.n16840 92.5
R31348 vdd.n16843 vdd.n16842 92.5
R31349 vdd.n16845 vdd.n16844 92.5
R31350 vdd.n16847 vdd.n16846 92.5
R31351 vdd.n16849 vdd.n16848 92.5
R31352 vdd.n16851 vdd.n16850 92.5
R31353 vdd.n16853 vdd.n16852 92.5
R31354 vdd.n16863 vdd.n16862 92.5
R31355 vdd.n16864 vdd.n16863 92.5
R31356 vdd.n16867 vdd.n16866 92.5
R31357 vdd.n16868 vdd.n16867 92.5
R31358 vdd.n16881 vdd.n16880 92.5
R31359 vdd.n16882 vdd.n16881 92.5
R31360 vdd.n16897 vdd.n16896 92.5
R31361 vdd.n16898 vdd.n16897 92.5
R31362 vdd.n16913 vdd.n16912 92.5
R31363 vdd.n16914 vdd.n16913 92.5
R31364 vdd.n16929 vdd.n16928 92.5
R31365 vdd.n16930 vdd.n16929 92.5
R31366 vdd.n16945 vdd.n16944 92.5
R31367 vdd.n16946 vdd.n16945 92.5
R31368 vdd.n16961 vdd.n16960 92.5
R31369 vdd.n16962 vdd.n16961 92.5
R31370 vdd.n16975 vdd.n16974 92.5
R31371 vdd.n16976 vdd.n16975 92.5
R31372 vdd.n16989 vdd.n16988 92.5
R31373 vdd.n16990 vdd.n16989 92.5
R31374 vdd.n17005 vdd.n17004 92.5
R31375 vdd.n17006 vdd.n17005 92.5
R31376 vdd.n17021 vdd.n17020 92.5
R31377 vdd.n17022 vdd.n17021 92.5
R31378 vdd.n17037 vdd.n17036 92.5
R31379 vdd.n17038 vdd.n17037 92.5
R31380 vdd.n17053 vdd.n17052 92.5
R31381 vdd.n17054 vdd.n17053 92.5
R31382 vdd.n17069 vdd.n17068 92.5
R31383 vdd.n17070 vdd.n17069 92.5
R31384 vdd.n17085 vdd.n17084 92.5
R31385 vdd.n17086 vdd.n17085 92.5
R31386 vdd.n17101 vdd.n17100 92.5
R31387 vdd.n17102 vdd.n17101 92.5
R31388 vdd.n17117 vdd.n17116 92.5
R31389 vdd.n17118 vdd.n17117 92.5
R31390 vdd.n17121 vdd.n17120 92.5
R31391 vdd.n17122 vdd.n17121 92.5
R31392 vdd.n17137 vdd.n17136 92.5
R31393 vdd.n17138 vdd.n17137 92.5
R31394 vdd.n17153 vdd.n17152 92.5
R31395 vdd.n17154 vdd.n17153 92.5
R31396 vdd.n17169 vdd.n17168 92.5
R31397 vdd.n17170 vdd.n17169 92.5
R31398 vdd.n17185 vdd.n17184 92.5
R31399 vdd.n17186 vdd.n17185 92.5
R31400 vdd.n17201 vdd.n17200 92.5
R31401 vdd.n17202 vdd.n17201 92.5
R31402 vdd.n17217 vdd.n17216 92.5
R31403 vdd.n17218 vdd.n17217 92.5
R31404 vdd.n17233 vdd.n17232 92.5
R31405 vdd.n17234 vdd.n17233 92.5
R31406 vdd.n17247 vdd.n17246 92.5
R31407 vdd.n17248 vdd.n17247 92.5
R31408 vdd.n17261 vdd.n17260 92.5
R31409 vdd.n17262 vdd.n17261 92.5
R31410 vdd.n17277 vdd.n17276 92.5
R31411 vdd.n17278 vdd.n17277 92.5
R31412 vdd.n17293 vdd.n17292 92.5
R31413 vdd.n17294 vdd.n17293 92.5
R31414 vdd.n17309 vdd.n17308 92.5
R31415 vdd.n17310 vdd.n17309 92.5
R31416 vdd.n17325 vdd.n17324 92.5
R31417 vdd.n17326 vdd.n17325 92.5
R31418 vdd.n17341 vdd.n17340 92.5
R31419 vdd.n17342 vdd.n17341 92.5
R31420 vdd.n17357 vdd.n17356 92.5
R31421 vdd.n17358 vdd.n17357 92.5
R31422 vdd.n17373 vdd.n17372 92.5
R31423 vdd.n17374 vdd.n17373 92.5
R31424 vdd.n17389 vdd.n17388 92.5
R31425 vdd.n17390 vdd.n17389 92.5
R31426 vdd.n17393 vdd.n17392 92.5
R31427 vdd.n17394 vdd.n17393 92.5
R31428 vdd.n17409 vdd.n17408 92.5
R31429 vdd.n17410 vdd.n17409 92.5
R31430 vdd.n17425 vdd.n17424 92.5
R31431 vdd.n17426 vdd.n17425 92.5
R31432 vdd.n17441 vdd.n17440 92.5
R31433 vdd.n17442 vdd.n17441 92.5
R31434 vdd.n17457 vdd.n17456 92.5
R31435 vdd.n17458 vdd.n17457 92.5
R31436 vdd.n17473 vdd.n17472 92.5
R31437 vdd.n17474 vdd.n17473 92.5
R31438 vdd.n17489 vdd.n17488 92.5
R31439 vdd.n17490 vdd.n17489 92.5
R31440 vdd.n17505 vdd.n17504 92.5
R31441 vdd.n17506 vdd.n17505 92.5
R31442 vdd.n17519 vdd.n17518 92.5
R31443 vdd.n17520 vdd.n17519 92.5
R31444 vdd.n17533 vdd.n17532 92.5
R31445 vdd.n17534 vdd.n17533 92.5
R31446 vdd.n17549 vdd.n17548 92.5
R31447 vdd.n17550 vdd.n17549 92.5
R31448 vdd.n17565 vdd.n17564 92.5
R31449 vdd.n17566 vdd.n17565 92.5
R31450 vdd.n17581 vdd.n17580 92.5
R31451 vdd.n17582 vdd.n17581 92.5
R31452 vdd.n16826 vdd.n16825 92.5
R31453 vdd.n16827 vdd.n16826 92.5
R31454 vdd.n17599 vdd.n17598 92.5
R31455 vdd.n17600 vdd.n17599 92.5
R31456 vdd.n17615 vdd.n17614 92.5
R31457 vdd.n17616 vdd.n17615 92.5
R31458 vdd.n17631 vdd.n17630 92.5
R31459 vdd.n17632 vdd.n17631 92.5
R31460 vdd.n17647 vdd.n17646 92.5
R31461 vdd.n17648 vdd.n17647 92.5
R31462 vdd.n17651 vdd.n17650 92.5
R31463 vdd.n17652 vdd.n17651 92.5
R31464 vdd.n17667 vdd.n17666 92.5
R31465 vdd.n17668 vdd.n17667 92.5
R31466 vdd.n17683 vdd.n17682 92.5
R31467 vdd.n17684 vdd.n17683 92.5
R31468 vdd.n17699 vdd.n17698 92.5
R31469 vdd.n17700 vdd.n17699 92.5
R31470 vdd.n17715 vdd.n17714 92.5
R31471 vdd.n17716 vdd.n17715 92.5
R31472 vdd.n17731 vdd.n17730 92.5
R31473 vdd.n17732 vdd.n17731 92.5
R31474 vdd.n17747 vdd.n17746 92.5
R31475 vdd.n17748 vdd.n17747 92.5
R31476 vdd.n17763 vdd.n17762 92.5
R31477 vdd.n17764 vdd.n17763 92.5
R31478 vdd.n17777 vdd.n17776 92.5
R31479 vdd.n17778 vdd.n17777 92.5
R31480 vdd.n17791 vdd.n17790 92.5
R31481 vdd.n17792 vdd.n17791 92.5
R31482 vdd.n17807 vdd.n17806 92.5
R31483 vdd.n17808 vdd.n17807 92.5
R31484 vdd.n17823 vdd.n17822 92.5
R31485 vdd.n17824 vdd.n17823 92.5
R31486 vdd.n17839 vdd.n17838 92.5
R31487 vdd.n17840 vdd.n17839 92.5
R31488 vdd.n17855 vdd.n17854 92.5
R31489 vdd.n17856 vdd.n17855 92.5
R31490 vdd.n17871 vdd.n17870 92.5
R31491 vdd.n17872 vdd.n17871 92.5
R31492 vdd.n17886 vdd.n17885 92.5
R31493 vdd.n17887 vdd.n17886 92.5
R31494 vdd.n17902 vdd.n17901 92.5
R31495 vdd.n17903 vdd.n17902 92.5
R31496 vdd.n17918 vdd.n17917 92.5
R31497 vdd.n17919 vdd.n17918 92.5
R31498 vdd.n17922 vdd.n17921 92.5
R31499 vdd.n17923 vdd.n17922 92.5
R31500 vdd.n17938 vdd.n17937 92.5
R31501 vdd.n17939 vdd.n17938 92.5
R31502 vdd.n17954 vdd.n17953 92.5
R31503 vdd.n17955 vdd.n17954 92.5
R31504 vdd.n17970 vdd.n17969 92.5
R31505 vdd.n17971 vdd.n17970 92.5
R31506 vdd.n17986 vdd.n17985 92.5
R31507 vdd.n17987 vdd.n17986 92.5
R31508 vdd.n18002 vdd.n18001 92.5
R31509 vdd.n18003 vdd.n18002 92.5
R31510 vdd.n18018 vdd.n18017 92.5
R31511 vdd.n18019 vdd.n18018 92.5
R31512 vdd.n18034 vdd.n18033 92.5
R31513 vdd.n18035 vdd.n18034 92.5
R31514 vdd.n18048 vdd.n18047 92.5
R31515 vdd.n18049 vdd.n18048 92.5
R31516 vdd.n18062 vdd.n18061 92.5
R31517 vdd.n18063 vdd.n18062 92.5
R31518 vdd.n18078 vdd.n18077 92.5
R31519 vdd.n18079 vdd.n18078 92.5
R31520 vdd.n18094 vdd.n18093 92.5
R31521 vdd.n18095 vdd.n18094 92.5
R31522 vdd.n18110 vdd.n18109 92.5
R31523 vdd.n18111 vdd.n18110 92.5
R31524 vdd.n18126 vdd.n18125 92.5
R31525 vdd.n18127 vdd.n18126 92.5
R31526 vdd.n18142 vdd.n18141 92.5
R31527 vdd.n18143 vdd.n18142 92.5
R31528 vdd.n18158 vdd.n18157 92.5
R31529 vdd.n18159 vdd.n18158 92.5
R31530 vdd.n18174 vdd.n18173 92.5
R31531 vdd.n18175 vdd.n18174 92.5
R31532 vdd.n18190 vdd.n18189 92.5
R31533 vdd.n18191 vdd.n18190 92.5
R31534 vdd.n18194 vdd.n18193 92.5
R31535 vdd.n18195 vdd.n18194 92.5
R31536 vdd.n18210 vdd.n18209 92.5
R31537 vdd.n18211 vdd.n18210 92.5
R31538 vdd.n18226 vdd.n18225 92.5
R31539 vdd.n18241 vdd.n18240 92.5
R31540 vdd.n18256 vdd.n18255 92.5
R31541 vdd.n18271 vdd.n18270 92.5
R31542 vdd.n18286 vdd.n18285 92.5
R31543 vdd.n18301 vdd.n18300 92.5
R31544 vdd.n16815 vdd.n16814 92.5
R31545 vdd.n15033 vdd.n15032 92.5
R31546 vdd.n18326 vdd.n18325 92.5
R31547 vdd.n18343 vdd.n18342 92.5
R31548 vdd.n14988 vdd.n14987 92.5
R31549 vdd.n14990 vdd.n14989 92.5
R31550 vdd.n14992 vdd.n14991 92.5
R31551 vdd.n14994 vdd.n14993 92.5
R31552 vdd.n14996 vdd.n14995 92.5
R31553 vdd.n14998 vdd.n14997 92.5
R31554 vdd.n15000 vdd.n14999 92.5
R31555 vdd.n18496 vdd.n18495 92.5
R31556 vdd.n18510 vdd.n18509 92.5
R31557 vdd.n18529 vdd.n18528 92.5
R31558 vdd.n18545 vdd.n18544 92.5
R31559 vdd.n18561 vdd.n18560 92.5
R31560 vdd.n18577 vdd.n18576 92.5
R31561 vdd.n18593 vdd.n18592 92.5
R31562 vdd.n18609 vdd.n18608 92.5
R31563 vdd.n18625 vdd.n18624 92.5
R31564 vdd.n18643 vdd.n18642 92.5
R31565 vdd.n18659 vdd.n18658 92.5
R31566 vdd.n18675 vdd.n18674 92.5
R31567 vdd.n18691 vdd.n18690 92.5
R31568 vdd.n18707 vdd.n18706 92.5
R31569 vdd.n18723 vdd.n18722 92.5
R31570 vdd.n18739 vdd.n18738 92.5
R31571 vdd.n18755 vdd.n18754 92.5
R31572 vdd.n18769 vdd.n18768 92.5
R31573 vdd.n18788 vdd.n18787 92.5
R31574 vdd.n18804 vdd.n18803 92.5
R31575 vdd.n18820 vdd.n18819 92.5
R31576 vdd.n18836 vdd.n18835 92.5
R31577 vdd.n18852 vdd.n18851 92.5
R31578 vdd.n18868 vdd.n18867 92.5
R31579 vdd.n18884 vdd.n18883 92.5
R31580 vdd.n18902 vdd.n18901 92.5
R31581 vdd.n18918 vdd.n18917 92.5
R31582 vdd.n18934 vdd.n18933 92.5
R31583 vdd.n18950 vdd.n18949 92.5
R31584 vdd.n18966 vdd.n18965 92.5
R31585 vdd.n18982 vdd.n18981 92.5
R31586 vdd.n18998 vdd.n18997 92.5
R31587 vdd.n19014 vdd.n19013 92.5
R31588 vdd.n19028 vdd.n19027 92.5
R31589 vdd.n19047 vdd.n19046 92.5
R31590 vdd.n19063 vdd.n19062 92.5
R31591 vdd.n19079 vdd.n19078 92.5
R31592 vdd.n19095 vdd.n19094 92.5
R31593 vdd.n19111 vdd.n19110 92.5
R31594 vdd.n19126 vdd.n19125 92.5
R31595 vdd.n21003 vdd.n21002 92.5
R31596 vdd.n19151 vdd.n19150 92.5
R31597 vdd.n21025 vdd.n21024 92.5
R31598 vdd.n21041 vdd.n21040 92.5
R31599 vdd.n21057 vdd.n21056 92.5
R31600 vdd.n21073 vdd.n21072 92.5
R31601 vdd.n21085 vdd.n21084 92.5
R31602 vdd.n21105 vdd.n21104 92.5
R31603 vdd.n21121 vdd.n21120 92.5
R31604 vdd.n21135 vdd.n21134 92.5
R31605 vdd.n21154 vdd.n21153 92.5
R31606 vdd.n21170 vdd.n21169 92.5
R31607 vdd.n21186 vdd.n21185 92.5
R31608 vdd.n21202 vdd.n21201 92.5
R31609 vdd.n21218 vdd.n21217 92.5
R31610 vdd.n21234 vdd.n21233 92.5
R31611 vdd.n21250 vdd.n21249 92.5
R31612 vdd.n21268 vdd.n21267 92.5
R31613 vdd.n21284 vdd.n21283 92.5
R31614 vdd.n21300 vdd.n21299 92.5
R31615 vdd.n21316 vdd.n21315 92.5
R31616 vdd.n21332 vdd.n21331 92.5
R31617 vdd.n21348 vdd.n21347 92.5
R31618 vdd.n21364 vdd.n21363 92.5
R31619 vdd.n21380 vdd.n21379 92.5
R31620 vdd.n21394 vdd.n21393 92.5
R31621 vdd.n21413 vdd.n21412 92.5
R31622 vdd.n21429 vdd.n21428 92.5
R31623 vdd.n21445 vdd.n21444 92.5
R31624 vdd.n21461 vdd.n21460 92.5
R31625 vdd.n21477 vdd.n21476 92.5
R31626 vdd.n21493 vdd.n21492 92.5
R31627 vdd.n21509 vdd.n21508 92.5
R31628 vdd.n21527 vdd.n21526 92.5
R31629 vdd.n21543 vdd.n21542 92.5
R31630 vdd.n21559 vdd.n21558 92.5
R31631 vdd.n21575 vdd.n21574 92.5
R31632 vdd.n21591 vdd.n21590 92.5
R31633 vdd.n21615 vdd.n21614 92.5
R31634 vdd.n21609 vdd.n21608 92.5
R31635 vdd.n21672 vdd.n21671 92.5
R31636 vdd.n18477 vdd.n18476 92.5
R31637 vdd.n18479 vdd.n18478 92.5
R31638 vdd.n18472 vdd.n18471 92.5
R31639 vdd.n18474 vdd.n18473 92.5
R31640 vdd.n18467 vdd.n18466 92.5
R31641 vdd.n21667 vdd.n21666 92.5
R31642 vdd.n21668 vdd.n21667 92.5
R31643 vdd.n21671 vdd.n21670 92.5
R31644 vdd.n21614 vdd.n21613 92.5
R31645 vdd.n21590 vdd.n21589 92.5
R31646 vdd.n21574 vdd.n21573 92.5
R31647 vdd.n21558 vdd.n21557 92.5
R31648 vdd.n21542 vdd.n21541 92.5
R31649 vdd.n21526 vdd.n21525 92.5
R31650 vdd.n21515 vdd.n21514 92.5
R31651 vdd.n21516 vdd.n21515 92.5
R31652 vdd.n21508 vdd.n21507 92.5
R31653 vdd.n21492 vdd.n21491 92.5
R31654 vdd.n21476 vdd.n21475 92.5
R31655 vdd.n21460 vdd.n21459 92.5
R31656 vdd.n21444 vdd.n21443 92.5
R31657 vdd.n21428 vdd.n21427 92.5
R31658 vdd.n21412 vdd.n21411 92.5
R31659 vdd.n21393 vdd.n21392 92.5
R31660 vdd.n21396 vdd.n21395 92.5
R31661 vdd.n21397 vdd.n21396 92.5
R31662 vdd.n21379 vdd.n21378 92.5
R31663 vdd.n21363 vdd.n21362 92.5
R31664 vdd.n21347 vdd.n21346 92.5
R31665 vdd.n21331 vdd.n21330 92.5
R31666 vdd.n21315 vdd.n21314 92.5
R31667 vdd.n21299 vdd.n21298 92.5
R31668 vdd.n21283 vdd.n21282 92.5
R31669 vdd.n21267 vdd.n21266 92.5
R31670 vdd.n21256 vdd.n21255 92.5
R31671 vdd.n21257 vdd.n21256 92.5
R31672 vdd.n21249 vdd.n21248 92.5
R31673 vdd.n21233 vdd.n21232 92.5
R31674 vdd.n21217 vdd.n21216 92.5
R31675 vdd.n21201 vdd.n21200 92.5
R31676 vdd.n21185 vdd.n21184 92.5
R31677 vdd.n21169 vdd.n21168 92.5
R31678 vdd.n21153 vdd.n21152 92.5
R31679 vdd.n21134 vdd.n21133 92.5
R31680 vdd.n21137 vdd.n21136 92.5
R31681 vdd.n21138 vdd.n21137 92.5
R31682 vdd.n21120 vdd.n21119 92.5
R31683 vdd.n21104 vdd.n21103 92.5
R31684 vdd.n21084 vdd.n21083 92.5
R31685 vdd.n21072 vdd.n21071 92.5
R31686 vdd.n21056 vdd.n21055 92.5
R31687 vdd.n21040 vdd.n21039 92.5
R31688 vdd.n19150 vdd.n19149 92.5
R31689 vdd.n21008 vdd.n21007 92.5
R31690 vdd.n21009 vdd.n21008 92.5
R31691 vdd.n19110 vdd.n19109 92.5
R31692 vdd.n19094 vdd.n19093 92.5
R31693 vdd.n19078 vdd.n19077 92.5
R31694 vdd.n19062 vdd.n19061 92.5
R31695 vdd.n19046 vdd.n19045 92.5
R31696 vdd.n19027 vdd.n19026 92.5
R31697 vdd.n19030 vdd.n19029 92.5
R31698 vdd.n19031 vdd.n19030 92.5
R31699 vdd.n19013 vdd.n19012 92.5
R31700 vdd.n18997 vdd.n18996 92.5
R31701 vdd.n18981 vdd.n18980 92.5
R31702 vdd.n18965 vdd.n18964 92.5
R31703 vdd.n18949 vdd.n18948 92.5
R31704 vdd.n18933 vdd.n18932 92.5
R31705 vdd.n18917 vdd.n18916 92.5
R31706 vdd.n18901 vdd.n18900 92.5
R31707 vdd.n18890 vdd.n18889 92.5
R31708 vdd.n18891 vdd.n18890 92.5
R31709 vdd.n18883 vdd.n18882 92.5
R31710 vdd.n18867 vdd.n18866 92.5
R31711 vdd.n18851 vdd.n18850 92.5
R31712 vdd.n18835 vdd.n18834 92.5
R31713 vdd.n18819 vdd.n18818 92.5
R31714 vdd.n18803 vdd.n18802 92.5
R31715 vdd.n18787 vdd.n18786 92.5
R31716 vdd.n18768 vdd.n18767 92.5
R31717 vdd.n18771 vdd.n18770 92.5
R31718 vdd.n18772 vdd.n18771 92.5
R31719 vdd.n18754 vdd.n18753 92.5
R31720 vdd.n18738 vdd.n18737 92.5
R31721 vdd.n18722 vdd.n18721 92.5
R31722 vdd.n18706 vdd.n18705 92.5
R31723 vdd.n18690 vdd.n18689 92.5
R31724 vdd.n18674 vdd.n18673 92.5
R31725 vdd.n18658 vdd.n18657 92.5
R31726 vdd.n18642 vdd.n18641 92.5
R31727 vdd.n18631 vdd.n18630 92.5
R31728 vdd.n18632 vdd.n18631 92.5
R31729 vdd.n18624 vdd.n18623 92.5
R31730 vdd.n18608 vdd.n18607 92.5
R31731 vdd.n18592 vdd.n18591 92.5
R31732 vdd.n18576 vdd.n18575 92.5
R31733 vdd.n18560 vdd.n18559 92.5
R31734 vdd.n18544 vdd.n18543 92.5
R31735 vdd.n18528 vdd.n18527 92.5
R31736 vdd.n18509 vdd.n18508 92.5
R31737 vdd.n18512 vdd.n18511 92.5
R31738 vdd.n18513 vdd.n18512 92.5
R31739 vdd.n18495 vdd.n18494 92.5
R31740 vdd.n18469 vdd.n18468 92.5
R31741 vdd.n18460 vdd.n18459 92.5
R31742 vdd.n18449 vdd.n18448 92.5
R31743 vdd.n18445 vdd.n18444 92.5
R31744 vdd.n18441 vdd.n18440 92.5
R31745 vdd.n18437 vdd.n18436 92.5
R31746 vdd.n18433 vdd.n18432 92.5
R31747 vdd.n21634 vdd.n21633 92.5
R31748 vdd.n21728 vdd.n21727 92.5
R31749 vdd.n21726 vdd.n21725 92.5
R31750 vdd.n21723 vdd.n21722 92.5
R31751 vdd.n21721 vdd.n21720 92.5
R31752 vdd.n21718 vdd.n21717 92.5
R31753 vdd.n21716 vdd.n21715 92.5
R31754 vdd.n21713 vdd.n21712 92.5
R31755 vdd.n21711 vdd.n21710 92.5
R31756 vdd.n21660 vdd.n21659 92.5
R31757 vdd.n20543 vdd.n20542 92.5
R31758 vdd.n20559 vdd.n20558 92.5
R31759 vdd.n20575 vdd.n20574 92.5
R31760 vdd.n20591 vdd.n20590 92.5
R31761 vdd.n20607 vdd.n20606 92.5
R31762 vdd.n20623 vdd.n20622 92.5
R31763 vdd.n20637 vdd.n20636 92.5
R31764 vdd.n20656 vdd.n20655 92.5
R31765 vdd.n20672 vdd.n20671 92.5
R31766 vdd.n20688 vdd.n20687 92.5
R31767 vdd.n20704 vdd.n20703 92.5
R31768 vdd.n20719 vdd.n20718 92.5
R31769 vdd.n19944 vdd.n19943 92.5
R31770 vdd.n19932 vdd.n19931 92.5
R31771 vdd.n19920 vdd.n19919 92.5
R31772 vdd.n19908 vdd.n19907 92.5
R31773 vdd.n20749 vdd.n20748 92.5
R31774 vdd.n20765 vdd.n20764 92.5
R31775 vdd.n20780 vdd.n20779 92.5
R31776 vdd.n20796 vdd.n20795 92.5
R31777 vdd.n20812 vdd.n20811 92.5
R31778 vdd.n20825 vdd.n20824 92.5
R31779 vdd.n20839 vdd.n20838 92.5
R31780 vdd.n20855 vdd.n20854 92.5
R31781 vdd.n19889 vdd.n19888 92.5
R31782 vdd.n20876 vdd.n20875 92.5
R31783 vdd.n20892 vdd.n20891 92.5
R31784 vdd.n20908 vdd.n20907 92.5
R31785 vdd.n19876 vdd.n19875 92.5
R31786 vdd.n19864 vdd.n19863 92.5
R31787 vdd.n19852 vdd.n19851 92.5
R31788 vdd.n19839 vdd.n19838 92.5
R31789 vdd.n20939 vdd.n20938 92.5
R31790 vdd.n20955 vdd.n20954 92.5
R31791 vdd.n20971 vdd.n20970 92.5
R31792 vdd.n20987 vdd.n20986 92.5
R31793 vdd.n19156 vdd.n19155 92.5
R31794 vdd.n19169 vdd.n19168 92.5
R31795 vdd.n19819 vdd.n19818 92.5
R31796 vdd.n19806 vdd.n19805 92.5
R31797 vdd.n19790 vdd.n19789 92.5
R31798 vdd.n19774 vdd.n19773 92.5
R31799 vdd.n19758 vdd.n19757 92.5
R31800 vdd.n19742 vdd.n19741 92.5
R31801 vdd.n19185 vdd.n19184 92.5
R31802 vdd.n19198 vdd.n19197 92.5
R31803 vdd.n19210 vdd.n19209 92.5
R31804 vdd.n19222 vdd.n19221 92.5
R31805 vdd.n19711 vdd.n19710 92.5
R31806 vdd.n19695 vdd.n19694 92.5
R31807 vdd.n19679 vdd.n19678 92.5
R31808 vdd.n19663 vdd.n19662 92.5
R31809 vdd.n19647 vdd.n19646 92.5
R31810 vdd.n19634 vdd.n19633 92.5
R31811 vdd.n19617 vdd.n19616 92.5
R31812 vdd.n19604 vdd.n19603 92.5
R31813 vdd.n19588 vdd.n19587 92.5
R31814 vdd.n19572 vdd.n19571 92.5
R31815 vdd.n19556 vdd.n19555 92.5
R31816 vdd.n19540 vdd.n19539 92.5
R31817 vdd.n19242 vdd.n19241 92.5
R31818 vdd.n19254 vdd.n19253 92.5
R31819 vdd.n19266 vdd.n19265 92.5
R31820 vdd.n19278 vdd.n19277 92.5
R31821 vdd.n19510 vdd.n19509 92.5
R31822 vdd.n19495 vdd.n19494 92.5
R31823 vdd.n19479 vdd.n19478 92.5
R31824 vdd.n19463 vdd.n19462 92.5
R31825 vdd.n19447 vdd.n19446 92.5
R31826 vdd.n19431 vdd.n19430 92.5
R31827 vdd.n19414 vdd.n19413 92.5
R31828 vdd.n19398 vdd.n19397 92.5
R31829 vdd.n19382 vdd.n19381 92.5
R31830 vdd.n19366 vdd.n19365 92.5
R31831 vdd.n19350 vdd.n19349 92.5
R31832 vdd.n20517 vdd.n20516 92.5
R31833 vdd.n20520 vdd.n20519 92.5
R31834 vdd.n19963 vdd.n19962 92.5
R31835 vdd.n19965 vdd.n19964 92.5
R31836 vdd.n19967 vdd.n19966 92.5
R31837 vdd.n19287 vdd.n19286 92.5
R31838 vdd.n19231 vdd.n19230 92.5
R31839 vdd.n19175 vdd.n19174 92.5
R31840 vdd.n19895 vdd.n19894 92.5
R31841 vdd.n19952 vdd.n19951 92.5
R31842 vdd.n20513 vdd.n20512 92.5
R31843 vdd.n20539 vdd.n20513 92.5
R31844 vdd.n20542 vdd.n20541 92.5
R31845 vdd.n20558 vdd.n20557 92.5
R31846 vdd.n20574 vdd.n20573 92.5
R31847 vdd.n20590 vdd.n20589 92.5
R31848 vdd.n20606 vdd.n20605 92.5
R31849 vdd.n20622 vdd.n20621 92.5
R31850 vdd.n20639 vdd.n20638 92.5
R31851 vdd.n20640 vdd.n20639 92.5
R31852 vdd.n20636 vdd.n20635 92.5
R31853 vdd.n20655 vdd.n20654 92.5
R31854 vdd.n20671 vdd.n20670 92.5
R31855 vdd.n20687 vdd.n20686 92.5
R31856 vdd.n20703 vdd.n20702 92.5
R31857 vdd.n20718 vdd.n20717 92.5
R31858 vdd.n19943 vdd.n19942 92.5
R31859 vdd.n19931 vdd.n19930 92.5
R31860 vdd.n20731 vdd.n20730 92.5
R31861 vdd.n20732 vdd.n20731 92.5
R31862 vdd.n19919 vdd.n19918 92.5
R31863 vdd.n19907 vdd.n19906 92.5
R31864 vdd.n20748 vdd.n20747 92.5
R31865 vdd.n20764 vdd.n20763 92.5
R31866 vdd.n20779 vdd.n20778 92.5
R31867 vdd.n20795 vdd.n20794 92.5
R31868 vdd.n20811 vdd.n20810 92.5
R31869 vdd.n20824 vdd.n20823 92.5
R31870 vdd.n20841 vdd.n20840 92.5
R31871 vdd.n20842 vdd.n20841 92.5
R31872 vdd.n20838 vdd.n20837 92.5
R31873 vdd.n20854 vdd.n20853 92.5
R31874 vdd.n19888 vdd.n19887 92.5
R31875 vdd.n20875 vdd.n20874 92.5
R31876 vdd.n20891 vdd.n20890 92.5
R31877 vdd.n20907 vdd.n20906 92.5
R31878 vdd.n19875 vdd.n19874 92.5
R31879 vdd.n19863 vdd.n19862 92.5
R31880 vdd.n20920 vdd.n20919 92.5
R31881 vdd.n20921 vdd.n20920 92.5
R31882 vdd.n19851 vdd.n19850 92.5
R31883 vdd.n19838 vdd.n19837 92.5
R31884 vdd.n20938 vdd.n20937 92.5
R31885 vdd.n20954 vdd.n20953 92.5
R31886 vdd.n20970 vdd.n20969 92.5
R31887 vdd.n20986 vdd.n20985 92.5
R31888 vdd.n19155 vdd.n19154 92.5
R31889 vdd.n19168 vdd.n19167 92.5
R31890 vdd.n19821 vdd.n19820 92.5
R31891 vdd.n19822 vdd.n19821 92.5
R31892 vdd.n19818 vdd.n19817 92.5
R31893 vdd.n19805 vdd.n19804 92.5
R31894 vdd.n19789 vdd.n19788 92.5
R31895 vdd.n19773 vdd.n19772 92.5
R31896 vdd.n19757 vdd.n19756 92.5
R31897 vdd.n19741 vdd.n19740 92.5
R31898 vdd.n19184 vdd.n19183 92.5
R31899 vdd.n19197 vdd.n19196 92.5
R31900 vdd.n19723 vdd.n19722 92.5
R31901 vdd.n19724 vdd.n19723 92.5
R31902 vdd.n19209 vdd.n19208 92.5
R31903 vdd.n19221 vdd.n19220 92.5
R31904 vdd.n19710 vdd.n19709 92.5
R31905 vdd.n19694 vdd.n19693 92.5
R31906 vdd.n19678 vdd.n19677 92.5
R31907 vdd.n19662 vdd.n19661 92.5
R31908 vdd.n19646 vdd.n19645 92.5
R31909 vdd.n19633 vdd.n19632 92.5
R31910 vdd.n19619 vdd.n19618 92.5
R31911 vdd.n19620 vdd.n19619 92.5
R31912 vdd.n19616 vdd.n19615 92.5
R31913 vdd.n19603 vdd.n19602 92.5
R31914 vdd.n19587 vdd.n19586 92.5
R31915 vdd.n19571 vdd.n19570 92.5
R31916 vdd.n19555 vdd.n19554 92.5
R31917 vdd.n19539 vdd.n19538 92.5
R31918 vdd.n19241 vdd.n19240 92.5
R31919 vdd.n19253 vdd.n19252 92.5
R31920 vdd.n19522 vdd.n19521 92.5
R31921 vdd.n19523 vdd.n19522 92.5
R31922 vdd.n19265 vdd.n19264 92.5
R31923 vdd.n19277 vdd.n19276 92.5
R31924 vdd.n19509 vdd.n19508 92.5
R31925 vdd.n19494 vdd.n19493 92.5
R31926 vdd.n19478 vdd.n19477 92.5
R31927 vdd.n19462 vdd.n19461 92.5
R31928 vdd.n19446 vdd.n19445 92.5
R31929 vdd.n19430 vdd.n19429 92.5
R31930 vdd.n19416 vdd.n19415 92.5
R31931 vdd.n19417 vdd.n19416 92.5
R31932 vdd.n19413 vdd.n19412 92.5
R31933 vdd.n19397 vdd.n19396 92.5
R31934 vdd.n19381 vdd.n19380 92.5
R31935 vdd.n19365 vdd.n19364 92.5
R31936 vdd.n19349 vdd.n19348 92.5
R31937 vdd.n19315 vdd.n19314 92.5
R31938 vdd.n19317 vdd.n19316 92.5
R31939 vdd.n19310 vdd.n19309 92.5
R31940 vdd.n19312 vdd.n19311 92.5
R31941 vdd.n19305 vdd.n19304 92.5
R31942 vdd.n19307 vdd.n19306 92.5
R31943 vdd.n19334 vdd.n19333 92.5
R31944 vdd.n19333 vdd.n19332 92.5
R31945 vdd.n19297 vdd.n19296 92.5
R31946 vdd.n20057 vdd.n20056 92.5
R31947 vdd.n20052 vdd.n20051 92.5
R31948 vdd.n20050 vdd.n20049 92.5
R31949 vdd.n20047 vdd.n20046 92.5
R31950 vdd.n20045 vdd.n20044 92.5
R31951 vdd.n20024 vdd.n20023 92.5
R31952 vdd.n20055 vdd.n20054 92.5
R31953 vdd.n20032 vdd.n20031 92.5
R31954 vdd.n20061 vdd.n20032 92.5
R31955 vdd.n20075 vdd.n20074 92.5
R31956 vdd.n20077 vdd.n20075 92.5
R31957 vdd.n20091 vdd.n20090 92.5
R31958 vdd.n20093 vdd.n20091 92.5
R31959 vdd.n20107 vdd.n20106 92.5
R31960 vdd.n20109 vdd.n20107 92.5
R31961 vdd.n20123 vdd.n20122 92.5
R31962 vdd.n20125 vdd.n20123 92.5
R31963 vdd.n20142 vdd.n20141 92.5
R31964 vdd.n20144 vdd.n20142 92.5
R31965 vdd.n20139 vdd.n20138 92.5
R31966 vdd.n20140 vdd.n20139 92.5
R31967 vdd.n20166 vdd.n20165 92.5
R31968 vdd.n20167 vdd.n20166 92.5
R31969 vdd.n20163 vdd.n20162 92.5
R31970 vdd.n20164 vdd.n20163 92.5
R31971 vdd.n20182 vdd.n20181 92.5
R31972 vdd.n20183 vdd.n20182 92.5
R31973 vdd.n20198 vdd.n20197 92.5
R31974 vdd.n20199 vdd.n20198 92.5
R31975 vdd.n20214 vdd.n20213 92.5
R31976 vdd.n20215 vdd.n20214 92.5
R31977 vdd.n20230 vdd.n20229 92.5
R31978 vdd.n20231 vdd.n20230 92.5
R31979 vdd.n20246 vdd.n20245 92.5
R31980 vdd.n20247 vdd.n20246 92.5
R31981 vdd.n20262 vdd.n20261 92.5
R31982 vdd.n20263 vdd.n20262 92.5
R31983 vdd.n20008 vdd.n20007 92.5
R31984 vdd.n20009 vdd.n20008 92.5
R31985 vdd.n19995 vdd.n19994 92.5
R31986 vdd.n19997 vdd.n19995 92.5
R31987 vdd.n20279 vdd.n20278 92.5
R31988 vdd.n20281 vdd.n20279 92.5
R31989 vdd.n20295 vdd.n20294 92.5
R31990 vdd.n20297 vdd.n20295 92.5
R31991 vdd.n20311 vdd.n20310 92.5
R31992 vdd.n20313 vdd.n20311 92.5
R31993 vdd.n20327 vdd.n20326 92.5
R31994 vdd.n20329 vdd.n20327 92.5
R31995 vdd.n20343 vdd.n20342 92.5
R31996 vdd.n20345 vdd.n20343 92.5
R31997 vdd.n20359 vdd.n20358 92.5
R31998 vdd.n20361 vdd.n20359 92.5
R31999 vdd.n20378 vdd.n20377 92.5
R32000 vdd.n20380 vdd.n20378 92.5
R32001 vdd.n20375 vdd.n20374 92.5
R32002 vdd.n20376 vdd.n20375 92.5
R32003 vdd.n20402 vdd.n20401 92.5
R32004 vdd.n20403 vdd.n20402 92.5
R32005 vdd.n20399 vdd.n20398 92.5
R32006 vdd.n20400 vdd.n20399 92.5
R32007 vdd.n20418 vdd.n20417 92.5
R32008 vdd.n20419 vdd.n20418 92.5
R32009 vdd.n20434 vdd.n20433 92.5
R32010 vdd.n20435 vdd.n20434 92.5
R32011 vdd.n20450 vdd.n20449 92.5
R32012 vdd.n19977 vdd.n19975 92.5
R32013 vdd.n20471 vdd.n19974 92.5
R32014 vdd.n20507 vdd.n20506 92.5
R32015 vdd.n20502 vdd.n20501 92.5
R32016 vdd.n20504 vdd.n20503 92.5
R32017 vdd.n20497 vdd.n20496 92.5
R32018 vdd.n20499 vdd.n20498 92.5
R32019 vdd.n20492 vdd.n20491 92.5
R32020 vdd.n20494 vdd.n20493 92.5
R32021 vdd.n20487 vdd.n20486 92.5
R32022 vdd.n20489 vdd.n20488 92.5
R32023 vdd.n20482 vdd.n20481 92.5
R32024 vdd.n20484 vdd.n20483 92.5
R32025 vdd.n20474 vdd.n20473 92.5
R32026 vdd.n20479 vdd.n20478 92.5
R32027 vdd.n20509 vdd.n20508 92.5
R32028 vdd.n20387 vdd.n20386 92.5
R32029 vdd.n20389 vdd.n20388 92.5
R32030 vdd.n20151 vdd.n20150 92.5
R32031 vdd.n20153 vdd.n20152 92.5
R32032 vdd.n24671 vdd.n24636 92.5
R32033 vdd.n24670 vdd.n24669 92.5
R32034 vdd.n24668 vdd.n24667 92.5
R32035 vdd.n24666 vdd.n24665 92.5
R32036 vdd.n24664 vdd.n24663 92.5
R32037 vdd.n24662 vdd.n24661 92.5
R32038 vdd.n24660 vdd.n24659 92.5
R32039 vdd.n24658 vdd.n24657 92.5
R32040 vdd.n24656 vdd.n24655 92.5
R32041 vdd.n24654 vdd.n24653 92.5
R32042 vdd.n24652 vdd.n24651 92.5
R32043 vdd.n24650 vdd.n24649 92.5
R32044 vdd.n24648 vdd.n24647 92.5
R32045 vdd.n24646 vdd.n24645 92.5
R32046 vdd.n24427 vdd.n24426 92.5
R32047 vdd.n24425 vdd.n24424 92.5
R32048 vdd.n24430 vdd.n24429 92.5
R32049 vdd.n24436 vdd.n24435 92.5
R32050 vdd.n24434 vdd.n24433 92.5
R32051 vdd.n24439 vdd.n24438 92.5
R32052 vdd.n24442 vdd.n24441 92.5
R32053 vdd.n24445 vdd.n24444 92.5
R32054 vdd.n24448 vdd.n24447 92.5
R32055 vdd.n24451 vdd.n24450 92.5
R32056 vdd.n24454 vdd.n24453 92.5
R32057 vdd.n24457 vdd.n24456 92.5
R32058 vdd.n24461 vdd.n24460 92.5
R32059 vdd.n24464 vdd.n24463 92.5
R32060 vdd.n24469 vdd.n24468 92.5
R32061 vdd.n24467 vdd.n24466 92.5
R32062 vdd.n24473 vdd.n24472 92.5
R32063 vdd.n24490 vdd.n24411 92.5
R32064 vdd.n25063 vdd.n25062 92.5
R32065 vdd.n25065 vdd.n25064 92.5
R32066 vdd.n25067 vdd.n25066 92.5
R32067 vdd.n25069 vdd.n25068 92.5
R32068 vdd.n25071 vdd.n25070 92.5
R32069 vdd.n25073 vdd.n25072 92.5
R32070 vdd.n25075 vdd.n25074 92.5
R32071 vdd.n25077 vdd.n25076 92.5
R32072 vdd.n25079 vdd.n25078 92.5
R32073 vdd.n25081 vdd.n25080 92.5
R32074 vdd.n25083 vdd.n25082 92.5
R32075 vdd.n25085 vdd.n25084 92.5
R32076 vdd.n25087 vdd.n25086 92.5
R32077 vdd.n25089 vdd.n25088 92.5
R32078 vdd.n24198 vdd.n24197 90.476
R32079 vdd.n23976 vdd.n23975 90.476
R32080 vdd.n23966 vdd.n23965 90.476
R32081 vdd.n23744 vdd.n23743 90.476
R32082 vdd.n23734 vdd.n23733 90.476
R32083 vdd.n23056 vdd.n23055 90.476
R32084 vdd.n23278 vdd.n23277 90.476
R32085 vdd.n23288 vdd.n23287 90.476
R32086 vdd.n23510 vdd.n23509 90.476
R32087 vdd.n23520 vdd.n23519 90.476
R32088 vdd.n22477 vdd.n22476 90.476
R32089 vdd.n22699 vdd.n22698 90.476
R32090 vdd.n22709 vdd.n22708 90.476
R32091 vdd.n22931 vdd.n22930 90.476
R32092 vdd.n22941 vdd.n22940 90.476
R32093 vdd.n22181 vdd.n22180 90.476
R32094 vdd.n22264 vdd.n22263 90.476
R32095 vdd.n22275 vdd.n22274 90.476
R32096 vdd.n22149 vdd.n22148 90.476
R32097 vdd.n22160 vdd.n22159 90.476
R32098 vdd.n11659 vdd.n11658 89.664
R32099 vdd.n24101 vdd.n24100 84.821
R32100 vdd.n24075 vdd.n24074 84.821
R32101 vdd.n23869 vdd.n23868 84.821
R32102 vdd.n23843 vdd.n23842 84.821
R32103 vdd.n23637 vdd.n23636 84.821
R32104 vdd.n23155 vdd.n23154 84.821
R32105 vdd.n23181 vdd.n23180 84.821
R32106 vdd.n23387 vdd.n23386 84.821
R32107 vdd.n23413 vdd.n23412 84.821
R32108 vdd.n23619 vdd.n23618 84.821
R32109 vdd.n22576 vdd.n22575 84.821
R32110 vdd.n22602 vdd.n22601 84.821
R32111 vdd.n22808 vdd.n22807 84.821
R32112 vdd.n22834 vdd.n22833 84.821
R32113 vdd.n23040 vdd.n23039 84.821
R32114 vdd.n22192 vdd.n22191 84.821
R32115 vdd.n22050 vdd.n22049 84.821
R32116 vdd.n22171 vdd.n22170 84.821
R32117 vdd.n14503 vdd.n14502 84.328
R32118 vdd.n13115 vdd.n13114 84.328
R32119 vdd.t82 vdd.t56 83.254
R32120 vdd.t339 vdd.t341 83.254
R32121 vdd.n14658 vdd.n8143 82.822
R32122 vdd.n14945 vdd.n14944 82.822
R32123 vdd.n20478 vdd.n20477 82.822
R32124 vdd.n24646 vdd.n24644 82.822
R32125 vdd.n25063 vdd.n25061 82.822
R32126 vdd.n10444 vdd.n10291 82.468
R32127 vdd.n13041 vdd.n9330 82.468
R32128 vdd.n12937 vdd.n9517 82.468
R32129 vdd.n12833 vdd.n9690 82.468
R32130 vdd.n12729 vdd.n9877 82.468
R32131 vdd.n12625 vdd.n10048 82.468
R32132 vdd.n24184 vdd.n24183 79.166
R32133 vdd.n23990 vdd.n23989 79.166
R32134 vdd.n23952 vdd.n23951 79.166
R32135 vdd.n23758 vdd.n23757 79.166
R32136 vdd.n23720 vdd.n23719 79.166
R32137 vdd.n23070 vdd.n23069 79.166
R32138 vdd.n23264 vdd.n23263 79.166
R32139 vdd.n23302 vdd.n23301 79.166
R32140 vdd.n23496 vdd.n23495 79.166
R32141 vdd.n23534 vdd.n23533 79.166
R32142 vdd.n22491 vdd.n22490 79.166
R32143 vdd.n22685 vdd.n22684 79.166
R32144 vdd.n22723 vdd.n22722 79.166
R32145 vdd.n22917 vdd.n22916 79.166
R32146 vdd.n22955 vdd.n22954 79.166
R32147 vdd.n22461 vdd.n22460 79.166
R32148 vdd.n22317 vdd.n22316 79.166
R32149 vdd.n24289 vdd.n24288 79.166
R32150 vdd.n13082 vdd.n9288 79.102
R32151 vdd.n9323 vdd.n9288 79.102
R32152 vdd.n9323 vdd.n9321 79.102
R32153 vdd.n13048 vdd.n9321 79.102
R32154 vdd.n13048 vdd.n9322 79.102
R32155 vdd.n13044 vdd.n9322 79.102
R32156 vdd.n13044 vdd.n9327 79.102
R32157 vdd.n13029 vdd.n9327 79.102
R32158 vdd.n13029 vdd.n9356 79.102
R32159 vdd.n13025 vdd.n9356 79.102
R32160 vdd.n13025 vdd.n9358 79.102
R32161 vdd.n9409 vdd.n9358 79.102
R32162 vdd.n12999 vdd.n9409 79.102
R32163 vdd.n12999 vdd.n9410 79.102
R32164 vdd.n12995 vdd.n9410 79.102
R32165 vdd.n12995 vdd.n9413 79.102
R32166 vdd.n9469 vdd.n9413 79.102
R32167 vdd.n9469 vdd.n9467 79.102
R32168 vdd.n12961 vdd.n9467 79.102
R32169 vdd.n12961 vdd.n9468 79.102
R32170 vdd.n12957 vdd.n9468 79.102
R32171 vdd.n12957 vdd.n9473 79.102
R32172 vdd.n9520 vdd.n9473 79.102
R32173 vdd.n12934 vdd.n9520 79.102
R32174 vdd.n12934 vdd.n9521 79.102
R32175 vdd.n12930 vdd.n9521 79.102
R32176 vdd.n12930 vdd.n9524 79.102
R32177 vdd.n9565 vdd.n9524 79.102
R32178 vdd.n12904 vdd.n9565 79.102
R32179 vdd.n12904 vdd.n9566 79.102
R32180 vdd.n12900 vdd.n9566 79.102
R32181 vdd.n12900 vdd.n9569 79.102
R32182 vdd.n9616 vdd.n9569 79.102
R32183 vdd.n12878 vdd.n9616 79.102
R32184 vdd.n12878 vdd.n9617 79.102
R32185 vdd.n12874 vdd.n9617 79.102
R32186 vdd.n12874 vdd.n9620 79.102
R32187 vdd.n9683 vdd.n9620 79.102
R32188 vdd.n9683 vdd.n9681 79.102
R32189 vdd.n12840 vdd.n9681 79.102
R32190 vdd.n12840 vdd.n9682 79.102
R32191 vdd.n12836 vdd.n9682 79.102
R32192 vdd.n12836 vdd.n9687 79.102
R32193 vdd.n12821 vdd.n9687 79.102
R32194 vdd.n12821 vdd.n9716 79.102
R32195 vdd.n12817 vdd.n9716 79.102
R32196 vdd.n12817 vdd.n9718 79.102
R32197 vdd.n9770 vdd.n9718 79.102
R32198 vdd.n12791 vdd.n9770 79.102
R32199 vdd.n12791 vdd.n9771 79.102
R32200 vdd.n12787 vdd.n9771 79.102
R32201 vdd.n12787 vdd.n9774 79.102
R32202 vdd.n9829 vdd.n9774 79.102
R32203 vdd.n9829 vdd.n9827 79.102
R32204 vdd.n12753 vdd.n9827 79.102
R32205 vdd.n12753 vdd.n9828 79.102
R32206 vdd.n12749 vdd.n9828 79.102
R32207 vdd.n12749 vdd.n9833 79.102
R32208 vdd.n9880 vdd.n9833 79.102
R32209 vdd.n12726 vdd.n9880 79.102
R32210 vdd.n12726 vdd.n9881 79.102
R32211 vdd.n12722 vdd.n9881 79.102
R32212 vdd.n12722 vdd.n9884 79.102
R32213 vdd.n9924 vdd.n9884 79.102
R32214 vdd.n12696 vdd.n9924 79.102
R32215 vdd.n12696 vdd.n9925 79.102
R32216 vdd.n12692 vdd.n9925 79.102
R32217 vdd.n12692 vdd.n9928 79.102
R32218 vdd.n9976 vdd.n9928 79.102
R32219 vdd.n12670 vdd.n9976 79.102
R32220 vdd.n12670 vdd.n9977 79.102
R32221 vdd.n12666 vdd.n9977 79.102
R32222 vdd.n12666 vdd.n9980 79.102
R32223 vdd.n10042 vdd.n9980 79.102
R32224 vdd.n10042 vdd.n10040 79.102
R32225 vdd.n12632 vdd.n10040 79.102
R32226 vdd.n12632 vdd.n10041 79.102
R32227 vdd.n12628 vdd.n10041 79.102
R32228 vdd.n12628 vdd.n10046 79.102
R32229 vdd.n12612 vdd.n10046 79.102
R32230 vdd.n12612 vdd.n10058 79.102
R32231 vdd.n12608 vdd.n10058 79.102
R32232 vdd.n12608 vdd.n10060 79.102
R32233 vdd.n10113 vdd.n10060 79.102
R32234 vdd.n12593 vdd.n10113 79.102
R32235 vdd.n12593 vdd.n10114 79.102
R32236 vdd.n12589 vdd.n10114 79.102
R32237 vdd.n12589 vdd.n10117 79.102
R32238 vdd.n10495 vdd.n10117 79.102
R32239 vdd.n12565 vdd.n10495 79.102
R32240 vdd.n12565 vdd.n10496 79.102
R32241 vdd.n12561 vdd.n10496 79.102
R32242 vdd.n12561 vdd.n10499 79.102
R32243 vdd.n12557 vdd.n10499 79.102
R32244 vdd.n12557 vdd.n10502 79.102
R32245 vdd.n12553 vdd.n10502 79.102
R32246 vdd.n12553 vdd.n10504 79.102
R32247 vdd.n12549 vdd.n10504 79.102
R32248 vdd.n12549 vdd.n10506 79.102
R32249 vdd.n12545 vdd.n10506 79.102
R32250 vdd.n12545 vdd.n10508 79.102
R32251 vdd.n12541 vdd.n10508 79.102
R32252 vdd.n12541 vdd.n10509 79.102
R32253 vdd.n12537 vdd.n10509 79.102
R32254 vdd.n12537 vdd.n10511 79.102
R32255 vdd.n12533 vdd.n10511 79.102
R32256 vdd.n12533 vdd.n10514 79.102
R32257 vdd.n12529 vdd.n10514 79.102
R32258 vdd.n12529 vdd.n10516 79.102
R32259 vdd.n12518 vdd.n10516 79.102
R32260 vdd.n12518 vdd.n10525 79.102
R32261 vdd.n12514 vdd.n10525 79.102
R32262 vdd.n12514 vdd.n10527 79.102
R32263 vdd.n10578 vdd.n10527 79.102
R32264 vdd.n12487 vdd.n10578 79.102
R32265 vdd.n12487 vdd.n10579 79.102
R32266 vdd.n12483 vdd.n10579 79.102
R32267 vdd.n12483 vdd.n10582 79.102
R32268 vdd.n10617 vdd.n10582 79.102
R32269 vdd.n12458 vdd.n10617 79.102
R32270 vdd.n12458 vdd.n10618 79.102
R32271 vdd.n12454 vdd.n10618 79.102
R32272 vdd.n12454 vdd.n10621 79.102
R32273 vdd.n10666 vdd.n10621 79.102
R32274 vdd.n12430 vdd.n10666 79.102
R32275 vdd.n12430 vdd.n10667 79.102
R32276 vdd.n12426 vdd.n10667 79.102
R32277 vdd.n12426 vdd.n10670 79.102
R32278 vdd.n10714 vdd.n10670 79.102
R32279 vdd.n12399 vdd.n10714 79.102
R32280 vdd.n12399 vdd.n10715 79.102
R32281 vdd.n12395 vdd.n10715 79.102
R32282 vdd.n12395 vdd.n10718 79.102
R32283 vdd.n10768 vdd.n10718 79.102
R32284 vdd.n10768 vdd.n10766 79.102
R32285 vdd.n12369 vdd.n10766 79.102
R32286 vdd.n12369 vdd.n10767 79.102
R32287 vdd.n12365 vdd.n10767 79.102
R32288 vdd.n12365 vdd.n10772 79.102
R32289 vdd.n10819 vdd.n10772 79.102
R32290 vdd.n12340 vdd.n10819 79.102
R32291 vdd.n12340 vdd.n10820 79.102
R32292 vdd.n12336 vdd.n10820 79.102
R32293 vdd.n12336 vdd.n10823 79.102
R32294 vdd.n12322 vdd.n10823 79.102
R32295 vdd.n12322 vdd.n10863 79.102
R32296 vdd.n12318 vdd.n10863 79.102
R32297 vdd.n12318 vdd.n10865 79.102
R32298 vdd.n10910 vdd.n10865 79.102
R32299 vdd.n12291 vdd.n10910 79.102
R32300 vdd.n12291 vdd.n10911 79.102
R32301 vdd.n12287 vdd.n10911 79.102
R32302 vdd.n12287 vdd.n10914 79.102
R32303 vdd.n10954 vdd.n10914 79.102
R32304 vdd.n12268 vdd.n10954 79.102
R32305 vdd.n12268 vdd.n10955 79.102
R32306 vdd.n12264 vdd.n10955 79.102
R32307 vdd.n12264 vdd.n10958 79.102
R32308 vdd.n11006 vdd.n10958 79.102
R32309 vdd.n12239 vdd.n11006 79.102
R32310 vdd.n12239 vdd.n11007 79.102
R32311 vdd.n12235 vdd.n11007 79.102
R32312 vdd.n12235 vdd.n11010 79.102
R32313 vdd.n11051 vdd.n11010 79.102
R32314 vdd.n12208 vdd.n11051 79.102
R32315 vdd.n12208 vdd.n11052 79.102
R32316 vdd.n12204 vdd.n11052 79.102
R32317 vdd.n12204 vdd.n11055 79.102
R32318 vdd.n11100 vdd.n11055 79.102
R32319 vdd.n12178 vdd.n11100 79.102
R32320 vdd.n12178 vdd.n11101 79.102
R32321 vdd.n12174 vdd.n11101 79.102
R32322 vdd.n12174 vdd.n11104 79.102
R32323 vdd.n11140 vdd.n11104 79.102
R32324 vdd.n12149 vdd.n11140 79.102
R32325 vdd.n12149 vdd.n11141 79.102
R32326 vdd.n12145 vdd.n11141 79.102
R32327 vdd.n12145 vdd.n11144 79.102
R32328 vdd.n11186 vdd.n11144 79.102
R32329 vdd.n12120 vdd.n11186 79.102
R32330 vdd.n12120 vdd.n11187 79.102
R32331 vdd.n12116 vdd.n11187 79.102
R32332 vdd.n12116 vdd.n11190 79.102
R32333 vdd.n11235 vdd.n11190 79.102
R32334 vdd.n12089 vdd.n11235 79.102
R32335 vdd.n12089 vdd.n11236 79.102
R32336 vdd.n12085 vdd.n11236 79.102
R32337 vdd.n12085 vdd.n11239 79.102
R32338 vdd.n11276 vdd.n11239 79.102
R32339 vdd.n12063 vdd.n11276 79.102
R32340 vdd.n12063 vdd.n11277 79.102
R32341 vdd.n12059 vdd.n11277 79.102
R32342 vdd.n12059 vdd.n11280 79.102
R32343 vdd.n11328 vdd.n11280 79.102
R32344 vdd.n12034 vdd.n11328 79.102
R32345 vdd.n12034 vdd.n11329 79.102
R32346 vdd.n12030 vdd.n11329 79.102
R32347 vdd.n12030 vdd.n11332 79.102
R32348 vdd.n12016 vdd.n11332 79.102
R32349 vdd.n12016 vdd.n11372 79.102
R32350 vdd.n12012 vdd.n11372 79.102
R32351 vdd.n12012 vdd.n11374 79.102
R32352 vdd.n11419 vdd.n11374 79.102
R32353 vdd.n11985 vdd.n11419 79.102
R32354 vdd.n11985 vdd.n11420 79.102
R32355 vdd.n11981 vdd.n11420 79.102
R32356 vdd.n11981 vdd.n11423 79.102
R32357 vdd.n11439 vdd.n11423 79.102
R32358 vdd.n11962 vdd.n11439 79.102
R32359 vdd.n11962 vdd.n11440 79.102
R32360 vdd.n11958 vdd.n11440 79.102
R32361 vdd.n11958 vdd.n11443 79.102
R32362 vdd.n11932 vdd.n11443 79.102
R32363 vdd.n11932 vdd.n11561 79.102
R32364 vdd.n11928 vdd.n11561 79.102
R32365 vdd.n11928 vdd.n11563 79.102
R32366 vdd.n14617 vdd.n8170 79.058
R32367 vdd.n11631 vdd.n11577 79.058
R32368 vdd.n11924 vdd.n11563 78.549
R32369 vdd.n10477 vdd.t82 75.509
R32370 vdd.n15260 vdd.t339 75.509
R32371 vdd.n24115 vdd.n24114 73.511
R32372 vdd.n24061 vdd.n24060 73.511
R32373 vdd.n23883 vdd.n23882 73.511
R32374 vdd.n23829 vdd.n23828 73.511
R32375 vdd.n23651 vdd.n23650 73.511
R32376 vdd.n23141 vdd.n23140 73.511
R32377 vdd.n23195 vdd.n23194 73.511
R32378 vdd.n23373 vdd.n23372 73.511
R32379 vdd.n23427 vdd.n23426 73.511
R32380 vdd.n23605 vdd.n23604 73.511
R32381 vdd.n22562 vdd.n22561 73.511
R32382 vdd.n22616 vdd.n22615 73.511
R32383 vdd.n22794 vdd.n22793 73.511
R32384 vdd.n22848 vdd.n22847 73.511
R32385 vdd.n23026 vdd.n23025 73.511
R32386 vdd.n22389 vdd.n22388 73.511
R32387 vdd.n22359 vdd.n22358 73.511
R32388 vdd.n24334 vdd.n24333 73.511
R32389 vdd.n22088 vdd.n22087 73.511
R32390 vdd.n24217 vdd.n24216 73.511
R32391 vdd.n18493 vdd.n18492 71.074
R32392 vdd.n14782 vdd.n8075 70.758
R32393 vdd.n30500 vdd.n30351 67.954
R32394 vdd.n30500 vdd.n30354 67.954
R32395 vdd.n30500 vdd.n30356 67.954
R32396 vdd.n30500 vdd.n30358 67.954
R32397 vdd.n30500 vdd.n30359 67.954
R32398 vdd.n30500 vdd.n30363 67.954
R32399 vdd.n30500 vdd.n30366 67.954
R32400 vdd.n30500 vdd.n30367 67.954
R32401 vdd.n30500 vdd.n30372 67.954
R32402 vdd.n30500 vdd.n30375 67.954
R32403 vdd.n30500 vdd.n30378 67.954
R32404 vdd.n30500 vdd.n30381 67.954
R32405 vdd.n30500 vdd.n30384 67.954
R32406 vdd.n30500 vdd.n30387 67.954
R32407 vdd.n30500 vdd.n30388 67.954
R32408 vdd.n30500 vdd.n30391 67.954
R32409 vdd.n30500 vdd.n30396 67.954
R32410 vdd.n30500 vdd.n30397 67.954
R32411 vdd.n30500 vdd.n30400 67.954
R32412 vdd.n30500 vdd.n30405 67.954
R32413 vdd.n30500 vdd.n30406 67.954
R32414 vdd.n30500 vdd.n30411 67.954
R32415 vdd.n30500 vdd.n30412 67.954
R32416 vdd.n30500 vdd.n30415 67.954
R32417 vdd.n30500 vdd.n30420 67.954
R32418 vdd.n30500 vdd.n30423 67.954
R32419 vdd.n30500 vdd.n30424 67.954
R32420 vdd.n30500 vdd.n30429 67.954
R32421 vdd.n30500 vdd.n30432 67.954
R32422 vdd.n30500 vdd.n30433 67.954
R32423 vdd.n30500 vdd.n30438 67.954
R32424 vdd.n30500 vdd.n30439 67.954
R32425 vdd.n30500 vdd.n30442 67.954
R32426 vdd.n30500 vdd.n30447 67.954
R32427 vdd.n30500 vdd.n30450 67.954
R32428 vdd.n30500 vdd.n30451 67.954
R32429 vdd.n30500 vdd.n30456 67.954
R32430 vdd.n30500 vdd.n30457 67.954
R32431 vdd.n30500 vdd.n30462 67.954
R32432 vdd.n30500 vdd.n30465 67.954
R32433 vdd.n30500 vdd.n30466 67.954
R32434 vdd.n30500 vdd.n30469 67.954
R32435 vdd.n30500 vdd.n30474 67.954
R32436 vdd.n30500 vdd.n30477 67.954
R32437 vdd.n30500 vdd.n30480 67.954
R32438 vdd.n30500 vdd.n30483 67.954
R32439 vdd.n30500 vdd.n30485 67.954
R32440 vdd.n30500 vdd.n30487 67.954
R32441 vdd.n30500 vdd.n30488 67.954
R32442 vdd.n30500 vdd.n30490 67.954
R32443 vdd.n30500 vdd.n30493 67.954
R32444 vdd.n30500 vdd.n30495 67.954
R32445 vdd.n30500 vdd.n30496 67.954
R32446 vdd.n14969 vdd.n7990 67.954
R32447 vdd.n14969 vdd.n7991 67.954
R32448 vdd.n14969 vdd.n7992 67.954
R32449 vdd.n14969 vdd.n7993 67.954
R32450 vdd.n14969 vdd.n7994 67.954
R32451 vdd.n14969 vdd.n7995 67.954
R32452 vdd.n14969 vdd.n7996 67.954
R32453 vdd.n14969 vdd.n7997 67.954
R32454 vdd.n14969 vdd.n7998 67.954
R32455 vdd.n14969 vdd.n14968 67.954
R32456 vdd.n14530 vdd.n8200 67.954
R32457 vdd.n14530 vdd.n8201 67.954
R32458 vdd.n14530 vdd.n8202 67.954
R32459 vdd.n14530 vdd.n8203 67.954
R32460 vdd.n14530 vdd.n8204 67.954
R32461 vdd.n14530 vdd.n8205 67.954
R32462 vdd.n14530 vdd.n8206 67.954
R32463 vdd.n14530 vdd.n8207 67.954
R32464 vdd.n14530 vdd.n8208 67.954
R32465 vdd.n14530 vdd.n8209 67.954
R32466 vdd.n20539 vdd.n20521 67.954
R32467 vdd.n20539 vdd.n20522 67.954
R32468 vdd.n20539 vdd.n20524 67.954
R32469 vdd.n20539 vdd.n20527 67.954
R32470 vdd.n20539 vdd.n20529 67.954
R32471 vdd.n20539 vdd.n20530 67.954
R32472 vdd.n20539 vdd.n20532 67.954
R32473 vdd.n20539 vdd.n20534 67.954
R32474 vdd.n20539 vdd.n20536 67.954
R32475 vdd.n20539 vdd.n20537 67.954
R32476 vdd.n24490 vdd.n24416 67.954
R32477 vdd.n24490 vdd.n24418 67.954
R32478 vdd.n24490 vdd.n24419 67.954
R32479 vdd.n24490 vdd.n24421 67.954
R32480 vdd.n24490 vdd.n24423 67.954
R32481 vdd.n24490 vdd.n24428 67.954
R32482 vdd.n24490 vdd.n24431 67.954
R32483 vdd.n24490 vdd.n24432 67.954
R32484 vdd.n24490 vdd.n24437 67.954
R32485 vdd.n24490 vdd.n24440 67.954
R32486 vdd.n24490 vdd.n24443 67.954
R32487 vdd.n24490 vdd.n24446 67.954
R32488 vdd.n24490 vdd.n24449 67.954
R32489 vdd.n24490 vdd.n24452 67.954
R32490 vdd.n24490 vdd.n24455 67.954
R32491 vdd.n24490 vdd.n24458 67.954
R32492 vdd.n24490 vdd.n24459 67.954
R32493 vdd.n24490 vdd.n24462 67.954
R32494 vdd.n24490 vdd.n24465 67.954
R32495 vdd.n24490 vdd.n24470 67.954
R32496 vdd.n24490 vdd.n24471 67.954
R32497 vdd.n24490 vdd.n24474 67.954
R32498 vdd.n24490 vdd.n24476 67.954
R32499 vdd.n24490 vdd.n24478 67.954
R32500 vdd.n24490 vdd.n24481 67.954
R32501 vdd.n24490 vdd.n24482 67.954
R32502 vdd.n24490 vdd.n24485 67.954
R32503 vdd.n24490 vdd.n24486 67.954
R32504 vdd.n24170 vdd.n24169 67.857
R32505 vdd.n24004 vdd.n24003 67.857
R32506 vdd.n23938 vdd.n23937 67.857
R32507 vdd.n23772 vdd.n23771 67.857
R32508 vdd.n23706 vdd.n23705 67.857
R32509 vdd.n23084 vdd.n23083 67.857
R32510 vdd.n23250 vdd.n23249 67.857
R32511 vdd.n23316 vdd.n23315 67.857
R32512 vdd.n23482 vdd.n23481 67.857
R32513 vdd.n23548 vdd.n23547 67.857
R32514 vdd.n22505 vdd.n22504 67.857
R32515 vdd.n22671 vdd.n22670 67.857
R32516 vdd.n22737 vdd.n22736 67.857
R32517 vdd.n22903 vdd.n22902 67.857
R32518 vdd.n22969 vdd.n22968 67.857
R32519 vdd.n22445 vdd.n22444 67.857
R32520 vdd.n22250 vdd.n22249 67.857
R32521 vdd.n22301 vdd.n22300 67.857
R32522 vdd.n22126 vdd.n22125 67.857
R32523 vdd.n24273 vdd.n24272 67.857
R32524 vdd.n11924 vdd.n11566 66.787
R32525 vdd.n15005 vdd.n15004 66.787
R32526 vdd.n12526 vdd.n10517 65.489
R32527 vdd.n11600 vdd.n11559 65.489
R32528 vdd.n16870 vdd.n16835 65.489
R32529 vdd.n24741 vdd.n24740 64.569
R32530 vdd.n25173 vdd.n25172 64.569
R32531 vdd.n12522 vdd.n10522 64.276
R32532 vdd.n10551 vdd.n10537 64.276
R32533 vdd.n10555 vdd.n10530 64.276
R32534 vdd.n12504 vdd.n10531 64.276
R32535 vdd.n12500 vdd.n10565 64.276
R32536 vdd.n12490 vdd.n10571 64.276
R32537 vdd.n10599 vdd.n10595 64.276
R32538 vdd.n12473 vdd.n10586 64.276
R32539 vdd.n12469 vdd.n10606 64.276
R32540 vdd.n12462 vdd.n10613 64.276
R32541 vdd.n10644 vdd.n10632 64.276
R32542 vdd.n10648 vdd.n10624 64.276
R32543 vdd.n12444 vdd.n10625 64.276
R32544 vdd.n12440 vdd.n10657 64.276
R32545 vdd.n10691 vdd.n10673 64.276
R32546 vdd.n12416 vdd.n10674 64.276
R32547 vdd.n12412 vdd.n10700 64.276
R32548 vdd.n12402 vdd.n10706 64.276
R32549 vdd.n10736 vdd.n10728 64.276
R32550 vdd.n10740 vdd.n10721 64.276
R32551 vdd.n12385 vdd.n10722 64.276
R32552 vdd.n12381 vdd.n10750 64.276
R32553 vdd.n12373 vdd.n10756 64.276
R32554 vdd.n10795 vdd.n10783 64.276
R32555 vdd.n10799 vdd.n10775 64.276
R32556 vdd.n12355 vdd.n10776 64.276
R32557 vdd.n12351 vdd.n10808 64.276
R32558 vdd.n12344 vdd.n10815 64.276
R32559 vdd.n10843 vdd.n10842 64.276
R32560 vdd.n12325 vdd.n10856 64.276
R32561 vdd.n10883 vdd.n10875 64.276
R32562 vdd.n10887 vdd.n10868 64.276
R32563 vdd.n12308 vdd.n10869 64.276
R32564 vdd.n12304 vdd.n10897 64.276
R32565 vdd.n12294 vdd.n10903 64.276
R32566 vdd.n10936 vdd.n10928 64.276
R32567 vdd.n10940 vdd.n10916 64.276
R32568 vdd.n12276 vdd.n10921 64.276
R32569 vdd.n12272 vdd.n10951 64.276
R32570 vdd.n10982 vdd.n10969 64.276
R32571 vdd.n10986 vdd.n10961 64.276
R32572 vdd.n12254 vdd.n10962 64.276
R32573 vdd.n12250 vdd.n10995 64.276
R32574 vdd.n12243 vdd.n11002 64.276
R32575 vdd.n12225 vdd.n11014 64.276
R32576 vdd.n12221 vdd.n11037 64.276
R32577 vdd.n12211 vdd.n11043 64.276
R32578 vdd.n11073 vdd.n11065 64.276
R32579 vdd.n11077 vdd.n11058 64.276
R32580 vdd.n12194 vdd.n11059 64.276
R32581 vdd.n12190 vdd.n11087 64.276
R32582 vdd.n12180 vdd.n11093 64.276
R32583 vdd.n11120 vdd.n11107 64.276
R32584 vdd.n12164 vdd.n11108 64.276
R32585 vdd.n12160 vdd.n11129 64.276
R32586 vdd.n12153 vdd.n11136 64.276
R32587 vdd.n11167 vdd.n11155 64.276
R32588 vdd.n11170 vdd.n11147 64.276
R32589 vdd.n12135 vdd.n11148 64.276
R32590 vdd.n11208 vdd.n11200 64.276
R32591 vdd.n11212 vdd.n11193 64.276
R32592 vdd.n12106 vdd.n11194 64.276
R32593 vdd.n12102 vdd.n11222 64.276
R32594 vdd.n12092 vdd.n11228 64.276
R32595 vdd.n11257 vdd.n11249 64.276
R32596 vdd.n11261 vdd.n11242 64.276
R32597 vdd.n12075 vdd.n11243 64.276
R32598 vdd.n12067 vdd.n11272 64.276
R32599 vdd.n11304 vdd.n11291 64.276
R32600 vdd.n11308 vdd.n11283 64.276
R32601 vdd.n12049 vdd.n11284 64.276
R32602 vdd.n12045 vdd.n11317 64.276
R32603 vdd.n12038 vdd.n11324 64.276
R32604 vdd.n11352 vdd.n11351 64.276
R32605 vdd.n12019 vdd.n11365 64.276
R32606 vdd.n11392 vdd.n11384 64.276
R32607 vdd.n11396 vdd.n11377 64.276
R32608 vdd.n12002 vdd.n11378 64.276
R32609 vdd.n11998 vdd.n11406 64.276
R32610 vdd.n11988 vdd.n11412 64.276
R32611 vdd.n11480 vdd.n11472 64.276
R32612 vdd.n11484 vdd.n11425 64.276
R32613 vdd.n11970 vdd.n11430 64.276
R32614 vdd.n11966 vdd.n11436 64.276
R32615 vdd.n11524 vdd.n11523 64.276
R32616 vdd.n11525 vdd.n11446 64.276
R32617 vdd.n11947 vdd.n11447 64.276
R32618 vdd.n11943 vdd.n11550 64.276
R32619 vdd.n10474 vdd.n10273 64.276
R32620 vdd.n10468 vdd.n10278 64.276
R32621 vdd.n10456 vdd.n10280 64.276
R32622 vdd.n10452 vdd.n10291 64.276
R32623 vdd.n10444 vdd.n10296 64.276
R32624 vdd.n10432 vdd.n10298 64.276
R32625 vdd.n10428 vdd.n10308 64.276
R32626 vdd.n10418 vdd.n10314 64.276
R32627 vdd.n10414 vdd.n10321 64.276
R32628 vdd.n10402 vdd.n10325 64.276
R32629 vdd.n10395 vdd.n10336 64.276
R32630 vdd.n10390 vdd.n10337 64.276
R32631 vdd.n10378 vdd.n10345 64.276
R32632 vdd.n10371 vdd.n10356 64.276
R32633 vdd.n13079 vdd.n9291 64.276
R32634 vdd.n13075 vdd.n9296 64.276
R32635 vdd.n13062 vdd.n9299 64.276
R32636 vdd.n13058 vdd.n9309 64.276
R32637 vdd.n13051 vdd.n9316 64.276
R32638 vdd.n9344 vdd.n9330 64.276
R32639 vdd.n13041 vdd.n9331 64.276
R32640 vdd.n9375 vdd.n9353 64.276
R32641 vdd.n9382 vdd.n9367 64.276
R32642 vdd.n13022 vdd.n9361 64.276
R32643 vdd.n13015 vdd.n9397 64.276
R32644 vdd.n13011 vdd.n9402 64.276
R32645 vdd.n13002 vdd.n9408 64.276
R32646 vdd.n9443 vdd.n9433 64.276
R32647 vdd.n12988 vdd.n9420 64.276
R32648 vdd.n12975 vdd.n9422 64.276
R32649 vdd.n12971 vdd.n9456 64.276
R32650 vdd.n12964 vdd.n9463 64.276
R32651 vdd.n9495 vdd.n9482 64.276
R32652 vdd.n12954 vdd.n9476 64.276
R32653 vdd.n12950 vdd.n9507 64.276
R32654 vdd.n12937 vdd.n9509 64.276
R32655 vdd.n9537 vdd.n9517 64.276
R32656 vdd.n12927 vdd.n9526 64.276
R32657 vdd.n12920 vdd.n9552 64.276
R32658 vdd.n12916 vdd.n9557 64.276
R32659 vdd.n12907 vdd.n9563 64.276
R32660 vdd.n9592 vdd.n9578 64.276
R32661 vdd.n12897 vdd.n9572 64.276
R32662 vdd.n12890 vdd.n9606 64.276
R32663 vdd.n9636 vdd.n9613 64.276
R32664 vdd.n9645 vdd.n9629 64.276
R32665 vdd.n12871 vdd.n9623 64.276
R32666 vdd.n12867 vdd.n9657 64.276
R32667 vdd.n12854 vdd.n9659 64.276
R32668 vdd.n12850 vdd.n9670 64.276
R32669 vdd.n12843 vdd.n9677 64.276
R32670 vdd.n9704 vdd.n9690 64.276
R32671 vdd.n12833 vdd.n9691 64.276
R32672 vdd.n9735 vdd.n9713 64.276
R32673 vdd.n9742 vdd.n9727 64.276
R32674 vdd.n12814 vdd.n9721 64.276
R32675 vdd.n12807 vdd.n9757 64.276
R32676 vdd.n12803 vdd.n9762 64.276
R32677 vdd.n12794 vdd.n9768 64.276
R32678 vdd.n9802 vdd.n9793 64.276
R32679 vdd.n12780 vdd.n9781 64.276
R32680 vdd.n12767 vdd.n9782 64.276
R32681 vdd.n12763 vdd.n9816 64.276
R32682 vdd.n12756 vdd.n9823 64.276
R32683 vdd.n9855 vdd.n9842 64.276
R32684 vdd.n12746 vdd.n9836 64.276
R32685 vdd.n12742 vdd.n9867 64.276
R32686 vdd.n12729 vdd.n9869 64.276
R32687 vdd.n9898 vdd.n9877 64.276
R32688 vdd.n12719 vdd.n9887 64.276
R32689 vdd.n12712 vdd.n9912 64.276
R32690 vdd.n12708 vdd.n9916 64.276
R32691 vdd.n12699 vdd.n9921 64.276
R32692 vdd.n9952 vdd.n9937 64.276
R32693 vdd.n12689 vdd.n9931 64.276
R32694 vdd.n12682 vdd.n9966 64.276
R32695 vdd.n9996 vdd.n9973 64.276
R32696 vdd.n10005 vdd.n9989 64.276
R32697 vdd.n12663 vdd.n9983 64.276
R32698 vdd.n12659 vdd.n10017 64.276
R32699 vdd.n12646 vdd.n10019 64.276
R32700 vdd.n12642 vdd.n10030 64.276
R32701 vdd.n12635 vdd.n10037 64.276
R32702 vdd.n10158 vdd.n10048 64.276
R32703 vdd.n12625 vdd.n10049 64.276
R32704 vdd.n10140 vdd.n10055 64.276
R32705 vdd.n10187 vdd.n10138 64.276
R32706 vdd.n12605 vdd.n10063 64.276
R32707 vdd.n10108 vdd.n10064 64.276
R32708 vdd.n10110 vdd.n10099 64.276
R32709 vdd.n10229 vdd.n10101 64.276
R32710 vdd.n10245 vdd.n10238 64.276
R32711 vdd.n10483 vdd.n10481 64.276
R32712 vdd.n10492 vdd.n10489 64.276
R32713 vdd.n15304 vdd.n15299 64.276
R32714 vdd.n15325 vdd.n15318 64.276
R32715 vdd.n15532 vdd.n15524 64.276
R32716 vdd.n15559 vdd.n15546 64.276
R32717 vdd.n15788 vdd.n15780 64.276
R32718 vdd.n15815 vdd.n15802 64.276
R32719 vdd.n16044 vdd.n16036 64.276
R32720 vdd.n16071 vdd.n16058 64.276
R32721 vdd.n16300 vdd.n16292 64.276
R32722 vdd.n16327 vdd.n16314 64.276
R32723 vdd.n16572 vdd.n16547 64.276
R32724 vdd.n14641 vdd.n8169 63.999
R32725 vdd.n11655 vdd.n11576 63.999
R32726 vdd.n18461 vdd.n18460 63.999
R32727 vdd.n21643 vdd.n21642 63.999
R32728 vdd.n31141 vdd.n31140 63.623
R32729 vdd.n30332 vdd.n30331 63.623
R32730 vdd.n35706 vdd.n35705 63.623
R32731 vdd.n2735 vdd.n2734 63.623
R32732 vdd.n12433 vdd.n10664 63.063
R32733 vdd.n10687 vdd.n10664 63.063
R32734 vdd.n12334 vdd.n10826 63.063
R32735 vdd.n12334 vdd.n10827 63.063
R32736 vdd.n11029 vdd.n11027 63.063
R32737 vdd.n11029 vdd.n11013 63.063
R32738 vdd.n12131 vdd.n11178 63.063
R32739 vdd.n12123 vdd.n11178 63.063
R32740 vdd.n12028 vdd.n11335 63.063
R32741 vdd.n12028 vdd.n11336 63.063
R32742 vdd.n17124 vdd.n17113 63.063
R32743 vdd.n17396 vdd.n17385 63.063
R32744 vdd.n17654 vdd.n17643 63.063
R32745 vdd.n17925 vdd.n17914 63.063
R32746 vdd.n18197 vdd.n18186 63.063
R32747 vdd.n11844 vdd.t224 62.35
R32748 vdd.n21935 vdd.t194 62.35
R32749 vdd.n11701 vdd.t185 62.347
R32750 vdd.n21772 vdd.t176 62.347
R32751 vdd.n11701 vdd.t189 62.339
R32752 vdd.n21772 vdd.t219 62.339
R32753 vdd.n11844 vdd.t211 62.336
R32754 vdd.n21935 vdd.t180 62.336
R32755 vdd.n24129 vdd.n24128 62.202
R32756 vdd.n24047 vdd.n24046 62.202
R32757 vdd.n23897 vdd.n23896 62.202
R32758 vdd.n23815 vdd.n23814 62.202
R32759 vdd.n23665 vdd.n23664 62.202
R32760 vdd.n23127 vdd.n23126 62.202
R32761 vdd.n23209 vdd.n23208 62.202
R32762 vdd.n23359 vdd.n23358 62.202
R32763 vdd.n23441 vdd.n23440 62.202
R32764 vdd.n23591 vdd.n23590 62.202
R32765 vdd.n22548 vdd.n22547 62.202
R32766 vdd.n22630 vdd.n22629 62.202
R32767 vdd.n22780 vdd.n22779 62.202
R32768 vdd.n22862 vdd.n22861 62.202
R32769 vdd.n23012 vdd.n23011 62.202
R32770 vdd.n22401 vdd.n22400 62.202
R32771 vdd.n22208 vdd.n22207 62.202
R32772 vdd.n24346 vdd.n24345 62.202
R32773 vdd.n22072 vdd.n22071 62.202
R32774 vdd.n24229 vdd.n24228 62.202
R32775 vdd.n10473 vdd.n10271 61.933
R32776 vdd.n14527 vdd.n8212 61.74
R32777 vdd.n13107 vdd.n13087 61.74
R32778 vdd.n19298 vdd.n19297 61.74
R32779 vdd.n19968 vdd.n19967 61.74
R32780 vdd.n11600 vdd.n11598 61.667
R32781 vdd.n11600 vdd.n11599 61.667
R32782 vdd.n19331 vdd.n19330 61.574
R32783 vdd.n20540 vdd.n20539 61.574
R32784 vdd.n30499 vdd.n30497 60.14
R32785 vdd.n14970 vdd.n7986 60.14
R32786 vdd.n14529 vdd.n8210 60.14
R32787 vdd.n24489 vdd.n24487 60.14
R32788 vdd.n30350 vdd.n30348 60.139
R32789 vdd.n14948 vdd.n7989 60.139
R32790 vdd.n14506 vdd.n8199 60.139
R32791 vdd.n20518 vdd.n20514 60.139
R32792 vdd.n24414 vdd.n24412 60.139
R32793 vdd.n14599 vdd.n14575 59.481
R32794 vdd.n14973 vdd.n14972 59.481
R32795 vdd.n20025 vdd.n20024 59.481
R32796 vdd.n24672 vdd.n24671 59.481
R32797 vdd.n25090 vdd.n25089 59.481
R32798 vdd.n20511 vdd.n20472 58.641
R32799 vdd.n20060 vdd.n20059 58.641
R32800 vdd.n14969 vdd.n7987 58.497
R32801 vdd.n24156 vdd.n24155 56.547
R32802 vdd.n24018 vdd.n24017 56.547
R32803 vdd.n23924 vdd.n23923 56.547
R32804 vdd.n23786 vdd.n23785 56.547
R32805 vdd.n23692 vdd.n23691 56.547
R32806 vdd.n23098 vdd.n23097 56.547
R32807 vdd.n23236 vdd.n23235 56.547
R32808 vdd.n23330 vdd.n23329 56.547
R32809 vdd.n23468 vdd.n23467 56.547
R32810 vdd.n23562 vdd.n23561 56.547
R32811 vdd.n22519 vdd.n22518 56.547
R32812 vdd.n22657 vdd.n22656 56.547
R32813 vdd.n22751 vdd.n22750 56.547
R32814 vdd.n22889 vdd.n22888 56.547
R32815 vdd.n22983 vdd.n22982 56.547
R32816 vdd.n22430 vdd.n22429 56.547
R32817 vdd.n22286 vdd.n22285 56.547
R32818 vdd.n24258 vdd.n24257 56.547
R32819 vdd.n24196 vdd.n24195 56.47
R32820 vdd.n23974 vdd.n23973 56.47
R32821 vdd.n23964 vdd.n23963 56.47
R32822 vdd.n23742 vdd.n23741 56.47
R32823 vdd.n23732 vdd.n23731 56.47
R32824 vdd.n23054 vdd.n23053 56.47
R32825 vdd.n23276 vdd.n23275 56.47
R32826 vdd.n23286 vdd.n23285 56.47
R32827 vdd.n23508 vdd.n23507 56.47
R32828 vdd.n23518 vdd.n23517 56.47
R32829 vdd.n22475 vdd.n22474 56.47
R32830 vdd.n22697 vdd.n22696 56.47
R32831 vdd.n22707 vdd.n22706 56.47
R32832 vdd.n22929 vdd.n22928 56.47
R32833 vdd.n22939 vdd.n22938 56.47
R32834 vdd.n22179 vdd.n22178 56.47
R32835 vdd.n22261 vdd.n22260 56.47
R32836 vdd.n22273 vdd.n22272 56.47
R32837 vdd.n22146 vdd.n22145 56.47
R32838 vdd.n22158 vdd.n22157 56.47
R32839 vdd.n24102 vdd.n24098 52.941
R32840 vdd.n24076 vdd.n24072 52.941
R32841 vdd.n23870 vdd.n23866 52.941
R32842 vdd.n23844 vdd.n23840 52.941
R32843 vdd.n23638 vdd.n23634 52.941
R32844 vdd.n23156 vdd.n23152 52.941
R32845 vdd.n23182 vdd.n23178 52.941
R32846 vdd.n23388 vdd.n23384 52.941
R32847 vdd.n23414 vdd.n23410 52.941
R32848 vdd.n23620 vdd.n23616 52.941
R32849 vdd.n22577 vdd.n22573 52.941
R32850 vdd.n22603 vdd.n22599 52.941
R32851 vdd.n22809 vdd.n22805 52.941
R32852 vdd.n22835 vdd.n22831 52.941
R32853 vdd.n23041 vdd.n23037 52.941
R32854 vdd.n22193 vdd.n22189 52.941
R32855 vdd.n22200 vdd.n22199 52.941
R32856 vdd.n22051 vdd.n22047 52.941
R32857 vdd.n22058 vdd.n22057 52.941
R32858 vdd.n22172 vdd.n22168 52.941
R32859 vdd.n24143 vdd.n24142 50.892
R32860 vdd.n24033 vdd.n24032 50.892
R32861 vdd.n23911 vdd.n23910 50.892
R32862 vdd.n23801 vdd.n23800 50.892
R32863 vdd.n23679 vdd.n23678 50.892
R32864 vdd.n23113 vdd.n23112 50.892
R32865 vdd.n23223 vdd.n23222 50.892
R32866 vdd.n23345 vdd.n23344 50.892
R32867 vdd.n23455 vdd.n23454 50.892
R32868 vdd.n23577 vdd.n23576 50.892
R32869 vdd.n22534 vdd.n22533 50.892
R32870 vdd.n22644 vdd.n22643 50.892
R32871 vdd.n22766 vdd.n22765 50.892
R32872 vdd.n22876 vdd.n22875 50.892
R32873 vdd.n22998 vdd.n22997 50.892
R32874 vdd.n22416 vdd.n22415 50.892
R32875 vdd.n22225 vdd.n22224 50.892
R32876 vdd.n24361 vdd.n24360 50.892
R32877 vdd.n22101 vdd.n22100 50.892
R32878 vdd.n24244 vdd.n24243 50.892
R32879 vdd.n24182 vdd.n24181 49.411
R32880 vdd.n23988 vdd.n23987 49.411
R32881 vdd.n23950 vdd.n23949 49.411
R32882 vdd.n23756 vdd.n23755 49.411
R32883 vdd.n23718 vdd.n23717 49.411
R32884 vdd.n23068 vdd.n23067 49.411
R32885 vdd.n23262 vdd.n23261 49.411
R32886 vdd.n23300 vdd.n23299 49.411
R32887 vdd.n23494 vdd.n23493 49.411
R32888 vdd.n23532 vdd.n23531 49.411
R32889 vdd.n22489 vdd.n22488 49.411
R32890 vdd.n22683 vdd.n22682 49.411
R32891 vdd.n22721 vdd.n22720 49.411
R32892 vdd.n22915 vdd.n22914 49.411
R32893 vdd.n22953 vdd.n22952 49.411
R32894 vdd.n22459 vdd.n22458 49.411
R32895 vdd.n22336 vdd.n22335 49.411
R32896 vdd.n22315 vdd.n22314 49.411
R32897 vdd.n22138 vdd.n22137 49.411
R32898 vdd.n24287 vdd.n24286 49.411
R32899 vdd.n11739 vdd.n11738 49.396
R32900 vdd.n11823 vdd.n11822 49.396
R32901 vdd.n21818 vdd.n21816 49.396
R32902 vdd.n21914 vdd.n21913 49.396
R32903 vdd.n30493 vdd.n30492 49.094
R32904 vdd.n30490 vdd.n30489 49.094
R32905 vdd.n30474 vdd.n30473 49.094
R32906 vdd.n30469 vdd.n30468 49.094
R32907 vdd.n30462 vdd.n30461 49.094
R32908 vdd.n30456 vdd.n30455 49.094
R32909 vdd.n30447 vdd.n30446 49.094
R32910 vdd.n30442 vdd.n30441 49.094
R32911 vdd.n30438 vdd.n30437 49.094
R32912 vdd.n30429 vdd.n30428 49.094
R32913 vdd.n30420 vdd.n30419 49.094
R32914 vdd.n30415 vdd.n30414 49.094
R32915 vdd.n30411 vdd.n30410 49.094
R32916 vdd.n30405 vdd.n30404 49.094
R32917 vdd.n30400 vdd.n30399 49.094
R32918 vdd.n30396 vdd.n30395 49.094
R32919 vdd.n30391 vdd.n30390 49.094
R32920 vdd.n30372 vdd.n30371 49.094
R32921 vdd.n30363 vdd.n30362 49.094
R32922 vdd.n30354 vdd.n30353 49.094
R32923 vdd.n30354 vdd.n30352 49.094
R32924 vdd.n30356 vdd.n30355 49.094
R32925 vdd.n30358 vdd.n30357 49.094
R32926 vdd.n30363 vdd.n30361 49.094
R32927 vdd.n30366 vdd.n30365 49.094
R32928 vdd.n30372 vdd.n30369 49.094
R32929 vdd.n30375 vdd.n30374 49.094
R32930 vdd.n30378 vdd.n30377 49.094
R32931 vdd.n30381 vdd.n30380 49.094
R32932 vdd.n30384 vdd.n30383 49.094
R32933 vdd.n30387 vdd.n30386 49.094
R32934 vdd.n30396 vdd.n30393 49.094
R32935 vdd.n30405 vdd.n30402 49.094
R32936 vdd.n30411 vdd.n30408 49.094
R32937 vdd.n30420 vdd.n30417 49.094
R32938 vdd.n30423 vdd.n30422 49.094
R32939 vdd.n30429 vdd.n30426 49.094
R32940 vdd.n30432 vdd.n30431 49.094
R32941 vdd.n30438 vdd.n30435 49.094
R32942 vdd.n30447 vdd.n30444 49.094
R32943 vdd.n30450 vdd.n30449 49.094
R32944 vdd.n30456 vdd.n30453 49.094
R32945 vdd.n30462 vdd.n30459 49.094
R32946 vdd.n30465 vdd.n30464 49.094
R32947 vdd.n30474 vdd.n30471 49.094
R32948 vdd.n30477 vdd.n30476 49.094
R32949 vdd.n30480 vdd.n30479 49.094
R32950 vdd.n30483 vdd.n30482 49.094
R32951 vdd.n30485 vdd.n30484 49.094
R32952 vdd.n30487 vdd.n30486 49.094
R32953 vdd.n30493 vdd.n30491 49.094
R32954 vdd.n30495 vdd.n30494 49.094
R32955 vdd.n14524 vdd.n8209 49.094
R32956 vdd.n14522 vdd.n8208 49.094
R32957 vdd.n14520 vdd.n8207 49.094
R32958 vdd.n14518 vdd.n8206 49.094
R32959 vdd.n14516 vdd.n8205 49.094
R32960 vdd.n14514 vdd.n8204 49.094
R32961 vdd.n14512 vdd.n8203 49.094
R32962 vdd.n14510 vdd.n8202 49.094
R32963 vdd.n14508 vdd.n8201 49.094
R32964 vdd.n14506 vdd.n8200 49.094
R32965 vdd.n14968 vdd.n14967 49.094
R32966 vdd.n14964 vdd.n7998 49.094
R32967 vdd.n14962 vdd.n7997 49.094
R32968 vdd.n14960 vdd.n7996 49.094
R32969 vdd.n14958 vdd.n7995 49.094
R32970 vdd.n14956 vdd.n7994 49.094
R32971 vdd.n14954 vdd.n7993 49.094
R32972 vdd.n14952 vdd.n7992 49.094
R32973 vdd.n14950 vdd.n7991 49.094
R32974 vdd.n14948 vdd.n7990 49.094
R32975 vdd.n14950 vdd.n7990 49.094
R32976 vdd.n14952 vdd.n7991 49.094
R32977 vdd.n14954 vdd.n7992 49.094
R32978 vdd.n14956 vdd.n7993 49.094
R32979 vdd.n14958 vdd.n7994 49.094
R32980 vdd.n14960 vdd.n7995 49.094
R32981 vdd.n14962 vdd.n7996 49.094
R32982 vdd.n14964 vdd.n7997 49.094
R32983 vdd.n14967 vdd.n7998 49.094
R32984 vdd.n14968 vdd.n7986 49.094
R32985 vdd.n14508 vdd.n8200 49.094
R32986 vdd.n14510 vdd.n8201 49.094
R32987 vdd.n14512 vdd.n8202 49.094
R32988 vdd.n14514 vdd.n8203 49.094
R32989 vdd.n14516 vdd.n8204 49.094
R32990 vdd.n14518 vdd.n8205 49.094
R32991 vdd.n14520 vdd.n8206 49.094
R32992 vdd.n14522 vdd.n8207 49.094
R32993 vdd.n14524 vdd.n8208 49.094
R32994 vdd.n8210 vdd.n8209 49.094
R32995 vdd.n20536 vdd.n20535 49.094
R32996 vdd.n20534 vdd.n20533 49.094
R32997 vdd.n20532 vdd.n20531 49.094
R32998 vdd.n20527 vdd.n20526 49.094
R32999 vdd.n20524 vdd.n20523 49.094
R33000 vdd.n20521 vdd.n20520 49.094
R33001 vdd.n20527 vdd.n20525 49.094
R33002 vdd.n20529 vdd.n20528 49.094
R33003 vdd.n24485 vdd.n24484 49.094
R33004 vdd.n24481 vdd.n24480 49.094
R33005 vdd.n24478 vdd.n24477 49.094
R33006 vdd.n24476 vdd.n24475 49.094
R33007 vdd.n24474 vdd.n24473 49.094
R33008 vdd.n24470 vdd.n24469 49.094
R33009 vdd.n24465 vdd.n24464 49.094
R33010 vdd.n24462 vdd.n24461 49.094
R33011 vdd.n24437 vdd.n24436 49.094
R33012 vdd.n24428 vdd.n24427 49.094
R33013 vdd.n24423 vdd.n24422 49.094
R33014 vdd.n24421 vdd.n24420 49.094
R33015 vdd.n24416 vdd.n24415 49.094
R33016 vdd.n24418 vdd.n24417 49.094
R33017 vdd.n24428 vdd.n24425 49.094
R33018 vdd.n24431 vdd.n24430 49.094
R33019 vdd.n24437 vdd.n24434 49.094
R33020 vdd.n24440 vdd.n24439 49.094
R33021 vdd.n24443 vdd.n24442 49.094
R33022 vdd.n24446 vdd.n24445 49.094
R33023 vdd.n24449 vdd.n24448 49.094
R33024 vdd.n24452 vdd.n24451 49.094
R33025 vdd.n24455 vdd.n24454 49.094
R33026 vdd.n24458 vdd.n24457 49.094
R33027 vdd.n24470 vdd.n24467 49.094
R33028 vdd.n24481 vdd.n24479 49.094
R33029 vdd.n24485 vdd.n24483 49.094
R33030 vdd.n24509 vdd.n24504 47.085
R33031 vdd.n24491 vdd.n24490 47.085
R33032 vdd.n24116 vdd.n24112 45.882
R33033 vdd.n24062 vdd.n24058 45.882
R33034 vdd.n23884 vdd.n23880 45.882
R33035 vdd.n23830 vdd.n23826 45.882
R33036 vdd.n23652 vdd.n23648 45.882
R33037 vdd.n23142 vdd.n23138 45.882
R33038 vdd.n23196 vdd.n23192 45.882
R33039 vdd.n23374 vdd.n23370 45.882
R33040 vdd.n23428 vdd.n23424 45.882
R33041 vdd.n23606 vdd.n23602 45.882
R33042 vdd.n22563 vdd.n22559 45.882
R33043 vdd.n22617 vdd.n22613 45.882
R33044 vdd.n22795 vdd.n22791 45.882
R33045 vdd.n22849 vdd.n22845 45.882
R33046 vdd.n23027 vdd.n23023 45.882
R33047 vdd.n22390 vdd.n22386 45.882
R33048 vdd.n22360 vdd.n22354 45.882
R33049 vdd.n24335 vdd.n24331 45.882
R33050 vdd.n22089 vdd.n22083 45.882
R33051 vdd.n24218 vdd.n24214 45.882
R33052 vdd.n24142 vdd.n24141 45.238
R33053 vdd.n24032 vdd.n24031 45.238
R33054 vdd.n23910 vdd.n23909 45.238
R33055 vdd.n23800 vdd.n23799 45.238
R33056 vdd.n23678 vdd.n23677 45.238
R33057 vdd.n23112 vdd.n23111 45.238
R33058 vdd.n23222 vdd.n23221 45.238
R33059 vdd.n23344 vdd.n23343 45.238
R33060 vdd.n23454 vdd.n23453 45.238
R33061 vdd.n23576 vdd.n23575 45.238
R33062 vdd.n22533 vdd.n22532 45.238
R33063 vdd.n22643 vdd.n22642 45.238
R33064 vdd.n22765 vdd.n22764 45.238
R33065 vdd.n22875 vdd.n22874 45.238
R33066 vdd.n22997 vdd.n22996 45.238
R33067 vdd.n22415 vdd.n22414 45.238
R33068 vdd.n22224 vdd.n22223 45.238
R33069 vdd.n24360 vdd.n24359 45.238
R33070 vdd.n22100 vdd.n22099 45.238
R33071 vdd.n24243 vdd.n24242 45.238
R33072 vdd.n10596 vdd.n10585 43.659
R33073 vdd.n10761 vdd.n10758 43.659
R33074 vdd.n12284 vdd.n10918 43.659
R33075 vdd.n11116 vdd.n11094 43.659
R33076 vdd.n12071 vdd.n11269 43.659
R33077 vdd.n11978 vdd.n11427 43.659
R33078 vdd.n10382 vdd.n10340 43.659
R33079 vdd.n12992 vdd.n9416 43.659
R33080 vdd.n12886 vdd.n9611 43.659
R33081 vdd.n12784 vdd.n9777 43.659
R33082 vdd.n12678 vdd.n9971 43.659
R33083 vdd.n12586 vdd.n10120 43.659
R33084 vdd.n24168 vdd.n24167 42.352
R33085 vdd.n24002 vdd.n24001 42.352
R33086 vdd.n23936 vdd.n23935 42.352
R33087 vdd.n23770 vdd.n23769 42.352
R33088 vdd.n23704 vdd.n23703 42.352
R33089 vdd.n23082 vdd.n23081 42.352
R33090 vdd.n23248 vdd.n23247 42.352
R33091 vdd.n23314 vdd.n23313 42.352
R33092 vdd.n23480 vdd.n23479 42.352
R33093 vdd.n23546 vdd.n23545 42.352
R33094 vdd.n22503 vdd.n22502 42.352
R33095 vdd.n22669 vdd.n22668 42.352
R33096 vdd.n22735 vdd.n22734 42.352
R33097 vdd.n22901 vdd.n22900 42.352
R33098 vdd.n22967 vdd.n22966 42.352
R33099 vdd.n22443 vdd.n22442 42.352
R33100 vdd.n22247 vdd.n22246 42.352
R33101 vdd.n22299 vdd.n22298 42.352
R33102 vdd.n22123 vdd.n22122 42.352
R33103 vdd.n24271 vdd.n24270 42.352
R33104 vdd.n30500 vdd.n30499 41.621
R33105 vdd.n14970 vdd.n14969 41.621
R33106 vdd.n14530 vdd.n14529 41.621
R33107 vdd.n20539 vdd.n20538 41.621
R33108 vdd.n24490 vdd.n24489 41.621
R33109 vdd.n30500 vdd.n30350 41.621
R33110 vdd.n14969 vdd.n7989 41.621
R33111 vdd.n14530 vdd.n8199 41.621
R33112 vdd.n20539 vdd.n20518 41.621
R33113 vdd.n24490 vdd.n24414 41.621
R33114 vdd.n24509 vdd.n24506 41.621
R33115 vdd.n24509 vdd.n24508 41.621
R33116 vdd.n24157 vdd.n24156 39.583
R33117 vdd.n24019 vdd.n24018 39.583
R33118 vdd.n23925 vdd.n23924 39.583
R33119 vdd.n23787 vdd.n23786 39.583
R33120 vdd.n23693 vdd.n23692 39.583
R33121 vdd.n23099 vdd.n23098 39.583
R33122 vdd.n23237 vdd.n23236 39.583
R33123 vdd.n23331 vdd.n23330 39.583
R33124 vdd.n23469 vdd.n23468 39.583
R33125 vdd.n23563 vdd.n23562 39.583
R33126 vdd.n22520 vdd.n22519 39.583
R33127 vdd.n22658 vdd.n22657 39.583
R33128 vdd.n22752 vdd.n22751 39.583
R33129 vdd.n22890 vdd.n22889 39.583
R33130 vdd.n22984 vdd.n22983 39.583
R33131 vdd.n22431 vdd.n22430 39.583
R33132 vdd.n22233 vdd.n22232 39.583
R33133 vdd.n22287 vdd.n22286 39.583
R33134 vdd.n22109 vdd.n22108 39.583
R33135 vdd.n24259 vdd.n24258 39.583
R33136 vdd.n24838 vdd.t203 39.534
R33137 vdd.t297 vdd.n8113 39.193
R33138 vdd.t293 vdd.n14875 39.193
R33139 vdd.n24130 vdd.n24126 38.823
R33140 vdd.n24048 vdd.n24044 38.823
R33141 vdd.n23898 vdd.n23894 38.823
R33142 vdd.n23816 vdd.n23812 38.823
R33143 vdd.n23666 vdd.n23662 38.823
R33144 vdd.n23128 vdd.n23124 38.823
R33145 vdd.n23210 vdd.n23206 38.823
R33146 vdd.n23360 vdd.n23356 38.823
R33147 vdd.n23442 vdd.n23438 38.823
R33148 vdd.n23592 vdd.n23588 38.823
R33149 vdd.n22549 vdd.n22545 38.823
R33150 vdd.n22631 vdd.n22627 38.823
R33151 vdd.n22781 vdd.n22777 38.823
R33152 vdd.n22863 vdd.n22859 38.823
R33153 vdd.n23013 vdd.n23009 38.823
R33154 vdd.n22402 vdd.n22398 38.823
R33155 vdd.n22210 vdd.n22209 38.823
R33156 vdd.n24347 vdd.n24343 38.823
R33157 vdd.n22074 vdd.n22073 38.823
R33158 vdd.n24230 vdd.n24226 38.823
R33159 vdd.n14601 vdd.n14574 38.799
R33160 vdd.n14596 vdd.n14573 38.799
R33161 vdd.n14593 vdd.n14572 38.799
R33162 vdd.n14589 vdd.n14571 38.799
R33163 vdd.n14585 vdd.n14570 38.799
R33164 vdd.n14581 vdd.n14569 38.799
R33165 vdd.n14577 vdd.n14568 38.799
R33166 vdd.n13109 vdd.n9283 38.799
R33167 vdd.n13104 vdd.n9282 38.799
R33168 vdd.n13101 vdd.n9281 38.799
R33169 vdd.n13097 vdd.n9280 38.799
R33170 vdd.n13093 vdd.n9279 38.799
R33171 vdd.n13089 vdd.n9278 38.799
R33172 vdd.n13112 vdd.n13111 38.799
R33173 vdd.n14643 vdd.n8167 38.799
R33174 vdd.n14638 vdd.n8166 38.799
R33175 vdd.n14635 vdd.n8165 38.799
R33176 vdd.n14631 vdd.n8164 38.799
R33177 vdd.n14627 vdd.n8163 38.799
R33178 vdd.n14623 vdd.n8162 38.799
R33179 vdd.n14619 vdd.n8161 38.799
R33180 vdd.n11657 vdd.n11656 38.799
R33181 vdd.n18491 vdd.n18490 38.799
R33182 vdd.n18489 vdd.n18487 38.799
R33183 vdd.n18486 vdd.n18484 38.799
R33184 vdd.n18483 vdd.n18481 38.799
R33185 vdd.n18480 vdd.n18477 38.799
R33186 vdd.n18475 vdd.n18472 38.799
R33187 vdd.n18470 vdd.n18467 38.799
R33188 vdd.n21738 vdd.n21737 38.799
R33189 vdd.n19329 vdd.n19328 38.799
R33190 vdd.n19327 vdd.n19325 38.799
R33191 vdd.n19324 vdd.n19322 38.799
R33192 vdd.n19321 vdd.n19319 38.799
R33193 vdd.n19318 vdd.n19315 38.799
R33194 vdd.n19313 vdd.n19310 38.799
R33195 vdd.n19308 vdd.n19305 38.799
R33196 vdd.n20510 vdd.n20507 38.799
R33197 vdd.n20505 vdd.n20502 38.799
R33198 vdd.n20500 vdd.n20497 38.799
R33199 vdd.n20495 vdd.n20492 38.799
R33200 vdd.n20490 vdd.n20487 38.799
R33201 vdd.n20485 vdd.n20482 38.799
R33202 vdd.n20480 vdd.n20474 38.799
R33203 vdd.n14594 vdd.n14573 38.798
R33204 vdd.n14590 vdd.n14572 38.798
R33205 vdd.n14586 vdd.n14571 38.798
R33206 vdd.n14582 vdd.n14570 38.798
R33207 vdd.n14578 vdd.n14569 38.798
R33208 vdd.n14568 vdd.n8144 38.798
R33209 vdd.n14601 vdd.n14600 38.798
R33210 vdd.n13102 vdd.n9282 38.798
R33211 vdd.n13098 vdd.n9281 38.798
R33212 vdd.n13094 vdd.n9280 38.798
R33213 vdd.n13090 vdd.n9279 38.798
R33214 vdd.n9278 vdd.n9275 38.798
R33215 vdd.n13111 vdd.n9273 38.798
R33216 vdd.n13109 vdd.n13108 38.798
R33217 vdd.n14636 vdd.n8166 38.798
R33218 vdd.n14632 vdd.n8165 38.798
R33219 vdd.n14628 vdd.n8164 38.798
R33220 vdd.n14624 vdd.n8163 38.798
R33221 vdd.n14620 vdd.n8162 38.798
R33222 vdd.n14616 vdd.n8161 38.798
R33223 vdd.n14643 vdd.n14642 38.798
R33224 vdd.n18489 vdd.n18488 38.798
R33225 vdd.n18486 vdd.n18485 38.798
R33226 vdd.n18483 vdd.n18482 38.798
R33227 vdd.n18480 vdd.n18479 38.798
R33228 vdd.n18475 vdd.n18474 38.798
R33229 vdd.n18470 vdd.n18469 38.798
R33230 vdd.n19327 vdd.n19326 38.798
R33231 vdd.n19324 vdd.n19323 38.798
R33232 vdd.n19321 vdd.n19320 38.798
R33233 vdd.n19318 vdd.n19317 38.798
R33234 vdd.n19313 vdd.n19312 38.798
R33235 vdd.n19308 vdd.n19307 38.798
R33236 vdd.n20505 vdd.n20504 38.798
R33237 vdd.n20500 vdd.n20499 38.798
R33238 vdd.n20495 vdd.n20494 38.798
R33239 vdd.n20490 vdd.n20489 38.798
R33240 vdd.n20485 vdd.n20484 38.798
R33241 vdd.n20480 vdd.n20479 38.798
R33242 vdd.n20510 vdd.n20509 38.798
R33243 vdd.n11657 vdd.n11574 38.798
R33244 vdd.n21738 vdd.n21736 38.798
R33245 vdd.n35713 vdd.n35711 38.798
R33246 vdd.n35839 vdd.n35837 38.798
R33247 vdd.n35836 vdd.n35834 38.798
R33248 vdd.n35832 vdd.n35829 38.798
R33249 vdd.n35827 vdd.n35824 38.798
R33250 vdd.n35822 vdd.n35819 38.798
R33251 vdd.n35817 vdd.n35814 38.798
R33252 vdd.n35812 vdd.n35809 38.798
R33253 vdd.n35807 vdd.n35804 38.798
R33254 vdd.n35802 vdd.n35799 38.798
R33255 vdd.n35797 vdd.n35794 38.798
R33256 vdd.n35792 vdd.n35789 38.798
R33257 vdd.n35787 vdd.n35784 38.798
R33258 vdd.n35782 vdd.n35779 38.798
R33259 vdd.n35777 vdd.n35774 38.798
R33260 vdd.n35772 vdd.n35769 38.798
R33261 vdd.n35767 vdd.n35764 38.798
R33262 vdd.n35762 vdd.n35759 38.798
R33263 vdd.n35757 vdd.n35754 38.798
R33264 vdd.n35752 vdd.n35749 38.798
R33265 vdd.n35747 vdd.n35744 38.798
R33266 vdd.n35742 vdd.n35739 38.798
R33267 vdd.n35737 vdd.n35734 38.798
R33268 vdd.n35732 vdd.n35729 38.798
R33269 vdd.n35727 vdd.n35724 38.798
R33270 vdd.n35722 vdd.n35720 38.798
R33271 vdd.n35719 vdd.n35717 38.798
R33272 vdd.n35716 vdd.n35714 38.798
R33273 vdd.n35713 vdd.n35712 38.798
R33274 vdd.n35839 vdd.n35838 38.798
R33275 vdd.n35836 vdd.n35835 38.798
R33276 vdd.n35832 vdd.n35831 38.798
R33277 vdd.n35827 vdd.n35826 38.798
R33278 vdd.n35822 vdd.n35821 38.798
R33279 vdd.n35817 vdd.n35816 38.798
R33280 vdd.n35812 vdd.n35811 38.798
R33281 vdd.n35807 vdd.n35806 38.798
R33282 vdd.n35802 vdd.n35801 38.798
R33283 vdd.n35797 vdd.n35796 38.798
R33284 vdd.n35792 vdd.n35791 38.798
R33285 vdd.n35787 vdd.n35786 38.798
R33286 vdd.n35782 vdd.n35781 38.798
R33287 vdd.n35777 vdd.n35776 38.798
R33288 vdd.n35772 vdd.n35771 38.798
R33289 vdd.n35767 vdd.n35766 38.798
R33290 vdd.n35762 vdd.n35761 38.798
R33291 vdd.n35757 vdd.n35756 38.798
R33292 vdd.n35752 vdd.n35751 38.798
R33293 vdd.n35747 vdd.n35746 38.798
R33294 vdd.n35742 vdd.n35741 38.798
R33295 vdd.n35737 vdd.n35736 38.798
R33296 vdd.n35732 vdd.n35731 38.798
R33297 vdd.n35727 vdd.n35726 38.798
R33298 vdd.n35722 vdd.n35721 38.798
R33299 vdd.n35719 vdd.n35718 38.798
R33300 vdd.n35716 vdd.n35715 38.798
R33301 vdd.n11650 vdd.n11573 38.798
R33302 vdd.n11646 vdd.n11572 38.798
R33303 vdd.n11642 vdd.n11571 38.798
R33304 vdd.n11638 vdd.n11570 38.798
R33305 vdd.n11634 vdd.n11569 38.798
R33306 vdd.n11630 vdd.n11568 38.798
R33307 vdd.n11652 vdd.n11573 38.798
R33308 vdd.n11649 vdd.n11572 38.798
R33309 vdd.n11645 vdd.n11571 38.798
R33310 vdd.n11641 vdd.n11570 38.798
R33311 vdd.n11637 vdd.n11569 38.798
R33312 vdd.n11633 vdd.n11568 38.798
R33313 vdd.n21735 vdd.n21733 38.798
R33314 vdd.n21732 vdd.n21730 38.798
R33315 vdd.n21729 vdd.n21726 38.798
R33316 vdd.n21724 vdd.n21721 38.798
R33317 vdd.n21719 vdd.n21716 38.798
R33318 vdd.n21714 vdd.n21711 38.798
R33319 vdd.n21735 vdd.n21734 38.798
R33320 vdd.n21732 vdd.n21731 38.798
R33321 vdd.n21729 vdd.n21728 38.798
R33322 vdd.n21724 vdd.n21723 38.798
R33323 vdd.n21719 vdd.n21718 38.798
R33324 vdd.n21714 vdd.n21713 38.798
R33325 vdd.n20037 vdd.n20035 38.798
R33326 vdd.n20040 vdd.n20038 38.798
R33327 vdd.n20043 vdd.n20041 38.798
R33328 vdd.n20048 vdd.n20045 38.798
R33329 vdd.n20053 vdd.n20050 38.798
R33330 vdd.n20058 vdd.n20055 38.798
R33331 vdd.n20058 vdd.n20057 38.798
R33332 vdd.n20053 vdd.n20052 38.798
R33333 vdd.n20048 vdd.n20047 38.798
R33334 vdd.n20043 vdd.n20042 38.798
R33335 vdd.n20040 vdd.n20039 38.798
R33336 vdd.n20037 vdd.n20036 38.798
R33337 vdd.n20034 vdd.n20033 38.798
R33338 vdd.n21741 vdd.n21740 37.55
R33339 vdd.n21616 vdd.n21610 37.296
R33340 vdd.n19147 vdd.n19143 37.296
R33341 vdd.n21009 vdd.n21004 37.296
R33342 vdd.n21668 vdd.n21664 36.592
R33343 vdd.n21673 vdd.n21668 36.592
R33344 vdd.n21398 vdd.n21397 36.592
R33345 vdd.n19032 vdd.n19031 36.592
R33346 vdd.n18773 vdd.n18772 36.592
R33347 vdd.n18514 vdd.n18513 36.592
R33348 vdd.n24154 vdd.n24153 35.294
R33349 vdd.n24016 vdd.n24015 35.294
R33350 vdd.n23922 vdd.n23921 35.294
R33351 vdd.n23784 vdd.n23783 35.294
R33352 vdd.n23690 vdd.n23689 35.294
R33353 vdd.n23096 vdd.n23095 35.294
R33354 vdd.n23234 vdd.n23233 35.294
R33355 vdd.n23328 vdd.n23327 35.294
R33356 vdd.n23466 vdd.n23465 35.294
R33357 vdd.n23560 vdd.n23559 35.294
R33358 vdd.n22517 vdd.n22516 35.294
R33359 vdd.n22655 vdd.n22654 35.294
R33360 vdd.n22749 vdd.n22748 35.294
R33361 vdd.n22887 vdd.n22886 35.294
R33362 vdd.n22981 vdd.n22980 35.294
R33363 vdd.n22428 vdd.n22427 35.294
R33364 vdd.n22236 vdd.n22235 35.294
R33365 vdd.n22284 vdd.n22283 35.294
R33366 vdd.n22112 vdd.n22111 35.294
R33367 vdd.n24256 vdd.n24255 35.294
R33368 vdd.n24128 vdd.n24127 33.928
R33369 vdd.n24046 vdd.n24045 33.928
R33370 vdd.n23896 vdd.n23895 33.928
R33371 vdd.n23814 vdd.n23813 33.928
R33372 vdd.n23664 vdd.n23663 33.928
R33373 vdd.n23126 vdd.n23125 33.928
R33374 vdd.n23208 vdd.n23207 33.928
R33375 vdd.n23358 vdd.n23357 33.928
R33376 vdd.n23440 vdd.n23439 33.928
R33377 vdd.n23590 vdd.n23589 33.928
R33378 vdd.n22547 vdd.n22546 33.928
R33379 vdd.n22629 vdd.n22628 33.928
R33380 vdd.n22779 vdd.n22778 33.928
R33381 vdd.n22861 vdd.n22860 33.928
R33382 vdd.n23011 vdd.n23010 33.928
R33383 vdd.n22400 vdd.n22399 33.928
R33384 vdd.n24345 vdd.n24344 33.928
R33385 vdd.n24228 vdd.n24227 33.928
R33386 vdd.n11658 vdd.n11567 32.306
R33387 vdd.n24144 vdd.n24140 31.764
R33388 vdd.n24034 vdd.n24030 31.764
R33389 vdd.n23912 vdd.n23908 31.764
R33390 vdd.n23802 vdd.n23798 31.764
R33391 vdd.n23680 vdd.n23676 31.764
R33392 vdd.n23114 vdd.n23110 31.764
R33393 vdd.n23224 vdd.n23220 31.764
R33394 vdd.n23346 vdd.n23342 31.764
R33395 vdd.n23456 vdd.n23452 31.764
R33396 vdd.n23578 vdd.n23574 31.764
R33397 vdd.n22535 vdd.n22531 31.764
R33398 vdd.n22645 vdd.n22641 31.764
R33399 vdd.n22767 vdd.n22763 31.764
R33400 vdd.n22877 vdd.n22873 31.764
R33401 vdd.n22999 vdd.n22995 31.764
R33402 vdd.n22417 vdd.n22413 31.764
R33403 vdd.n22226 vdd.n22221 31.764
R33404 vdd.n24362 vdd.n24358 31.764
R33405 vdd.n22102 vdd.n22097 31.764
R33406 vdd.n24245 vdd.n24241 31.764
R33407 vdd.n35912 vdd.n35908 31.448
R33408 vdd.n35933 vdd.n35928 31.448
R33409 vdd.n36143 vdd.n36139 31.448
R33410 vdd.n36164 vdd.n36159 31.448
R33411 vdd.n36374 vdd.n36370 31.448
R33412 vdd.n36395 vdd.n36390 31.448
R33413 vdd.n36605 vdd.n36601 31.448
R33414 vdd.n36626 vdd.n36621 31.448
R33415 vdd.n36836 vdd.n36832 31.448
R33416 vdd.n36857 vdd.n36852 31.448
R33417 vdd.n33267 vdd.n33263 31.448
R33418 vdd.n33249 vdd.n33244 31.448
R33419 vdd.n33073 vdd.n33069 31.448
R33420 vdd.n37259 vdd.n37254 31.448
R33421 vdd.n37445 vdd.n37440 31.448
R33422 vdd.n32913 vdd.n32909 31.448
R33423 vdd.n38124 vdd.n38120 31.448
R33424 vdd.n38135 vdd.n38130 31.448
R33425 vdd.n37912 vdd.n37907 31.448
R33426 vdd.n37891 vdd.n37887 31.448
R33427 vdd.n37681 vdd.n37676 31.448
R33428 vdd.n37660 vdd.n37656 31.448
R33429 vdd.n28333 vdd.n28329 31.448
R33430 vdd.n28354 vdd.n28349 31.448
R33431 vdd.n28564 vdd.n28560 31.448
R33432 vdd.n28585 vdd.n28580 31.448
R33433 vdd.n28795 vdd.n28791 31.448
R33434 vdd.n28152 vdd.n28147 31.448
R33435 vdd.n27767 vdd.n27762 31.448
R33436 vdd.n31890 vdd.n31889 31.448
R33437 vdd.n32228 vdd.n32227 31.448
R33438 vdd.n29693 vdd.n29688 31.448
R33439 vdd.n30299 vdd.n30294 31.448
R33440 vdd.n30567 vdd.n30563 31.448
R33441 vdd.n2792 vdd.n2791 31.448
R33442 vdd.n2809 vdd.n2808 31.448
R33443 vdd.n2973 vdd.n2972 31.448
R33444 vdd.n2990 vdd.n2989 31.448
R33445 vdd.n3154 vdd.n3153 31.448
R33446 vdd.n3171 vdd.n3170 31.448
R33447 vdd.n3335 vdd.n3334 31.448
R33448 vdd.n3352 vdd.n3351 31.448
R33449 vdd.n3516 vdd.n3515 31.448
R33450 vdd.n3533 vdd.n3532 31.448
R33451 vdd.n3709 vdd.n3708 31.448
R33452 vdd.n4010 vdd.n4009 31.448
R33453 vdd.n2282 vdd.n2281 31.448
R33454 vdd.n2301 vdd.n2300 31.448
R33455 vdd.n1978 vdd.n1977 31.448
R33456 vdd.n1988 vdd.n1987 31.448
R33457 vdd.n1738 vdd.n1737 31.448
R33458 vdd.n1745 vdd.n1744 31.448
R33459 vdd.n1571 vdd.n1570 31.448
R33460 vdd.n1554 vdd.n1553 31.448
R33461 vdd.n1390 vdd.n1389 31.448
R33462 vdd.n1373 vdd.n1372 31.448
R33463 vdd.n26839 vdd.n26838 31.448
R33464 vdd.n26856 vdd.n26855 31.448
R33465 vdd.n27020 vdd.n27019 31.448
R33466 vdd.n27037 vdd.n27036 31.448
R33467 vdd.n27201 vdd.n27200 31.448
R33468 vdd.n26744 vdd.n26743 31.448
R33469 vdd.n31866 vdd.n31865 31.448
R33470 vdd.n31892 vdd.n31885 31.448
R33471 vdd.n32230 vdd.n32223 31.448
R33472 vdd.n32257 vdd.n32256 31.448
R33473 vdd.n31118 vdd.n31117 31.448
R33474 vdd.n31178 vdd.n31177 31.448
R33475 vdd.n13215 vdd.n9171 31.448
R33476 vdd.n9177 vdd.n9172 31.448
R33477 vdd.n13508 vdd.n8951 31.448
R33478 vdd.n8956 vdd.n8952 31.448
R33479 vdd.n8768 vdd.n8732 31.448
R33480 vdd.n8737 vdd.n8733 31.448
R33481 vdd.n14117 vdd.n8514 31.448
R33482 vdd.n14109 vdd.n8506 31.448
R33483 vdd.n14397 vdd.n8298 31.448
R33484 vdd.n14429 vdd.n8275 31.448
R33485 vdd.n14786 vdd.n8075 31.448
R33486 vdd.n14782 vdd.n8079 31.448
R33487 vdd.n11627 vdd.n11578 31.448
R33488 vdd.n13144 vdd.n9246 31.448
R33489 vdd.n13380 vdd.n9057 31.448
R33490 vdd.n13437 vdd.n9022 31.448
R33491 vdd.n13672 vdd.n8837 31.448
R33492 vdd.n13729 vdd.n8802 31.448
R33493 vdd.n13951 vdd.n8595 31.448
R33494 vdd.n13994 vdd.n8596 31.448
R33495 vdd.n14241 vdd.n8373 31.448
R33496 vdd.n14285 vdd.n8374 31.448
R33497 vdd.n14604 vdd.n8180 31.448
R33498 vdd.n14613 vdd.n8175 31.448
R33499 vdd.n19419 vdd.n19410 31.448
R33500 vdd.n19433 vdd.n19427 31.448
R33501 vdd.n19622 vdd.n19613 31.448
R33502 vdd.n19636 vdd.n19630 31.448
R33503 vdd.n19824 vdd.n19815 31.448
R33504 vdd.n19171 vdd.n19165 31.448
R33505 vdd.n20844 vdd.n20835 31.448
R33506 vdd.n20827 vdd.n20821 31.448
R33507 vdd.n20642 vdd.n20633 31.448
R33508 vdd.n20625 vdd.n20619 31.448
R33509 vdd.n21663 vdd.n21662 31.448
R33510 vdd.n21674 vdd.n21657 31.448
R33511 vdd.n21399 vdd.n21390 31.448
R33512 vdd.n21382 vdd.n21376 31.448
R33513 vdd.n21140 vdd.n21131 31.448
R33514 vdd.n21123 vdd.n21117 31.448
R33515 vdd.n19033 vdd.n19024 31.448
R33516 vdd.n19016 vdd.n19010 31.448
R33517 vdd.n18774 vdd.n18765 31.448
R33518 vdd.n18757 vdd.n18751 31.448
R33519 vdd.n18515 vdd.n18506 31.448
R33520 vdd.n18498 vdd.n18465 31.448
R33521 vdd.n19993 vdd.n19992 31.448
R33522 vdd.n20005 vdd.n20004 31.448
R33523 vdd.n24511 vdd.n24510 31.448
R33524 vdd.n20470 vdd.n19978 31.08
R33525 vdd.n20404 vdd.n20403 31.08
R33526 vdd.n20381 vdd.n20376 31.08
R33527 vdd.n20168 vdd.n20167 31.08
R33528 vdd.n20145 vdd.n20140 31.08
R33529 vdd.n14674 vdd.n8124 31.003
R33530 vdd.n14685 vdd.n8125 31.003
R33531 vdd.n14702 vdd.n8119 31.003
R33532 vdd.n14712 vdd.n8113 31.003
R33533 vdd.n14714 vdd.n8104 31.003
R33534 vdd.n14729 vdd.n8100 31.003
R33535 vdd.n14758 vdd.n8094 31.003
R33536 vdd.n14760 vdd.n8082 31.003
R33537 vdd.n14789 vdd.n14788 31.003
R33538 vdd.n14800 vdd.n8064 31.003
R33539 vdd.n14818 vdd.n8055 31.003
R33540 vdd.n14816 vdd.n8050 31.003
R33541 vdd.n14844 vdd.n8044 31.003
R33542 vdd.n14859 vdd.n8035 31.003
R33543 vdd.n14875 vdd.n8030 31.003
R33544 vdd.n14876 vdd.n8020 31.003
R33545 vdd.n14896 vdd.n8021 31.003
R33546 vdd.n14894 vdd.n8016 31.003
R33547 vdd.n14932 vdd.n14927 31.003
R33548 vdd.n14930 vdd.n8001 31.003
R33549 vdd.n19621 vdd.n19620 30.493
R33550 vdd.n19823 vdd.n19822 30.493
R33551 vdd.n20843 vdd.n20842 30.493
R33552 vdd.n20641 vdd.n20640 30.493
R33553 vdd.n30499 vdd.n30498 30.07
R33554 vdd.n14971 vdd.n14970 30.07
R33555 vdd.n14529 vdd.n14528 30.07
R33556 vdd.n24489 vdd.n24488 30.07
R33557 vdd.n30350 vdd.n30349 30.07
R33558 vdd.n14504 vdd.n8199 30.07
R33559 vdd.n14946 vdd.n7989 30.07
R33560 vdd.n20518 vdd.n20517 30.07
R33561 vdd.n24414 vdd.n24413 30.07
R33562 vdd.n24508 vdd.n24507 30.07
R33563 vdd.n24506 vdd.n24505 30.07
R33564 vdd.t307 vdd.n8105 29.833
R33565 vdd.t292 vdd.n8034 29.833
R33566 vdd.n36027 vdd.n36026 29.482
R33567 vdd.n36041 vdd.n36040 29.482
R33568 vdd.n36258 vdd.n36257 29.482
R33569 vdd.n36272 vdd.n36271 29.482
R33570 vdd.n36489 vdd.n36488 29.482
R33571 vdd.n36503 vdd.n36502 29.482
R33572 vdd.n36720 vdd.n36719 29.482
R33573 vdd.n36734 vdd.n36733 29.482
R33574 vdd.n36951 vdd.n36950 29.482
R33575 vdd.n36965 vdd.n36964 29.482
R33576 vdd.n33143 vdd.n33142 29.482
R33577 vdd.n35637 vdd.n35636 29.482
R33578 vdd.n37319 vdd.n37318 29.482
R33579 vdd.n37349 vdd.n37348 29.482
R33580 vdd.n35664 vdd.n35663 29.482
R33581 vdd.n32826 vdd.n32825 29.482
R33582 vdd.n38020 vdd.n38019 29.482
R33583 vdd.n38006 vdd.n38005 29.482
R33584 vdd.n37789 vdd.n37788 29.482
R33585 vdd.n37775 vdd.n37774 29.482
R33586 vdd.n28217 vdd.n28216 29.482
R33587 vdd.n28231 vdd.n28230 29.482
R33588 vdd.n28448 vdd.n28447 29.482
R33589 vdd.n28462 vdd.n28461 29.482
R33590 vdd.n28679 vdd.n28678 29.482
R33591 vdd.n28693 vdd.n28692 29.482
R33592 vdd.n26699 vdd.n26698 29.482
R33593 vdd.n26308 vdd.n26307 29.482
R33594 vdd.n27981 vdd.n27980 29.482
R33595 vdd.n27878 vdd.n27877 29.482
R33596 vdd.n31458 vdd.n31457 29.482
R33597 vdd.n32401 vdd.n32400 29.482
R33598 vdd.n2885 vdd.n2884 29.482
R33599 vdd.n2895 vdd.n2894 29.482
R33600 vdd.n3066 vdd.n3065 29.482
R33601 vdd.n3076 vdd.n3075 29.482
R33602 vdd.n3247 vdd.n3246 29.482
R33603 vdd.n3257 vdd.n3256 29.482
R33604 vdd.n3428 vdd.n3427 29.482
R33605 vdd.n3438 vdd.n3437 29.482
R33606 vdd.n3609 vdd.n3608 29.482
R33607 vdd.n3619 vdd.n3618 29.482
R33608 vdd.n3896 vdd.n3895 29.482
R33609 vdd.n3813 vdd.n3812 29.482
R33610 vdd.n2524 vdd.n2523 29.482
R33611 vdd.n2494 vdd.n2493 29.482
R33612 vdd.n1239 vdd.n1238 29.482
R33613 vdd.n1815 vdd.n1814 29.482
R33614 vdd.n1657 vdd.n1656 29.482
R33615 vdd.n1647 vdd.n1646 29.482
R33616 vdd.n1476 vdd.n1475 29.482
R33617 vdd.n1466 vdd.n1465 29.482
R33618 vdd.n1295 vdd.n1294 29.482
R33619 vdd.n26761 vdd.n26760 29.482
R33620 vdd.n26932 vdd.n26931 29.482
R33621 vdd.n26942 vdd.n26941 29.482
R33622 vdd.n27113 vdd.n27112 29.482
R33623 vdd.n27123 vdd.n27122 29.482
R33624 vdd.n26695 vdd.n26694 29.482
R33625 vdd.n26304 vdd.n26303 29.482
R33626 vdd.n31613 vdd.n31612 29.482
R33627 vdd.n31597 vdd.n31596 29.482
R33628 vdd.n31454 vdd.n31453 29.482
R33629 vdd.n32397 vdd.n32396 29.482
R33630 vdd.n13358 vdd.n9063 29.482
R33631 vdd.n13403 vdd.n9047 29.482
R33632 vdd.n13650 vdd.n8843 29.482
R33633 vdd.n13696 vdd.n8826 29.482
R33634 vdd.n13966 vdd.n8623 29.482
R33635 vdd.n8628 vdd.n8612 29.482
R33636 vdd.n14256 vdd.n8401 29.482
R33637 vdd.n8406 vdd.n8390 29.482
R33638 vdd.n14683 vdd.n8118 29.482
R33639 vdd.n14711 vdd.n8112 29.482
R33640 vdd.n14857 vdd.n14856 29.482
R33641 vdd.n14905 vdd.n8022 29.482
R33642 vdd.n13244 vdd.n9180 29.482
R33643 vdd.n13277 vdd.n9156 29.482
R33644 vdd.n13536 vdd.n8959 29.482
R33645 vdd.n13569 vdd.n8935 29.482
R33646 vdd.n13819 vdd.n8713 29.482
R33647 vdd.n13857 vdd.n8714 29.482
R33648 vdd.n8527 vdd.n8491 29.482
R33649 vdd.n14146 vdd.n8492 29.482
R33650 vdd.n8296 vdd.n8288 29.482
R33651 vdd.n8289 vdd.n8240 29.482
R33652 vdd.n19262 vdd.n19261 29.482
R33653 vdd.n19250 vdd.n19249 29.482
R33654 vdd.n19206 vdd.n19205 29.482
R33655 vdd.n19194 vdd.n19193 29.482
R33656 vdd.n19848 vdd.n19847 29.482
R33657 vdd.n19860 vdd.n19859 29.482
R33658 vdd.n19916 vdd.n19915 29.482
R33659 vdd.n19928 vdd.n19927 29.482
R33660 vdd.n21523 vdd.n21522 29.482
R33661 vdd.n21505 vdd.n21504 29.482
R33662 vdd.n21264 vdd.n21263 29.482
R33663 vdd.n21246 vdd.n21245 29.482
R33664 vdd.n19145 vdd.n19144 29.482
R33665 vdd.n19137 vdd.n19136 29.482
R33666 vdd.n18898 vdd.n18897 29.482
R33667 vdd.n18880 vdd.n18879 29.482
R33668 vdd.n18639 vdd.n18638 29.482
R33669 vdd.n18621 vdd.n18620 29.482
R33670 vdd.n20405 vdd.n20396 29.482
R33671 vdd.n20382 vdd.n20373 29.482
R33672 vdd.n20169 vdd.n20160 29.482
R33673 vdd.n20146 vdd.n20137 29.482
R33674 vdd.n24742 vdd.n24739 29.482
R33675 vdd.n25174 vdd.n25171 29.482
R33676 vdd.n19418 vdd.t242 28.734
R33677 vdd.n20624 vdd.t248 28.734
R33678 vdd.n24171 vdd.n24170 28.273
R33679 vdd.n24005 vdd.n24004 28.273
R33680 vdd.n23939 vdd.n23938 28.273
R33681 vdd.n23773 vdd.n23772 28.273
R33682 vdd.n23707 vdd.n23706 28.273
R33683 vdd.n23085 vdd.n23084 28.273
R33684 vdd.n23251 vdd.n23250 28.273
R33685 vdd.n23317 vdd.n23316 28.273
R33686 vdd.n23483 vdd.n23482 28.273
R33687 vdd.n23549 vdd.n23548 28.273
R33688 vdd.n22506 vdd.n22505 28.273
R33689 vdd.n22672 vdd.n22671 28.273
R33690 vdd.n22738 vdd.n22737 28.273
R33691 vdd.n22904 vdd.n22903 28.273
R33692 vdd.n22970 vdd.n22969 28.273
R33693 vdd.n22446 vdd.n22445 28.273
R33694 vdd.n22251 vdd.n22250 28.273
R33695 vdd.n22302 vdd.n22301 28.273
R33696 vdd.n22127 vdd.n22126 28.273
R33697 vdd.n24274 vdd.n24273 28.273
R33698 vdd.n24140 vdd.n24139 28.235
R33699 vdd.n24030 vdd.n24029 28.235
R33700 vdd.n23908 vdd.n23907 28.235
R33701 vdd.n23798 vdd.n23797 28.235
R33702 vdd.n23676 vdd.n23675 28.235
R33703 vdd.n23110 vdd.n23109 28.235
R33704 vdd.n23220 vdd.n23219 28.235
R33705 vdd.n23342 vdd.n23341 28.235
R33706 vdd.n23452 vdd.n23451 28.235
R33707 vdd.n23574 vdd.n23573 28.235
R33708 vdd.n22531 vdd.n22530 28.235
R33709 vdd.n22641 vdd.n22640 28.235
R33710 vdd.n22763 vdd.n22762 28.235
R33711 vdd.n22873 vdd.n22872 28.235
R33712 vdd.n22995 vdd.n22994 28.235
R33713 vdd.n22413 vdd.n22412 28.235
R33714 vdd.n22221 vdd.n22220 28.235
R33715 vdd.n24358 vdd.n24357 28.235
R33716 vdd.n22097 vdd.n22096 28.235
R33717 vdd.n24241 vdd.n24240 28.235
R33718 vdd.n24876 vdd.t101 28.21
R33719 vdd.n24865 vdd.t139 28.175
R33720 vdd.n10265 vdd.n10264 27.741
R33721 vdd.n35898 vdd.n35894 27.517
R33722 vdd.n35947 vdd.n35943 27.517
R33723 vdd.n36129 vdd.n36125 27.517
R33724 vdd.n36178 vdd.n36174 27.517
R33725 vdd.n36360 vdd.n36356 27.517
R33726 vdd.n36409 vdd.n36405 27.517
R33727 vdd.n36591 vdd.n36587 27.517
R33728 vdd.n36640 vdd.n36636 27.517
R33729 vdd.n36822 vdd.n36818 27.517
R33730 vdd.n36871 vdd.n36867 27.517
R33731 vdd.n37057 vdd.n37053 27.517
R33732 vdd.n37096 vdd.n37092 27.517
R33733 vdd.n37227 vdd.n37226 27.517
R33734 vdd.n33058 vdd.n33054 27.517
R33735 vdd.n32928 vdd.n32924 27.517
R33736 vdd.n37469 vdd.n37465 27.517
R33737 vdd.n38151 vdd.n38147 27.517
R33738 vdd.n38108 vdd.n38104 27.517
R33739 vdd.n37926 vdd.n37922 27.517
R33740 vdd.n37877 vdd.n37873 27.517
R33741 vdd.n37695 vdd.n37691 27.517
R33742 vdd.n37646 vdd.n37642 27.517
R33743 vdd.n28319 vdd.n28315 27.517
R33744 vdd.n28368 vdd.n28364 27.517
R33745 vdd.n28550 vdd.n28546 27.517
R33746 vdd.n28599 vdd.n28595 27.517
R33747 vdd.n28781 vdd.n28777 27.517
R33748 vdd.n28164 vdd.n28160 27.517
R33749 vdd.n31845 vdd.n31844 27.517
R33750 vdd.n29029 vdd.n29025 27.517
R33751 vdd.n29871 vdd.n29867 27.517
R33752 vdd.n29837 vdd.n29833 27.517
R33753 vdd.n31093 vdd.n31092 27.517
R33754 vdd.n30546 vdd.n30542 27.517
R33755 vdd.n2781 vdd.n2780 27.517
R33756 vdd.n2820 vdd.n2819 27.517
R33757 vdd.n2962 vdd.n2961 27.517
R33758 vdd.n3001 vdd.n3000 27.517
R33759 vdd.n3143 vdd.n3142 27.517
R33760 vdd.n3182 vdd.n3181 27.517
R33761 vdd.n3324 vdd.n3323 27.517
R33762 vdd.n3363 vdd.n3362 27.517
R33763 vdd.n3505 vdd.n3504 27.517
R33764 vdd.n3544 vdd.n3543 27.517
R33765 vdd.n3690 vdd.n3689 27.517
R33766 vdd.n3995 vdd.n3994 27.517
R33767 vdd.n2157 vdd.n2153 27.517
R33768 vdd.n2320 vdd.n2319 27.517
R33769 vdd.n2566 vdd.n2565 27.517
R33770 vdd.n2071 vdd.n2070 27.517
R33771 vdd.n1757 vdd.n1756 27.517
R33772 vdd.n1724 vdd.n1723 27.517
R33773 vdd.n1582 vdd.n1581 27.517
R33774 vdd.n1543 vdd.n1542 27.517
R33775 vdd.n1401 vdd.n1400 27.517
R33776 vdd.n1362 vdd.n1361 27.517
R33777 vdd.n26828 vdd.n26827 27.517
R33778 vdd.n26867 vdd.n26866 27.517
R33779 vdd.n27009 vdd.n27008 27.517
R33780 vdd.n27048 vdd.n27047 27.517
R33781 vdd.n27190 vdd.n27189 27.517
R33782 vdd.n26736 vdd.n26735 27.517
R33783 vdd.n31847 vdd.n31840 27.517
R33784 vdd.n31910 vdd.n31909 27.517
R33785 vdd.n32202 vdd.n32201 27.517
R33786 vdd.n32282 vdd.n32281 27.517
R33787 vdd.n31095 vdd.n31088 27.517
R33788 vdd.n31267 vdd.n31266 27.517
R33789 vdd.n13206 vdd.n9208 27.517
R33790 vdd.n13267 vdd.n9164 27.517
R33791 vdd.n13500 vdd.n8987 27.517
R33792 vdd.n13559 vdd.n8943 27.517
R33793 vdd.n13779 vdd.n8767 27.517
R33794 vdd.n13841 vdd.n8727 27.517
R33795 vdd.n14077 vdd.n8553 27.517
R33796 vdd.n14130 vdd.n14129 27.517
R33797 vdd.n14355 vdd.n8335 27.517
R33798 vdd.n14421 vdd.n8284 27.517
R33799 vdd.n14790 vdd.n8070 27.517
R33800 vdd.n14799 vdd.n8063 27.517
R33801 vdd.n13134 vdd.n9262 27.517
R33802 vdd.n9077 vdd.n9061 27.517
R33803 vdd.n13429 vdd.n9031 27.517
R33804 vdd.n8857 vdd.n8841 27.517
R33805 vdd.n13721 vdd.n8811 27.517
R33806 vdd.n13959 vdd.n8630 27.517
R33807 vdd.n14013 vdd.n8582 27.517
R33808 vdd.n14249 vdd.n8409 27.517
R33809 vdd.n14303 vdd.n8363 27.517
R33810 vdd.n14546 vdd.n14539 27.517
R33811 vdd.n19400 vdd.n19394 27.517
R33812 vdd.n19449 vdd.n19443 27.517
R33813 vdd.n19606 vdd.n19600 27.517
R33814 vdd.n19649 vdd.n19643 27.517
R33815 vdd.n19808 vdd.n19802 27.517
R33816 vdd.n20998 vdd.n19158 27.517
R33817 vdd.n20857 vdd.n20851 27.517
R33818 vdd.n20814 vdd.n20808 27.517
R33819 vdd.n20658 vdd.n20652 27.517
R33820 vdd.n20609 vdd.n20603 27.517
R33821 vdd.n21606 vdd.n21605 27.517
R33822 vdd.n21415 vdd.n21409 27.517
R33823 vdd.n21366 vdd.n21360 27.517
R33824 vdd.n21156 vdd.n21150 27.517
R33825 vdd.n21107 vdd.n21101 27.517
R33826 vdd.n19049 vdd.n19043 27.517
R33827 vdd.n19000 vdd.n18994 27.517
R33828 vdd.n18790 vdd.n18784 27.517
R33829 vdd.n18741 vdd.n18735 27.517
R33830 vdd.n18531 vdd.n18525 27.517
R33831 vdd.n20277 vdd.n20276 27.517
R33832 vdd.n20259 vdd.n20258 27.517
R33833 vdd.n24826 vdd.n24825 27.517
R33834 vdd.n14914 vdd.t300 27.493
R33835 vdd.n14602 vdd.n14573 26.852
R33836 vdd.n14602 vdd.n14572 26.852
R33837 vdd.n14602 vdd.n14571 26.852
R33838 vdd.n14602 vdd.n14570 26.852
R33839 vdd.n14602 vdd.n14569 26.852
R33840 vdd.n14602 vdd.n14568 26.852
R33841 vdd.n14602 vdd.n14601 26.852
R33842 vdd.n13110 vdd.n9282 26.852
R33843 vdd.n13110 vdd.n9281 26.852
R33844 vdd.n13110 vdd.n9280 26.852
R33845 vdd.n13110 vdd.n9279 26.852
R33846 vdd.n13110 vdd.n9278 26.852
R33847 vdd.n13111 vdd.n13110 26.852
R33848 vdd.n13110 vdd.n13109 26.852
R33849 vdd.n14644 vdd.n8166 26.852
R33850 vdd.n14644 vdd.n8165 26.852
R33851 vdd.n14644 vdd.n8164 26.852
R33852 vdd.n14644 vdd.n8163 26.852
R33853 vdd.n14644 vdd.n8162 26.852
R33854 vdd.n14644 vdd.n8161 26.852
R33855 vdd.n14644 vdd.n14643 26.852
R33856 vdd.n18492 vdd.n18489 26.852
R33857 vdd.n18492 vdd.n18486 26.852
R33858 vdd.n18492 vdd.n18483 26.852
R33859 vdd.n18492 vdd.n18480 26.852
R33860 vdd.n18492 vdd.n18475 26.852
R33861 vdd.n18492 vdd.n18470 26.852
R33862 vdd.n18492 vdd.n18491 26.852
R33863 vdd.n19330 vdd.n19327 26.852
R33864 vdd.n19330 vdd.n19324 26.852
R33865 vdd.n19330 vdd.n19321 26.852
R33866 vdd.n19330 vdd.n19318 26.852
R33867 vdd.n19330 vdd.n19313 26.852
R33868 vdd.n19330 vdd.n19308 26.852
R33869 vdd.n19330 vdd.n19329 26.852
R33870 vdd.n20511 vdd.n20505 26.852
R33871 vdd.n20511 vdd.n20500 26.852
R33872 vdd.n20511 vdd.n20495 26.852
R33873 vdd.n20511 vdd.n20490 26.852
R33874 vdd.n20511 vdd.n20485 26.852
R33875 vdd.n20511 vdd.n20480 26.852
R33876 vdd.n20511 vdd.n20510 26.852
R33877 vdd.n11658 vdd.n11657 26.852
R33878 vdd.n21739 vdd.n21738 26.852
R33879 vdd.n35841 vdd.n35839 26.852
R33880 vdd.n35841 vdd.n35836 26.852
R33881 vdd.n35841 vdd.n35832 26.852
R33882 vdd.n35841 vdd.n35827 26.852
R33883 vdd.n35841 vdd.n35822 26.852
R33884 vdd.n35841 vdd.n35817 26.852
R33885 vdd.n35841 vdd.n35812 26.852
R33886 vdd.n35841 vdd.n35807 26.852
R33887 vdd.n35841 vdd.n35802 26.852
R33888 vdd.n35841 vdd.n35797 26.852
R33889 vdd.n35841 vdd.n35792 26.852
R33890 vdd.n35841 vdd.n35787 26.852
R33891 vdd.n35841 vdd.n35782 26.852
R33892 vdd.n35841 vdd.n35777 26.852
R33893 vdd.n35841 vdd.n35772 26.852
R33894 vdd.n35841 vdd.n35767 26.852
R33895 vdd.n35841 vdd.n35762 26.852
R33896 vdd.n35841 vdd.n35757 26.852
R33897 vdd.n35841 vdd.n35752 26.852
R33898 vdd.n35841 vdd.n35747 26.852
R33899 vdd.n35841 vdd.n35742 26.852
R33900 vdd.n35841 vdd.n35737 26.852
R33901 vdd.n35841 vdd.n35732 26.852
R33902 vdd.n35841 vdd.n35727 26.852
R33903 vdd.n35841 vdd.n35722 26.852
R33904 vdd.n35841 vdd.n35719 26.852
R33905 vdd.n35841 vdd.n35716 26.852
R33906 vdd.n35841 vdd.n35713 26.852
R33907 vdd.n11658 vdd.n11573 26.852
R33908 vdd.n11658 vdd.n11572 26.852
R33909 vdd.n11658 vdd.n11571 26.852
R33910 vdd.n11658 vdd.n11570 26.852
R33911 vdd.n11658 vdd.n11569 26.852
R33912 vdd.n11658 vdd.n11568 26.852
R33913 vdd.n21739 vdd.n21735 26.852
R33914 vdd.n21739 vdd.n21732 26.852
R33915 vdd.n21739 vdd.n21729 26.852
R33916 vdd.n21739 vdd.n21724 26.852
R33917 vdd.n21739 vdd.n21719 26.852
R33918 vdd.n21739 vdd.n21714 26.852
R33919 vdd.n20059 vdd.n20053 26.852
R33920 vdd.n20059 vdd.n20048 26.852
R33921 vdd.n20059 vdd.n20043 26.852
R33922 vdd.n20059 vdd.n20040 26.852
R33923 vdd.n20059 vdd.n20037 26.852
R33924 vdd.n20059 vdd.n20034 26.852
R33925 vdd.n20059 vdd.n20058 26.852
R33926 vdd.n21074 vdd.t279 26.037
R33927 vdd.n24504 vdd.n24503 25.614
R33928 vdd.n24503 vdd.n24502 25.614
R33929 vdd.n24502 vdd.n24501 25.614
R33930 vdd.n24501 vdd.n24500 25.614
R33931 vdd.n24500 vdd.n24499 25.614
R33932 vdd.n24498 vdd.n24497 25.614
R33933 vdd.n24497 vdd.n24496 25.614
R33934 vdd.n24496 vdd.n24495 25.614
R33935 vdd.n24495 vdd.n24494 25.614
R33936 vdd.n24494 vdd.n24493 25.614
R33937 vdd.n24493 vdd.n24492 25.614
R33938 vdd.n24492 vdd.n24491 25.614
R33939 vdd.n30331 vdd.n30330 25.6
R33940 vdd.n30330 vdd.n30329 25.6
R33941 vdd.n30329 vdd.n30328 25.6
R33942 vdd.n30328 vdd.n30327 25.6
R33943 vdd.n30327 vdd.n30326 25.6
R33944 vdd.n30326 vdd.n30325 25.6
R33945 vdd.n30325 vdd.n30324 25.6
R33946 vdd.n31134 vdd.n31133 25.6
R33947 vdd.n31135 vdd.n31134 25.6
R33948 vdd.n31136 vdd.n31135 25.6
R33949 vdd.n31137 vdd.n31136 25.6
R33950 vdd.n31138 vdd.n31137 25.6
R33951 vdd.n31139 vdd.n31138 25.6
R33952 vdd.n31140 vdd.n31139 25.6
R33953 vdd.n35705 vdd.n35704 25.6
R33954 vdd.n35704 vdd.n35703 25.6
R33955 vdd.n35703 vdd.n35702 25.6
R33956 vdd.n35702 vdd.n35701 25.6
R33957 vdd.n35701 vdd.n35700 25.6
R33958 vdd.n2730 vdd.n2729 25.6
R33959 vdd.n2731 vdd.n2730 25.6
R33960 vdd.n2732 vdd.n2731 25.6
R33961 vdd.n2733 vdd.n2732 25.6
R33962 vdd.n2734 vdd.n2733 25.6
R33963 vdd.n14527 vdd.n14526 25.6
R33964 vdd.n14526 vdd.n14525 25.6
R33965 vdd.n14525 vdd.n14523 25.6
R33966 vdd.n14523 vdd.n14521 25.6
R33967 vdd.n14521 vdd.n14519 25.6
R33968 vdd.n14519 vdd.n14517 25.6
R33969 vdd.n14517 vdd.n14515 25.6
R33970 vdd.n14515 vdd.n14513 25.6
R33971 vdd.n14513 vdd.n14511 25.6
R33972 vdd.n14511 vdd.n14509 25.6
R33973 vdd.n14509 vdd.n14507 25.6
R33974 vdd.n14507 vdd.n14505 25.6
R33975 vdd.n14505 vdd.n14503 25.6
R33976 vdd.n13115 vdd.n9210 25.6
R33977 vdd.n13200 vdd.n9210 25.6
R33978 vdd.n13201 vdd.n13200 25.6
R33979 vdd.n13202 vdd.n13201 25.6
R33980 vdd.n13202 vdd.n9168 25.6
R33981 vdd.n13259 vdd.n9168 25.6
R33982 vdd.n13260 vdd.n13259 25.6
R33983 vdd.n13263 vdd.n13260 25.6
R33984 vdd.n13263 vdd.n13262 25.6
R33985 vdd.n13262 vdd.n13261 25.6
R33986 vdd.n13261 vdd.n9091 25.6
R33987 vdd.n13350 vdd.n9091 25.6
R33988 vdd.n13351 vdd.n13350 25.6
R33989 vdd.n13352 vdd.n13351 25.6
R33990 vdd.n13352 vdd.n9043 25.6
R33991 vdd.n13406 vdd.n9043 25.6
R33992 vdd.n13407 vdd.n13406 25.6
R33993 vdd.n13408 vdd.n13407 25.6
R33994 vdd.n13408 vdd.n8990 25.6
R33995 vdd.n13494 vdd.n8990 25.6
R33996 vdd.n13495 vdd.n13494 25.6
R33997 vdd.n13496 vdd.n13495 25.6
R33998 vdd.n13496 vdd.n8947 25.6
R33999 vdd.n13550 vdd.n8947 25.6
R34000 vdd.n13551 vdd.n13550 25.6
R34001 vdd.n13554 vdd.n13551 25.6
R34002 vdd.n13554 vdd.n13553 25.6
R34003 vdd.n13553 vdd.n13552 25.6
R34004 vdd.n13552 vdd.n8871 25.6
R34005 vdd.n13642 vdd.n8871 25.6
R34006 vdd.n13643 vdd.n13642 25.6
R34007 vdd.n13644 vdd.n13643 25.6
R34008 vdd.n13644 vdd.n8822 25.6
R34009 vdd.n13699 vdd.n8822 25.6
R34010 vdd.n13700 vdd.n13699 25.6
R34011 vdd.n13701 vdd.n13700 25.6
R34012 vdd.n13701 vdd.n8774 25.6
R34013 vdd.n13774 vdd.n8774 25.6
R34014 vdd.n13775 vdd.n13774 25.6
R34015 vdd.n13776 vdd.n13775 25.6
R34016 vdd.n13776 vdd.n8729 25.6
R34017 vdd.n13835 vdd.n8729 25.6
R34018 vdd.n13836 vdd.n13835 25.6
R34019 vdd.n13837 vdd.n13836 25.6
R34020 vdd.n13837 vdd.n8679 25.6
R34021 vdd.n13901 vdd.n8679 25.6
R34022 vdd.n13902 vdd.n13901 25.6
R34023 vdd.n13903 vdd.n13902 25.6
R34024 vdd.n13903 vdd.n8617 25.6
R34025 vdd.n13969 vdd.n8617 25.6
R34026 vdd.n13970 vdd.n13969 25.6
R34027 vdd.n13972 vdd.n13970 25.6
R34028 vdd.n13972 vdd.n13971 25.6
R34029 vdd.n13971 vdd.n8562 25.6
R34030 vdd.n14064 vdd.n8562 25.6
R34031 vdd.n14065 vdd.n14064 25.6
R34032 vdd.n14066 vdd.n14065 25.6
R34033 vdd.n14066 vdd.n8510 25.6
R34034 vdd.n14120 vdd.n8510 25.6
R34035 vdd.n14121 vdd.n14120 25.6
R34036 vdd.n14123 vdd.n14121 25.6
R34037 vdd.n14123 vdd.n14122 25.6
R34038 vdd.n14122 vdd.n8455 25.6
R34039 vdd.n14190 vdd.n8455 25.6
R34040 vdd.n14191 vdd.n14190 25.6
R34041 vdd.n14192 vdd.n14191 25.6
R34042 vdd.n14192 vdd.n8395 25.6
R34043 vdd.n14259 vdd.n8395 25.6
R34044 vdd.n14260 vdd.n14259 25.6
R34045 vdd.n14262 vdd.n14260 25.6
R34046 vdd.n14262 vdd.n14261 25.6
R34047 vdd.n14261 vdd.n8344 25.6
R34048 vdd.n14339 vdd.n8344 25.6
R34049 vdd.n14340 vdd.n14339 25.6
R34050 vdd.n14343 vdd.n14340 25.6
R34051 vdd.n14343 vdd.n14342 25.6
R34052 vdd.n14342 vdd.n14341 25.6
R34053 vdd.n14341 vdd.n8271 25.6
R34054 vdd.n14432 vdd.n8271 25.6
R34055 vdd.n14433 vdd.n14432 25.6
R34056 vdd.n14435 vdd.n14433 25.6
R34057 vdd.n14435 vdd.n14434 25.6
R34058 vdd.n14434 vdd.n8213 25.6
R34059 vdd.n14502 vdd.n8213 25.6
R34060 vdd.n13107 vdd.n13106 25.6
R34061 vdd.n13106 vdd.n13105 25.6
R34062 vdd.n13105 vdd.n13103 25.6
R34063 vdd.n13103 vdd.n13100 25.6
R34064 vdd.n13100 vdd.n13099 25.6
R34065 vdd.n13099 vdd.n13096 25.6
R34066 vdd.n13096 vdd.n13095 25.6
R34067 vdd.n13095 vdd.n13092 25.6
R34068 vdd.n13092 vdd.n13091 25.6
R34069 vdd.n13091 vdd.n13088 25.6
R34070 vdd.n13088 vdd.n9274 25.6
R34071 vdd.n13113 vdd.n9274 25.6
R34072 vdd.n13114 vdd.n13113 25.6
R34073 vdd.n14599 vdd.n14598 25.6
R34074 vdd.n14598 vdd.n14597 25.6
R34075 vdd.n14597 vdd.n14595 25.6
R34076 vdd.n14595 vdd.n14592 25.6
R34077 vdd.n14592 vdd.n14591 25.6
R34078 vdd.n14591 vdd.n14588 25.6
R34079 vdd.n14588 vdd.n14587 25.6
R34080 vdd.n14587 vdd.n14584 25.6
R34081 vdd.n14584 vdd.n14583 25.6
R34082 vdd.n14583 vdd.n14580 25.6
R34083 vdd.n14580 vdd.n14579 25.6
R34084 vdd.n14579 vdd.n14576 25.6
R34085 vdd.n14576 vdd.n8143 25.6
R34086 vdd.n14972 vdd.n7984 25.6
R34087 vdd.n14966 vdd.n7984 25.6
R34088 vdd.n14966 vdd.n14965 25.6
R34089 vdd.n14965 vdd.n14963 25.6
R34090 vdd.n14963 vdd.n14961 25.6
R34091 vdd.n14961 vdd.n14959 25.6
R34092 vdd.n14959 vdd.n14957 25.6
R34093 vdd.n14957 vdd.n14955 25.6
R34094 vdd.n14955 vdd.n14953 25.6
R34095 vdd.n14953 vdd.n14951 25.6
R34096 vdd.n14951 vdd.n14949 25.6
R34097 vdd.n14949 vdd.n14947 25.6
R34098 vdd.n14947 vdd.n14945 25.6
R34099 vdd.n14659 vdd.n14658 25.6
R34100 vdd.n14660 vdd.n14659 25.6
R34101 vdd.n14660 vdd.n8122 25.6
R34102 vdd.n14697 vdd.n8122 25.6
R34103 vdd.n14698 vdd.n14697 25.6
R34104 vdd.n14700 vdd.n14698 25.6
R34105 vdd.n14700 vdd.n14699 25.6
R34106 vdd.n14699 vdd.n8102 25.6
R34107 vdd.n14743 vdd.n8102 25.6
R34108 vdd.n14744 vdd.n14743 25.6
R34109 vdd.n14746 vdd.n14744 25.6
R34110 vdd.n14746 vdd.n14745 25.6
R34111 vdd.n14745 vdd.n8080 25.6
R34112 vdd.n14776 vdd.n8080 25.6
R34113 vdd.n14777 vdd.n14776 25.6
R34114 vdd.n14778 vdd.n14777 25.6
R34115 vdd.n14778 vdd.n8052 25.6
R34116 vdd.n14830 vdd.n8052 25.6
R34117 vdd.n14831 vdd.n14830 25.6
R34118 vdd.n14832 vdd.n14831 25.6
R34119 vdd.n14832 vdd.n8032 25.6
R34120 vdd.n14871 vdd.n8032 25.6
R34121 vdd.n14872 vdd.n14871 25.6
R34122 vdd.n14873 vdd.n14872 25.6
R34123 vdd.n14873 vdd.n8018 25.6
R34124 vdd.n14908 vdd.n8018 25.6
R34125 vdd.n14909 vdd.n14908 25.6
R34126 vdd.n14911 vdd.n14909 25.6
R34127 vdd.n14911 vdd.n14910 25.6
R34128 vdd.n14910 vdd.n7999 25.6
R34129 vdd.n14944 vdd.n7999 25.6
R34130 vdd.n14641 vdd.n14640 25.6
R34131 vdd.n14640 vdd.n14639 25.6
R34132 vdd.n14639 vdd.n14637 25.6
R34133 vdd.n14637 vdd.n14634 25.6
R34134 vdd.n14634 vdd.n14633 25.6
R34135 vdd.n14633 vdd.n14630 25.6
R34136 vdd.n14630 vdd.n14629 25.6
R34137 vdd.n14629 vdd.n14626 25.6
R34138 vdd.n14626 vdd.n14625 25.6
R34139 vdd.n14625 vdd.n14622 25.6
R34140 vdd.n14622 vdd.n14621 25.6
R34141 vdd.n14621 vdd.n14618 25.6
R34142 vdd.n14618 vdd.n14617 25.6
R34143 vdd.n11577 vdd.n9242 25.6
R34144 vdd.n13147 vdd.n9242 25.6
R34145 vdd.n13148 vdd.n13147 25.6
R34146 vdd.n13150 vdd.n13148 25.6
R34147 vdd.n13150 vdd.n13149 25.6
R34148 vdd.n13149 vdd.n9188 25.6
R34149 vdd.n13231 vdd.n9188 25.6
R34150 vdd.n13232 vdd.n13231 25.6
R34151 vdd.n13235 vdd.n13232 25.6
R34152 vdd.n13235 vdd.n13234 25.6
R34153 vdd.n13234 vdd.n13233 25.6
R34154 vdd.n13233 vdd.n9128 25.6
R34155 vdd.n13318 vdd.n9128 25.6
R34156 vdd.n13319 vdd.n13318 25.6
R34157 vdd.n13325 vdd.n13319 25.6
R34158 vdd.n13325 vdd.n13324 25.6
R34159 vdd.n13324 vdd.n13323 25.6
R34160 vdd.n13323 vdd.n13320 25.6
R34161 vdd.n13320 vdd.n9018 25.6
R34162 vdd.n13440 vdd.n9018 25.6
R34163 vdd.n13441 vdd.n13440 25.6
R34164 vdd.n13443 vdd.n13441 25.6
R34165 vdd.n13443 vdd.n13442 25.6
R34166 vdd.n13442 vdd.n8967 25.6
R34167 vdd.n13523 vdd.n8967 25.6
R34168 vdd.n13524 vdd.n13523 25.6
R34169 vdd.n13527 vdd.n13524 25.6
R34170 vdd.n13527 vdd.n13526 25.6
R34171 vdd.n13526 vdd.n13525 25.6
R34172 vdd.n13525 vdd.n8907 25.6
R34173 vdd.n13610 vdd.n8907 25.6
R34174 vdd.n13611 vdd.n13610 25.6
R34175 vdd.n13617 vdd.n13611 25.6
R34176 vdd.n13617 vdd.n13616 25.6
R34177 vdd.n13616 vdd.n13615 25.6
R34178 vdd.n13615 vdd.n13612 25.6
R34179 vdd.n13612 vdd.n8798 25.6
R34180 vdd.n13732 vdd.n8798 25.6
R34181 vdd.n13733 vdd.n13732 25.6
R34182 vdd.n13734 vdd.n13733 25.6
R34183 vdd.n13734 vdd.n8751 25.6
R34184 vdd.n13805 vdd.n8751 25.6
R34185 vdd.n13806 vdd.n13805 25.6
R34186 vdd.n13807 vdd.n13806 25.6
R34187 vdd.n13807 vdd.n8710 25.6
R34188 vdd.n13866 vdd.n8710 25.6
R34189 vdd.n13867 vdd.n13866 25.6
R34190 vdd.n13868 vdd.n13867 25.6
R34191 vdd.n13868 vdd.n8644 25.6
R34192 vdd.n13929 vdd.n8644 25.6
R34193 vdd.n13930 vdd.n13929 25.6
R34194 vdd.n13932 vdd.n13930 25.6
R34195 vdd.n13932 vdd.n13931 25.6
R34196 vdd.n13931 vdd.n8591 25.6
R34197 vdd.n14006 vdd.n8591 25.6
R34198 vdd.n14007 vdd.n14006 25.6
R34199 vdd.n14009 vdd.n14007 25.6
R34200 vdd.n14009 vdd.n14008 25.6
R34201 vdd.n14008 vdd.n8538 25.6
R34202 vdd.n14092 vdd.n8538 25.6
R34203 vdd.n14093 vdd.n14092 25.6
R34204 vdd.n14094 vdd.n14093 25.6
R34205 vdd.n14094 vdd.n8487 25.6
R34206 vdd.n14155 vdd.n8487 25.6
R34207 vdd.n14156 vdd.n14155 25.6
R34208 vdd.n14157 vdd.n14156 25.6
R34209 vdd.n14157 vdd.n8423 25.6
R34210 vdd.n14219 vdd.n8423 25.6
R34211 vdd.n14220 vdd.n14219 25.6
R34212 vdd.n14222 vdd.n14220 25.6
R34213 vdd.n14222 vdd.n14221 25.6
R34214 vdd.n14221 vdd.n8369 25.6
R34215 vdd.n14297 vdd.n8369 25.6
R34216 vdd.n14298 vdd.n14297 25.6
R34217 vdd.n14299 vdd.n14298 25.6
R34218 vdd.n14299 vdd.n8315 25.6
R34219 vdd.n14374 vdd.n8315 25.6
R34220 vdd.n14375 vdd.n14374 25.6
R34221 vdd.n14379 vdd.n14375 25.6
R34222 vdd.n14379 vdd.n14378 25.6
R34223 vdd.n14378 vdd.n14377 25.6
R34224 vdd.n14377 vdd.n8237 25.6
R34225 vdd.n14463 vdd.n8237 25.6
R34226 vdd.n14464 vdd.n14463 25.6
R34227 vdd.n14466 vdd.n14464 25.6
R34228 vdd.n14466 vdd.n14465 25.6
R34229 vdd.n14465 vdd.n8185 25.6
R34230 vdd.n14561 vdd.n8185 25.6
R34231 vdd.n14562 vdd.n14561 25.6
R34232 vdd.n14564 vdd.n14562 25.6
R34233 vdd.n14564 vdd.n14563 25.6
R34234 vdd.n14563 vdd.n8170 25.6
R34235 vdd.n11655 vdd.n11654 25.6
R34236 vdd.n11654 vdd.n11653 25.6
R34237 vdd.n11653 vdd.n11651 25.6
R34238 vdd.n11651 vdd.n11648 25.6
R34239 vdd.n11648 vdd.n11647 25.6
R34240 vdd.n11647 vdd.n11644 25.6
R34241 vdd.n11644 vdd.n11643 25.6
R34242 vdd.n11643 vdd.n11640 25.6
R34243 vdd.n11640 vdd.n11639 25.6
R34244 vdd.n11639 vdd.n11636 25.6
R34245 vdd.n11636 vdd.n11635 25.6
R34246 vdd.n11635 vdd.n11632 25.6
R34247 vdd.n11632 vdd.n11631 25.6
R34248 vdd.n19967 vdd.n19965 25.6
R34249 vdd.n19965 vdd.n19963 25.6
R34250 vdd.n19963 vdd.n19961 25.6
R34251 vdd.n19961 vdd.n19960 25.6
R34252 vdd.n19960 vdd.n19959 25.6
R34253 vdd.n19959 vdd.n19958 25.6
R34254 vdd.n19958 vdd.n19957 25.6
R34255 vdd.n19957 vdd.n19956 25.6
R34256 vdd.n19956 vdd.n19955 25.6
R34257 vdd.n20516 vdd.n20515 25.6
R34258 vdd.n19297 vdd.n19295 25.6
R34259 vdd.n19295 vdd.n19294 25.6
R34260 vdd.n19294 vdd.n19293 25.6
R34261 vdd.n19293 vdd.n19292 25.6
R34262 vdd.n19292 vdd.n19291 25.6
R34263 vdd.n19291 vdd.n19290 25.6
R34264 vdd.n19290 vdd.n19289 25.6
R34265 vdd.n18460 vdd.n18458 25.6
R34266 vdd.n18458 vdd.n18457 25.6
R34267 vdd.n18457 vdd.n18456 25.6
R34268 vdd.n18456 vdd.n18455 25.6
R34269 vdd.n18455 vdd.n18454 25.6
R34270 vdd.n18454 vdd.n18453 25.6
R34271 vdd.n18453 vdd.n18452 25.6
R34272 vdd.n21666 vdd.n21665 25.6
R34273 vdd.n21613 vdd.n21612 25.6
R34274 vdd.n19149 vdd.n19148 25.6
R34275 vdd.n21007 vdd.n21006 25.6
R34276 vdd.n21006 vdd.n21005 25.6
R34277 vdd.n21642 vdd.n21641 25.6
R34278 vdd.n21641 vdd.n21640 25.6
R34279 vdd.n21640 vdd.n21639 25.6
R34280 vdd.n21639 vdd.n21638 25.6
R34281 vdd.n21638 vdd.n21637 25.6
R34282 vdd.n20024 vdd.n20022 25.6
R34283 vdd.n20022 vdd.n20021 25.6
R34284 vdd.n20021 vdd.n20020 25.6
R34285 vdd.n20020 vdd.n20019 25.6
R34286 vdd.n20019 vdd.n20018 25.6
R34287 vdd.n20018 vdd.n20017 25.6
R34288 vdd.n20017 vdd.n20016 25.6
R34289 vdd.n20477 vdd.n20476 25.6
R34290 vdd.n20476 vdd.n20475 25.6
R34291 vdd.n24671 vdd.n24670 25.6
R34292 vdd.n24670 vdd.n24668 25.6
R34293 vdd.n24668 vdd.n24666 25.6
R34294 vdd.n24666 vdd.n24664 25.6
R34295 vdd.n24664 vdd.n24662 25.6
R34296 vdd.n24662 vdd.n24660 25.6
R34297 vdd.n24660 vdd.n24658 25.6
R34298 vdd.n24658 vdd.n24656 25.6
R34299 vdd.n24656 vdd.n24654 25.6
R34300 vdd.n24654 vdd.n24652 25.6
R34301 vdd.n24652 vdd.n24650 25.6
R34302 vdd.n24650 vdd.n24648 25.6
R34303 vdd.n24648 vdd.n24646 25.6
R34304 vdd.n24644 vdd.n24643 25.6
R34305 vdd.n24643 vdd.n24642 25.6
R34306 vdd.n24642 vdd.n24641 25.6
R34307 vdd.n24641 vdd.n24640 25.6
R34308 vdd.n24640 vdd.n24639 25.6
R34309 vdd.n24639 vdd.n24638 25.6
R34310 vdd.n24638 vdd.n24637 25.6
R34311 vdd.n25056 vdd.n25055 25.6
R34312 vdd.n25057 vdd.n25056 25.6
R34313 vdd.n25058 vdd.n25057 25.6
R34314 vdd.n25059 vdd.n25058 25.6
R34315 vdd.n25060 vdd.n25059 25.6
R34316 vdd.n25061 vdd.n25060 25.6
R34317 vdd.n25089 vdd.n25087 25.6
R34318 vdd.n25087 vdd.n25085 25.6
R34319 vdd.n25085 vdd.n25083 25.6
R34320 vdd.n25083 vdd.n25081 25.6
R34321 vdd.n25081 vdd.n25079 25.6
R34322 vdd.n25079 vdd.n25077 25.6
R34323 vdd.n25077 vdd.n25075 25.6
R34324 vdd.n25075 vdd.n25073 25.6
R34325 vdd.n25073 vdd.n25071 25.6
R34326 vdd.n25071 vdd.n25069 25.6
R34327 vdd.n25069 vdd.n25067 25.6
R34328 vdd.n25067 vdd.n25065 25.6
R34329 vdd.n25065 vdd.n25063 25.6
R34330 vdd.n36013 vdd.n36012 25.551
R34331 vdd.n36055 vdd.n36054 25.551
R34332 vdd.n36244 vdd.n36243 25.551
R34333 vdd.n36286 vdd.n36285 25.551
R34334 vdd.n36475 vdd.n36474 25.551
R34335 vdd.n36517 vdd.n36516 25.551
R34336 vdd.n36706 vdd.n36705 25.551
R34337 vdd.n36748 vdd.n36747 25.551
R34338 vdd.n36937 vdd.n36936 25.551
R34339 vdd.n35684 vdd.n35683 25.551
R34340 vdd.n37145 vdd.n37144 25.551
R34341 vdd.n37173 vdd.n37172 25.551
R34342 vdd.n32986 vdd.n32985 25.551
R34343 vdd.n32972 vdd.n32971 25.551
R34344 vdd.n37520 vdd.n37519 25.551
R34345 vdd.n37566 vdd.n37565 25.551
R34346 vdd.n38034 vdd.n38033 25.551
R34347 vdd.n37992 vdd.n37991 25.551
R34348 vdd.n37803 vdd.n37802 25.551
R34349 vdd.n37761 vdd.n37760 25.551
R34350 vdd.n28203 vdd.n28202 25.551
R34351 vdd.n28245 vdd.n28244 25.551
R34352 vdd.n28434 vdd.n28433 25.551
R34353 vdd.n28476 vdd.n28475 25.551
R34354 vdd.n28665 vdd.n28664 25.551
R34355 vdd.n28707 vdd.n28706 25.551
R34356 vdd.n28110 vdd.n28109 25.551
R34357 vdd.n28084 vdd.n28083 25.551
R34358 vdd.n31627 vdd.n31626 25.551
R34359 vdd.n32065 vdd.n32064 25.551
R34360 vdd.n29718 vdd.n29717 25.551
R34361 vdd.n30186 vdd.n30185 25.551
R34362 vdd.n2874 vdd.n2873 25.551
R34363 vdd.n2906 vdd.n2905 25.551
R34364 vdd.n3055 vdd.n3054 25.551
R34365 vdd.n3087 vdd.n3086 25.551
R34366 vdd.n3236 vdd.n3235 25.551
R34367 vdd.n3268 vdd.n3267 25.551
R34368 vdd.n3417 vdd.n3416 25.551
R34369 vdd.n3449 vdd.n3448 25.551
R34370 vdd.n3598 vdd.n3597 25.551
R34371 vdd.n3640 vdd.n3639 25.551
R34372 vdd.n3918 vdd.n3917 25.551
R34373 vdd.n3852 vdd.n3851 25.551
R34374 vdd.n2418 vdd.n2417 25.551
R34375 vdd.n2477 vdd.n2476 25.551
R34376 vdd.n1863 vdd.n1862 25.551
R34377 vdd.n1796 vdd.n1795 25.551
R34378 vdd.n1668 vdd.n1667 25.551
R34379 vdd.n1636 vdd.n1635 25.551
R34380 vdd.n1487 vdd.n1486 25.551
R34381 vdd.n1455 vdd.n1454 25.551
R34382 vdd.n1306 vdd.n1305 25.551
R34383 vdd.n26772 vdd.n26771 25.551
R34384 vdd.n26921 vdd.n26920 25.551
R34385 vdd.n26953 vdd.n26952 25.551
R34386 vdd.n27102 vdd.n27101 25.551
R34387 vdd.n27134 vdd.n27133 25.551
R34388 vdd.n26617 vdd.n26616 25.551
R34389 vdd.n26345 vdd.n26344 25.551
R34390 vdd.n31623 vdd.n31622 25.551
R34391 vdd.n32061 vdd.n32060 25.551
R34392 vdd.n31473 vdd.n31472 25.551
R34393 vdd.n32504 vdd.n32503 25.551
R34394 vdd.n13367 vdd.n9068 25.551
R34395 vdd.n9054 vdd.n9053 25.551
R34396 vdd.n13659 vdd.n8848 25.551
R34397 vdd.n8834 vdd.n8833 25.551
R34398 vdd.n8665 vdd.n8659 25.551
R34399 vdd.n13979 vdd.n13978 25.551
R34400 vdd.n8442 vdd.n8439 25.551
R34401 vdd.n14269 vdd.n14268 25.551
R34402 vdd.n14694 vdd.n8127 25.551
R34403 vdd.n14740 vdd.n8106 25.551
R34404 vdd.n14868 vdd.n8037 25.551
R34405 vdd.n14897 vdd.n14885 25.551
R34406 vdd.n9202 vdd.n9184 25.551
R34407 vdd.n13285 vdd.n9139 25.551
R34408 vdd.n8980 vdd.n8963 25.551
R34409 vdd.n13577 vdd.n8917 25.551
R34410 vdd.n8748 vdd.n8747 25.551
R34411 vdd.n13872 vdd.n8702 25.551
R34412 vdd.n8534 vdd.n8526 25.551
R34413 vdd.n14161 vdd.n8479 25.551
R34414 vdd.n8306 vdd.n8295 25.551
R34415 vdd.n14441 vdd.n8263 25.551
R34416 vdd.n19274 vdd.n19273 25.551
R34417 vdd.n19238 vdd.n19237 25.551
R34418 vdd.n19218 vdd.n19217 25.551
R34419 vdd.n19181 vdd.n19180 25.551
R34420 vdd.n19835 vdd.n19834 25.551
R34421 vdd.n19872 vdd.n19871 25.551
R34422 vdd.n19904 vdd.n19903 25.551
R34423 vdd.n19940 vdd.n19939 25.551
R34424 vdd.n21539 vdd.n21538 25.551
R34425 vdd.n21489 vdd.n21488 25.551
R34426 vdd.n21280 vdd.n21279 25.551
R34427 vdd.n21230 vdd.n21229 25.551
R34428 vdd.n21023 vdd.n21022 25.551
R34429 vdd.n19123 vdd.n19122 25.551
R34430 vdd.n18914 vdd.n18913 25.551
R34431 vdd.n18864 vdd.n18863 25.551
R34432 vdd.n18655 vdd.n18654 25.551
R34433 vdd.n18605 vdd.n18604 25.551
R34434 vdd.n20421 vdd.n20415 25.551
R34435 vdd.n20363 vdd.n20357 25.551
R34436 vdd.n20185 vdd.n20179 25.551
R34437 vdd.n20127 vdd.n20121 25.551
R34438 vdd.n24728 vdd.n24727 25.551
R34439 vdd.n25186 vdd.n25185 25.551
R34440 vdd.n24499 vdd.t200 24.861
R34441 vdd.n24158 vdd.n24154 24.705
R34442 vdd.n24020 vdd.n24016 24.705
R34443 vdd.n23926 vdd.n23922 24.705
R34444 vdd.n23788 vdd.n23784 24.705
R34445 vdd.n23694 vdd.n23690 24.705
R34446 vdd.n23100 vdd.n23096 24.705
R34447 vdd.n23238 vdd.n23234 24.705
R34448 vdd.n23332 vdd.n23328 24.705
R34449 vdd.n23470 vdd.n23466 24.705
R34450 vdd.n23564 vdd.n23560 24.705
R34451 vdd.n22521 vdd.n22517 24.705
R34452 vdd.n22659 vdd.n22655 24.705
R34453 vdd.n22753 vdd.n22749 24.705
R34454 vdd.n22891 vdd.n22887 24.705
R34455 vdd.n22985 vdd.n22981 24.705
R34456 vdd.n22432 vdd.n22428 24.705
R34457 vdd.n22235 vdd.n22234 24.705
R34458 vdd.n22288 vdd.n22284 24.705
R34459 vdd.n22111 vdd.n22110 24.705
R34460 vdd.n24260 vdd.n24256 24.705
R34461 vdd.n24755 vdd.n24754 24.373
R34462 vdd.n25157 vdd.n25156 24.373
R34463 vdd.n35842 vdd.n35841 24.364
R34464 vdd.n30501 vdd.n30500 24.364
R34465 vdd.n35884 vdd.n35880 23.586
R34466 vdd.n35961 vdd.n35957 23.586
R34467 vdd.n36115 vdd.n36111 23.586
R34468 vdd.n36192 vdd.n36188 23.586
R34469 vdd.n36346 vdd.n36342 23.586
R34470 vdd.n36423 vdd.n36419 23.586
R34471 vdd.n36577 vdd.n36573 23.586
R34472 vdd.n36654 vdd.n36650 23.586
R34473 vdd.n36808 vdd.n36804 23.586
R34474 vdd.n36885 vdd.n36881 23.586
R34475 vdd.n33282 vdd.n33281 23.586
R34476 vdd.n33219 vdd.n33215 23.586
R34477 vdd.n37218 vdd.n37217 23.586
R34478 vdd.n37278 vdd.n37274 23.586
R34479 vdd.n37419 vdd.n37415 23.586
R34480 vdd.n37481 vdd.n37477 23.586
R34481 vdd.n38167 vdd.n38163 23.586
R34482 vdd.n38094 vdd.n38090 23.586
R34483 vdd.n37940 vdd.n37936 23.586
R34484 vdd.n37863 vdd.n37859 23.586
R34485 vdd.n37709 vdd.n37705 23.586
R34486 vdd.n37632 vdd.n37628 23.586
R34487 vdd.n28305 vdd.n28301 23.586
R34488 vdd.n28382 vdd.n28378 23.586
R34489 vdd.n28536 vdd.n28532 23.586
R34490 vdd.n28613 vdd.n28609 23.586
R34491 vdd.n28767 vdd.n28763 23.586
R34492 vdd.n28174 vdd.n28170 23.586
R34493 vdd.n28989 vdd.n28985 23.586
R34494 vdd.n27793 vdd.n27789 23.586
R34495 vdd.n31571 vdd.n31570 23.586
R34496 vdd.n29818 vdd.n29814 23.586
R34497 vdd.n30273 vdd.n30269 23.586
R34498 vdd.n30529 vdd.n30528 23.586
R34499 vdd.n2770 vdd.n2769 23.586
R34500 vdd.n2831 vdd.n2830 23.586
R34501 vdd.n2951 vdd.n2950 23.586
R34502 vdd.n3012 vdd.n3011 23.586
R34503 vdd.n3132 vdd.n3131 23.586
R34504 vdd.n3193 vdd.n3192 23.586
R34505 vdd.n3313 vdd.n3312 23.586
R34506 vdd.n3374 vdd.n3373 23.586
R34507 vdd.n3494 vdd.n3493 23.586
R34508 vdd.n3555 vdd.n3554 23.586
R34509 vdd.n2721 vdd.n2717 23.586
R34510 vdd.n3980 vdd.n3979 23.586
R34511 vdd.n2178 vdd.n2174 23.586
R34512 vdd.n2339 vdd.n2338 23.586
R34513 vdd.n2654 vdd.n2653 23.586
R34514 vdd.n1937 vdd.n1936 23.586
R34515 vdd.n1768 vdd.n1767 23.586
R34516 vdd.n1713 vdd.n1712 23.586
R34517 vdd.n1593 vdd.n1592 23.586
R34518 vdd.n1532 vdd.n1531 23.586
R34519 vdd.n1412 vdd.n1411 23.586
R34520 vdd.n1351 vdd.n1350 23.586
R34521 vdd.n26817 vdd.n26816 23.586
R34522 vdd.n26878 vdd.n26877 23.586
R34523 vdd.n26998 vdd.n26997 23.586
R34524 vdd.n27059 vdd.n27058 23.586
R34525 vdd.n27179 vdd.n27178 23.586
R34526 vdd.n26753 vdd.n26752 23.586
R34527 vdd.n31822 vdd.n31821 23.586
R34528 vdd.n31673 vdd.n31672 23.586
R34529 vdd.n31573 vdd.n31566 23.586
R34530 vdd.n31523 vdd.n31522 23.586
R34531 vdd.n31047 vdd.n31046 23.586
R34532 vdd.n31259 vdd.n31255 23.586
R34533 vdd.n13185 vdd.n9221 23.586
R34534 vdd.n13275 vdd.n9149 23.586
R34535 vdd.n13479 vdd.n9001 23.586
R34536 vdd.n13567 vdd.n8928 23.586
R34537 vdd.n13759 vdd.n8784 23.586
R34538 vdd.n13855 vdd.n8722 23.586
R34539 vdd.n14070 vdd.n8558 23.586
R34540 vdd.n14144 vdd.n8501 23.586
R34541 vdd.n14346 vdd.n8334 23.586
R34542 vdd.n14460 vdd.n8243 23.586
R34543 vdd.n14655 vdd.n8147 23.586
R34544 vdd.n14772 vdd.n8085 23.586
R34545 vdd.n14827 vdd.n8056 23.586
R34546 vdd.n14941 vdd.n7985 23.586
R34547 vdd.n13154 vdd.n9234 23.586
R34548 vdd.n13360 vdd.n9073 23.586
R34549 vdd.n13447 vdd.n9010 23.586
R34550 vdd.n13652 vdd.n8853 23.586
R34551 vdd.n13738 vdd.n8791 23.586
R34552 vdd.n8641 vdd.n8620 23.586
R34553 vdd.n14023 vdd.n14022 23.586
R34554 vdd.n8419 vdd.n8398 23.586
R34555 vdd.n14311 vdd.n8358 23.586
R34556 vdd.n14558 vdd.n8190 23.586
R34557 vdd.n19384 vdd.n19378 23.586
R34558 vdd.n19465 vdd.n19459 23.586
R34559 vdd.n19590 vdd.n19584 23.586
R34560 vdd.n19665 vdd.n19659 23.586
R34561 vdd.n19792 vdd.n19786 23.586
R34562 vdd.n20989 vdd.n20983 23.586
R34563 vdd.n19891 vdd.n19885 23.586
R34564 vdd.n20798 vdd.n20792 23.586
R34565 vdd.n20674 vdd.n20668 23.586
R34566 vdd.n20593 vdd.n20587 23.586
R34567 vdd.n21617 vdd.n21603 23.586
R34568 vdd.n21431 vdd.n21425 23.586
R34569 vdd.n21350 vdd.n21344 23.586
R34570 vdd.n21172 vdd.n21166 23.586
R34571 vdd.n21087 vdd.n21081 23.586
R34572 vdd.n19065 vdd.n19059 23.586
R34573 vdd.n18984 vdd.n18978 23.586
R34574 vdd.n18806 vdd.n18800 23.586
R34575 vdd.n18725 vdd.n18719 23.586
R34576 vdd.n18547 vdd.n18541 23.586
R34577 vdd.n19980 vdd.n19979 23.586
R34578 vdd.n20293 vdd.n20292 23.586
R34579 vdd.n20243 vdd.n20242 23.586
R34580 vdd.n20030 vdd.n20029 23.586
R34581 vdd.n24814 vdd.n24813 23.586
R34582 vdd.n25095 vdd.n25094 23.586
R34583 vdd.n21349 vdd.t345 23.222
R34584 vdd.t351 vdd.n21138 23.222
R34585 vdd.n18805 vdd.t277 23.222
R34586 vdd.n24114 vdd.n24113 22.619
R34587 vdd.n24060 vdd.n24059 22.619
R34588 vdd.n23882 vdd.n23881 22.619
R34589 vdd.n23828 vdd.n23827 22.619
R34590 vdd.n23650 vdd.n23649 22.619
R34591 vdd.n23140 vdd.n23139 22.619
R34592 vdd.n23194 vdd.n23193 22.619
R34593 vdd.n23372 vdd.n23371 22.619
R34594 vdd.n23426 vdd.n23425 22.619
R34595 vdd.n23604 vdd.n23603 22.619
R34596 vdd.n22561 vdd.n22560 22.619
R34597 vdd.n22615 vdd.n22614 22.619
R34598 vdd.n22793 vdd.n22792 22.619
R34599 vdd.n22847 vdd.n22846 22.619
R34600 vdd.n23025 vdd.n23024 22.619
R34601 vdd.n22388 vdd.n22387 22.619
R34602 vdd.n22358 vdd.n22357 22.619
R34603 vdd.n24333 vdd.n24332 22.619
R34604 vdd.n22087 vdd.n22086 22.619
R34605 vdd.n24216 vdd.n24215 22.619
R34606 vdd.n12560 vdd.n10500 21.824
R34607 vdd.n12560 vdd.n12559 21.824
R34608 vdd.n12559 vdd.n12558 21.824
R34609 vdd.n12558 vdd.n10501 21.824
R34610 vdd.n12552 vdd.n10501 21.824
R34611 vdd.n12552 vdd.n12551 21.824
R34612 vdd.n12551 vdd.n12550 21.824
R34613 vdd.n12550 vdd.n10505 21.824
R34614 vdd.n12544 vdd.n10505 21.824
R34615 vdd.n12544 vdd.n12543 21.824
R34616 vdd.n12536 vdd.n10512 21.824
R34617 vdd.n12535 vdd.n12534 21.824
R34618 vdd.n12534 vdd.n10513 21.824
R34619 vdd.n12528 vdd.n10513 21.824
R34620 vdd.n11926 vdd.n11925 21.824
R34621 vdd.n15103 vdd.n15101 21.824
R34622 vdd.n15101 vdd.n15099 21.824
R34623 vdd.n15099 vdd.n15097 21.824
R34624 vdd.n15097 vdd.n15095 21.824
R34625 vdd.n15095 vdd.n15093 21.824
R34626 vdd.n15093 vdd.n15091 21.824
R34627 vdd.n15091 vdd.n15089 21.824
R34628 vdd.n15089 vdd.n15087 21.824
R34629 vdd.n16841 vdd.n16839 21.824
R34630 vdd.n16847 vdd.n16845 21.824
R34631 vdd.n16851 vdd.n16849 21.824
R34632 vdd.n16853 vdd.n16851 21.824
R34633 vdd.n16864 vdd.n16853 21.824
R34634 vdd.n21707 vdd.n21706 21.824
R34635 vdd.n21000 vdd.n19152 21.814
R34636 vdd.n11914 vdd.n11913 21.772
R34637 vdd.n35710 vdd.n35709 21.62
R34638 vdd.n35999 vdd.n35998 21.62
R34639 vdd.n36069 vdd.n36068 21.62
R34640 vdd.n36230 vdd.n36229 21.62
R34641 vdd.n36300 vdd.n36299 21.62
R34642 vdd.n36461 vdd.n36460 21.62
R34643 vdd.n36531 vdd.n36530 21.62
R34644 vdd.n36692 vdd.n36691 21.62
R34645 vdd.n36762 vdd.n36761 21.62
R34646 vdd.n36923 vdd.n36922 21.62
R34647 vdd.n37004 vdd.n37003 21.62
R34648 vdd.n33170 vdd.n33169 21.62
R34649 vdd.n33132 vdd.n33131 21.62
R34650 vdd.n37311 vdd.n37310 21.62
R34651 vdd.n37383 vdd.n37382 21.62
R34652 vdd.n32844 vdd.n32843 21.62
R34653 vdd.n38208 vdd.n38207 21.62
R34654 vdd.n38048 vdd.n38047 21.62
R34655 vdd.n37978 vdd.n37977 21.62
R34656 vdd.n37817 vdd.n37816 21.62
R34657 vdd.n37747 vdd.n37746 21.62
R34658 vdd.n28189 vdd.n28188 21.62
R34659 vdd.n28259 vdd.n28258 21.62
R34660 vdd.n28420 vdd.n28419 21.62
R34661 vdd.n28490 vdd.n28489 21.62
R34662 vdd.n28651 vdd.n28650 21.62
R34663 vdd.n28721 vdd.n28720 21.62
R34664 vdd.n26208 vdd.n26207 21.62
R34665 vdd.n31753 vdd.n31752 21.62
R34666 vdd.n27834 vdd.n27833 21.62
R34667 vdd.n27910 vdd.n27909 21.62
R34668 vdd.n31486 vdd.n31485 21.62
R34669 vdd.n30217 vdd.n30216 21.62
R34670 vdd.n30346 vdd.n30345 21.62
R34671 vdd.n2739 vdd.n2738 21.62
R34672 vdd.n2863 vdd.n2862 21.62
R34673 vdd.n2917 vdd.n2916 21.62
R34674 vdd.n3044 vdd.n3043 21.62
R34675 vdd.n3098 vdd.n3097 21.62
R34676 vdd.n3225 vdd.n3224 21.62
R34677 vdd.n3279 vdd.n3278 21.62
R34678 vdd.n3406 vdd.n3405 21.62
R34679 vdd.n3460 vdd.n3459 21.62
R34680 vdd.n3587 vdd.n3586 21.62
R34681 vdd.n3650 vdd.n3649 21.62
R34682 vdd.n3935 vdd.n3934 21.62
R34683 vdd.n2216 vdd.n2215 21.62
R34684 vdd.n2399 vdd.n2398 21.62
R34685 vdd.n2599 vdd.n2598 21.62
R34686 vdd.n1223 vdd.n1222 21.62
R34687 vdd.n1780 vdd.n1779 21.62
R34688 vdd.n1679 vdd.n1678 21.62
R34689 vdd.n1625 vdd.n1624 21.62
R34690 vdd.n1498 vdd.n1497 21.62
R34691 vdd.n1444 vdd.n1443 21.62
R34692 vdd.n1317 vdd.n1316 21.62
R34693 vdd.n26783 vdd.n26782 21.62
R34694 vdd.n26910 vdd.n26909 21.62
R34695 vdd.n26964 vdd.n26963 21.62
R34696 vdd.n27091 vdd.n27090 21.62
R34697 vdd.n27145 vdd.n27144 21.62
R34698 vdd.n26204 vdd.n26203 21.62
R34699 vdd.n31749 vdd.n31748 21.62
R34700 vdd.n31640 vdd.n31639 21.62
R34701 vdd.n32096 vdd.n32095 21.62
R34702 vdd.n31482 vdd.n31481 21.62
R34703 vdd.n32483 vdd.n32482 21.62
R34704 vdd.n31145 vdd.n31144 21.62
R34705 vdd.n13119 vdd.n9272 21.62
R34706 vdd.n13347 vdd.n9096 21.62
R34707 vdd.n13411 vdd.n9041 21.62
R34708 vdd.n13639 vdd.n8876 21.62
R34709 vdd.n13705 vdd.n8820 21.62
R34710 vdd.n13906 vdd.n8658 21.62
R34711 vdd.n13991 vdd.n8603 21.62
R34712 vdd.n14196 vdd.n8437 21.62
R34713 vdd.n14282 vdd.n8381 21.62
R34714 vdd.n14499 vdd.n8211 21.62
R34715 vdd.n14675 vdd.n8133 21.62
R34716 vdd.n14732 vdd.n14723 21.62
R34717 vdd.n14847 vdd.n8043 21.62
R34718 vdd.n14886 vdd.n8015 21.62
R34719 vdd.n13228 vdd.n9193 21.62
R34720 vdd.n13315 vdd.n9133 21.62
R34721 vdd.n13520 vdd.n8971 21.62
R34722 vdd.n13607 vdd.n8911 21.62
R34723 vdd.n8764 vdd.n8745 21.62
R34724 vdd.n13880 vdd.n8696 21.62
R34725 vdd.n8551 vdd.n8533 21.62
R34726 vdd.n14169 vdd.n8473 21.62
R34727 vdd.n14382 vdd.n8305 21.62
R34728 vdd.n14469 vdd.n8231 21.62
R34729 vdd.n19303 vdd.n19302 21.62
R34730 vdd.n19506 vdd.n19505 21.62
R34731 vdd.n19536 vdd.n19535 21.62
R34732 vdd.n19707 vdd.n19706 21.62
R34733 vdd.n19738 vdd.n19737 21.62
R34734 vdd.n20935 vdd.n20934 21.62
R34735 vdd.n20904 vdd.n20903 21.62
R34736 vdd.n20745 vdd.n20744 21.62
R34737 vdd.n20715 vdd.n20714 21.62
R34738 vdd.n19973 vdd.n19972 21.62
R34739 vdd.n21555 vdd.n21554 21.62
R34740 vdd.n21473 vdd.n21472 21.62
R34741 vdd.n21296 vdd.n21295 21.62
R34742 vdd.n21214 vdd.n21213 21.62
R34743 vdd.n21037 vdd.n21036 21.62
R34744 vdd.n19107 vdd.n19106 21.62
R34745 vdd.n18930 vdd.n18929 21.62
R34746 vdd.n18848 vdd.n18847 21.62
R34747 vdd.n18671 vdd.n18670 21.62
R34748 vdd.n18589 vdd.n18588 21.62
R34749 vdd.n20437 vdd.n20431 21.62
R34750 vdd.n20347 vdd.n20341 21.62
R34751 vdd.n20201 vdd.n20195 21.62
R34752 vdd.n20111 vdd.n20105 21.62
R34753 vdd.n24715 vdd.n24714 21.62
R34754 vdd.n25198 vdd.n25197 21.62
R34755 vdd.n24767 vdd.n24766 21.501
R34756 vdd.n25145 vdd.n25144 21.501
R34757 vdd.n10264 vdd.n10263 21.379
R34758 vdd.n24126 vdd.n24125 21.176
R34759 vdd.n24044 vdd.n24043 21.176
R34760 vdd.n23894 vdd.n23893 21.176
R34761 vdd.n23812 vdd.n23811 21.176
R34762 vdd.n23662 vdd.n23661 21.176
R34763 vdd.n23124 vdd.n23123 21.176
R34764 vdd.n23206 vdd.n23205 21.176
R34765 vdd.n23356 vdd.n23355 21.176
R34766 vdd.n23438 vdd.n23437 21.176
R34767 vdd.n23588 vdd.n23587 21.176
R34768 vdd.n22545 vdd.n22544 21.176
R34769 vdd.n22627 vdd.n22626 21.176
R34770 vdd.n22777 vdd.n22776 21.176
R34771 vdd.n22859 vdd.n22858 21.176
R34772 vdd.n23009 vdd.n23008 21.176
R34773 vdd.n22398 vdd.n22397 21.176
R34774 vdd.n24343 vdd.n24342 21.176
R34775 vdd.n24226 vdd.n24225 21.176
R34776 vdd.n14781 vdd.n8073 21.059
R34777 vdd.n10599 vdd.n10596 20.617
R34778 vdd.n10758 vdd.n10750 20.617
R34779 vdd.n12284 vdd.n10916 20.617
R34780 vdd.n12180 vdd.n11094 20.617
R34781 vdd.n12075 vdd.n11269 20.617
R34782 vdd.n11978 vdd.n11425 20.617
R34783 vdd.n11601 vdd.n11600 20.617
R34784 vdd.n16977 vdd.n16972 20.617
R34785 vdd.n17249 vdd.n17244 20.617
R34786 vdd.n17521 vdd.n17516 20.617
R34787 vdd.n17779 vdd.n17774 20.617
R34788 vdd.n18050 vdd.n18045 20.617
R34789 vdd.n16816 vdd.n16812 20.617
R34790 vdd.n21703 vdd.n15017 20.617
R34791 vdd.n18530 vdd.t243 20.407
R34792 vdd.n13373 vdd.n9064 19.952
R34793 vdd.n13373 vdd.n9049 19.952
R34794 vdd.n13665 vdd.n8844 19.952
R34795 vdd.n13665 vdd.n8828 19.952
R34796 vdd.n13964 vdd.n13963 19.952
R34797 vdd.n13963 vdd.n8626 19.952
R34798 vdd.n14254 vdd.n14253 19.952
R34799 vdd.n14253 vdd.n8404 19.952
R34800 vdd.n13243 vdd.n13242 19.952
R34801 vdd.n13242 vdd.n9155 19.952
R34802 vdd.n13535 vdd.n13534 19.952
R34803 vdd.n13534 vdd.n8934 19.952
R34804 vdd.n13862 vdd.n8715 19.952
R34805 vdd.n13862 vdd.n8716 19.952
R34806 vdd.n14151 vdd.n8493 19.952
R34807 vdd.n14151 vdd.n8494 19.952
R34808 vdd.n14417 vdd.n8290 19.952
R34809 vdd.n14417 vdd.n8291 19.952
R34810 vdd.n21011 vdd.n19141 19.952
R34811 vdd.n21011 vdd.n19142 19.952
R34812 vdd.t359 vdd.n12542 19.898
R34813 vdd.n16843 vdd.t22 19.898
R34814 vdd.n35870 vdd.n35866 19.655
R34815 vdd.n35975 vdd.n35971 19.655
R34816 vdd.n36101 vdd.n36097 19.655
R34817 vdd.n36206 vdd.n36202 19.655
R34818 vdd.n36332 vdd.n36328 19.655
R34819 vdd.n36437 vdd.n36433 19.655
R34820 vdd.n36563 vdd.n36559 19.655
R34821 vdd.n36668 vdd.n36664 19.655
R34822 vdd.n36794 vdd.n36790 19.655
R34823 vdd.n36899 vdd.n36895 19.655
R34824 vdd.n37039 vdd.n37038 19.655
R34825 vdd.n37112 vdd.n37111 19.655
R34826 vdd.n33113 vdd.n33112 19.655
R34827 vdd.n33034 vdd.n33033 19.655
R34828 vdd.n37408 vdd.n37404 19.655
R34829 vdd.n32867 vdd.n32866 19.655
R34830 vdd.n38181 vdd.n38180 19.655
R34831 vdd.n38080 vdd.n38076 19.655
R34832 vdd.n37954 vdd.n37950 19.655
R34833 vdd.n37849 vdd.n37845 19.655
R34834 vdd.n37723 vdd.n37719 19.655
R34835 vdd.n37618 vdd.n37614 19.655
R34836 vdd.n28291 vdd.n28287 19.655
R34837 vdd.n28396 vdd.n28392 19.655
R34838 vdd.n28522 vdd.n28518 19.655
R34839 vdd.n28627 vdd.n28623 19.655
R34840 vdd.n28753 vdd.n28749 19.655
R34841 vdd.n28139 vdd.n28135 19.655
R34842 vdd.n28967 vdd.n28963 19.655
R34843 vdd.n27810 vdd.n27806 19.655
R34844 vdd.n29885 vdd.n29884 19.655
R34845 vdd.n31511 vdd.n31510 19.655
R34846 vdd.n32446 vdd.n32445 19.655
R34847 vdd.n30515 vdd.n30514 19.655
R34848 vdd.n2759 vdd.n2758 19.655
R34849 vdd.n2842 vdd.n2841 19.655
R34850 vdd.n2940 vdd.n2939 19.655
R34851 vdd.n3023 vdd.n3022 19.655
R34852 vdd.n3121 vdd.n3120 19.655
R34853 vdd.n3204 vdd.n3203 19.655
R34854 vdd.n3302 vdd.n3301 19.655
R34855 vdd.n3385 vdd.n3384 19.655
R34856 vdd.n3483 vdd.n3482 19.655
R34857 vdd.n3566 vdd.n3565 19.655
R34858 vdd.n2055 vdd.n2051 19.655
R34859 vdd.n2013 vdd.n2009 19.655
R34860 vdd.n2195 vdd.n2191 19.655
R34861 vdd.n2039 vdd.n2035 19.655
R34862 vdd.n2635 vdd.n2634 19.655
R34863 vdd.n1196 vdd.n1192 19.655
R34864 vdd.n1283 vdd.n1279 19.655
R34865 vdd.n1702 vdd.n1701 19.655
R34866 vdd.n1604 vdd.n1603 19.655
R34867 vdd.n1521 vdd.n1520 19.655
R34868 vdd.n1423 vdd.n1422 19.655
R34869 vdd.n1340 vdd.n1339 19.655
R34870 vdd.n26806 vdd.n26805 19.655
R34871 vdd.n26889 vdd.n26888 19.655
R34872 vdd.n26987 vdd.n26986 19.655
R34873 vdd.n27070 vdd.n27069 19.655
R34874 vdd.n27168 vdd.n27167 19.655
R34875 vdd.n27236 vdd.n27235 19.655
R34876 vdd.n31802 vdd.n31801 19.655
R34877 vdd.n31667 vdd.n31666 19.655
R34878 vdd.n32157 vdd.n32153 19.655
R34879 vdd.n31513 vdd.n31506 19.655
R34880 vdd.n32448 vdd.n32441 19.655
R34881 vdd.n31276 vdd.n31272 19.655
R34882 vdd.n13197 vdd.n9215 19.655
R34883 vdd.n13302 vdd.n9143 19.655
R34884 vdd.n13491 vdd.n8995 19.655
R34885 vdd.n13594 vdd.n8922 19.655
R34886 vdd.n13771 vdd.n8778 19.655
R34887 vdd.n13898 vdd.n8683 19.655
R34888 vdd.n14049 vdd.n8573 19.655
R34889 vdd.n14187 vdd.n8459 19.655
R34890 vdd.n14324 vdd.n8356 19.655
R34891 vdd.n14453 vdd.n8252 19.655
R34892 vdd.n14647 vdd.n8154 19.655
R34893 vdd.n14761 vdd.n8093 19.655
R34894 vdd.n14819 vdd.n14810 19.655
R34895 vdd.n14929 vdd.n8008 19.655
R34896 vdd.n13163 vdd.n13161 19.655
R34897 vdd.n9111 vdd.n9072 19.655
R34898 vdd.n13457 vdd.n13456 19.655
R34899 vdd.n8890 vdd.n8852 19.655
R34900 vdd.n13747 vdd.n8786 19.655
R34901 vdd.n8655 vdd.n8640 19.655
R34902 vdd.n14037 vdd.n8577 19.655
R34903 vdd.n8435 vdd.n8418 19.655
R34904 vdd.n14371 vdd.n8319 19.655
R34905 vdd.n14532 vdd.n8196 19.655
R34906 vdd.n19368 vdd.n19362 19.655
R34907 vdd.n19481 vdd.n19475 19.655
R34908 vdd.n19574 vdd.n19568 19.655
R34909 vdd.n19681 vdd.n19675 19.655
R34910 vdd.n19776 vdd.n19770 19.655
R34911 vdd.n20973 vdd.n20967 19.655
R34912 vdd.n20878 vdd.n20872 19.655
R34913 vdd.n20782 vdd.n20776 19.655
R34914 vdd.n20690 vdd.n20684 19.655
R34915 vdd.n20577 vdd.n20571 19.655
R34916 vdd.n21593 vdd.n21587 19.655
R34917 vdd.n21447 vdd.n21441 19.655
R34918 vdd.n21334 vdd.n21328 19.655
R34919 vdd.n21188 vdd.n21182 19.655
R34920 vdd.n21075 vdd.n21069 19.655
R34921 vdd.n19081 vdd.n19075 19.655
R34922 vdd.n18968 vdd.n18962 19.655
R34923 vdd.n18822 vdd.n18816 19.655
R34924 vdd.n18709 vdd.n18703 19.655
R34925 vdd.n18563 vdd.n18557 19.655
R34926 vdd.n20461 vdd.n20460 19.655
R34927 vdd.n20309 vdd.n20308 19.655
R34928 vdd.n20227 vdd.n20226 19.655
R34929 vdd.n20073 vdd.n20072 19.655
R34930 vdd.n24802 vdd.n24801 19.655
R34931 vdd.n25107 vdd.n25106 19.655
R34932 vdd.n11717 vdd.n11716 19.652
R34933 vdd.n11705 vdd.n11692 19.652
R34934 vdd.n11863 vdd.n11861 19.652
R34935 vdd.n11848 vdd.n11843 19.652
R34936 vdd.n21954 vdd.n21952 19.652
R34937 vdd.n21939 vdd.n21934 19.652
R34938 vdd.n12433 vdd.n10663 19.404
R34939 vdd.n10687 vdd.n10679 19.404
R34940 vdd.n10846 vdd.n10826 19.404
R34941 vdd.n10859 vdd.n10827 19.404
R34942 vdd.n11027 vdd.n11005 19.404
R34943 vdd.n12233 vdd.n11013 19.404
R34944 vdd.n12131 vdd.n11177 19.404
R34945 vdd.n12123 vdd.n11183 19.404
R34946 vdd.n11355 vdd.n11335 19.404
R34947 vdd.n11368 vdd.n11336 19.404
R34948 vdd.n10386 vdd.n10340 19.404
R34949 vdd.n10382 vdd.n10343 19.404
R34950 vdd.n9438 vdd.n9416 19.404
R34951 vdd.n12992 vdd.n9417 19.404
R34952 vdd.n12886 vdd.n9607 19.404
R34953 vdd.n12882 vdd.n9611 19.404
R34954 vdd.n9797 vdd.n9777 19.404
R34955 vdd.n12784 vdd.n9778 19.404
R34956 vdd.n12678 vdd.n9967 19.404
R34957 vdd.n12674 vdd.n9971 19.404
R34958 vdd.n10240 vdd.n10120 19.404
R34959 vdd.n12586 vdd.n10121 19.404
R34960 vdd.n17104 vdd.n17098 19.404
R34961 vdd.n17124 vdd.n17115 19.404
R34962 vdd.n17376 vdd.n17370 19.404
R34963 vdd.n17396 vdd.n17387 19.404
R34964 vdd.n17634 vdd.n17628 19.404
R34965 vdd.n17654 vdd.n17645 19.404
R34966 vdd.n17905 vdd.n17899 19.404
R34967 vdd.n17925 vdd.n17916 19.404
R34968 vdd.n18177 vdd.n18171 19.404
R34969 vdd.n18197 vdd.n18188 19.404
R34970 vdd.n15249 vdd.n15248 19.404
R34971 vdd.n15238 vdd.n15237 19.404
R34972 vdd.n15224 vdd.n15223 19.404
R34973 vdd.n15210 vdd.n15209 19.404
R34974 vdd.n15184 vdd.n15183 19.404
R34975 vdd.n15189 vdd.n15188 19.404
R34976 vdd.n15168 vdd.n15167 19.404
R34977 vdd.n15154 vdd.n15153 19.404
R34978 vdd.n15140 vdd.n15139 19.404
R34979 vdd.n15126 vdd.n15125 19.404
R34980 vdd.n16667 vdd.n16666 19.404
R34981 vdd.n16654 vdd.n16653 19.404
R34982 vdd.n19724 vdd.t142 19.351
R34983 vdd.n20921 vdd.t146 19.351
R34984 vdd.n12542 vdd.t362 19.256
R34985 vdd.n12536 vdd.t371 19.256
R34986 vdd.t6 vdd.n16843 19.256
R34987 vdd.t24 vdd.n16847 19.256
R34988 vdd.n14575 vdd.n8149 18.823
R34989 vdd.n14973 vdd.n7983 18.823
R34990 vdd.n25391 vdd.n25390 18.822
R34991 vdd.n11925 vdd.n11565 18.614
R34992 vdd.n21708 vdd.n21707 18.614
R34993 vdd.n24779 vdd.n24778 18.525
R34994 vdd.n25132 vdd.n25131 18.525
R34995 vdd.n13087 vdd.n9271 18.447
R34996 vdd.n14497 vdd.n8212 18.447
R34997 vdd.n10595 vdd.n10572 18.191
R34998 vdd.n12481 vdd.n10585 18.191
R34999 vdd.n12381 vdd.n10748 18.191
R35000 vdd.n10761 vdd.n10755 18.191
R35001 vdd.n10940 vdd.n10939 18.191
R35002 vdd.n12280 vdd.n10918 18.191
R35003 vdd.n11098 vdd.n11093 18.191
R35004 vdd.n11116 vdd.n11114 18.191
R35005 vdd.n12083 vdd.n11243 18.191
R35006 vdd.n12071 vdd.n11270 18.191
R35007 vdd.n11484 vdd.n11483 18.191
R35008 vdd.n11974 vdd.n11427 18.191
R35009 vdd.n10452 vdd.n10289 18.191
R35010 vdd.n10440 vdd.n10296 18.191
R35011 vdd.n9344 vdd.n9340 18.191
R35012 vdd.n13033 vdd.n9331 18.191
R35013 vdd.n12945 vdd.n9509 18.191
R35014 vdd.n9542 vdd.n9537 18.191
R35015 vdd.n9704 vdd.n9700 18.191
R35016 vdd.n12825 vdd.n9691 18.191
R35017 vdd.n12737 vdd.n9869 18.191
R35018 vdd.n9902 vdd.n9898 18.191
R35019 vdd.n10158 vdd.n10153 18.191
R35020 vdd.n12616 vdd.n10049 18.191
R35021 vdd.n16958 vdd.n16957 18.191
R35022 vdd.n16986 vdd.n16985 18.191
R35023 vdd.n17230 vdd.n17229 18.191
R35024 vdd.n17258 vdd.n17257 18.191
R35025 vdd.n17502 vdd.n17501 18.191
R35026 vdd.n17530 vdd.n17529 18.191
R35027 vdd.n17760 vdd.n17759 18.191
R35028 vdd.n17788 vdd.n17787 18.191
R35029 vdd.n18031 vdd.n18030 18.191
R35030 vdd.n18059 vdd.n18058 18.191
R35031 vdd.n18298 vdd.n18297 18.191
R35032 vdd.n15030 vdd.n15029 18.191
R35033 vdd.n15304 vdd.n15298 18.191
R35034 vdd.n15325 vdd.n15320 18.191
R35035 vdd.n15532 vdd.n15523 18.191
R35036 vdd.n15559 vdd.n15548 18.191
R35037 vdd.n15788 vdd.n15779 18.191
R35038 vdd.n15815 vdd.n15804 18.191
R35039 vdd.n16044 vdd.n16035 18.191
R35040 vdd.n16071 vdd.n16060 18.191
R35041 vdd.n16300 vdd.n16291 18.191
R35042 vdd.n16327 vdd.n16316 18.191
R35043 vdd.n16572 vdd.n16546 18.191
R35044 vdd.n13083 vdd.n9286 18.133
R35045 vdd.n9324 vdd.n9286 18.133
R35046 vdd.n9325 vdd.n9324 18.133
R35047 vdd.n13047 vdd.n9325 18.133
R35048 vdd.n13047 vdd.n13046 18.133
R35049 vdd.n13046 vdd.n13045 18.133
R35050 vdd.n13045 vdd.n9326 18.133
R35051 vdd.n13028 vdd.n9326 18.133
R35052 vdd.n13028 vdd.n13027 18.133
R35053 vdd.n13027 vdd.n13026 18.133
R35054 vdd.n13026 vdd.n9357 18.133
R35055 vdd.n9411 vdd.n9357 18.133
R35056 vdd.n12998 vdd.n9411 18.133
R35057 vdd.n12998 vdd.n12997 18.133
R35058 vdd.n12997 vdd.n12996 18.133
R35059 vdd.n12996 vdd.n9412 18.133
R35060 vdd.n9470 vdd.n9412 18.133
R35061 vdd.n9471 vdd.n9470 18.133
R35062 vdd.n12960 vdd.n9471 18.133
R35063 vdd.n12960 vdd.n12959 18.133
R35064 vdd.n12959 vdd.n12958 18.133
R35065 vdd.n12958 vdd.n9472 18.133
R35066 vdd.n9522 vdd.n9472 18.133
R35067 vdd.n12933 vdd.n9522 18.133
R35068 vdd.n12933 vdd.n12932 18.133
R35069 vdd.n12932 vdd.n12931 18.133
R35070 vdd.n12931 vdd.n9523 18.133
R35071 vdd.n9567 vdd.n9523 18.133
R35072 vdd.n12903 vdd.n9567 18.133
R35073 vdd.n12903 vdd.n12902 18.133
R35074 vdd.n12902 vdd.n12901 18.133
R35075 vdd.n12901 vdd.n9568 18.133
R35076 vdd.n9618 vdd.n9568 18.133
R35077 vdd.n12877 vdd.n9618 18.133
R35078 vdd.n12877 vdd.n12876 18.133
R35079 vdd.n12876 vdd.n12875 18.133
R35080 vdd.n12875 vdd.n9619 18.133
R35081 vdd.n9684 vdd.n9619 18.133
R35082 vdd.n9685 vdd.n9684 18.133
R35083 vdd.n12839 vdd.n9685 18.133
R35084 vdd.n12839 vdd.n12838 18.133
R35085 vdd.n12838 vdd.n12837 18.133
R35086 vdd.n12837 vdd.n9686 18.133
R35087 vdd.n12820 vdd.n9686 18.133
R35088 vdd.n12820 vdd.n12819 18.133
R35089 vdd.n12819 vdd.n12818 18.133
R35090 vdd.n12818 vdd.n9717 18.133
R35091 vdd.n9772 vdd.n9717 18.133
R35092 vdd.n12790 vdd.n9772 18.133
R35093 vdd.n12790 vdd.n12789 18.133
R35094 vdd.n12789 vdd.n12788 18.133
R35095 vdd.n12788 vdd.n9773 18.133
R35096 vdd.n9830 vdd.n9773 18.133
R35097 vdd.n9831 vdd.n9830 18.133
R35098 vdd.n12752 vdd.n9831 18.133
R35099 vdd.n12752 vdd.n12751 18.133
R35100 vdd.n12751 vdd.n12750 18.133
R35101 vdd.n12750 vdd.n9832 18.133
R35102 vdd.n9882 vdd.n9832 18.133
R35103 vdd.n12725 vdd.n9882 18.133
R35104 vdd.n12725 vdd.n12724 18.133
R35105 vdd.n12724 vdd.n12723 18.133
R35106 vdd.n12723 vdd.n9883 18.133
R35107 vdd.n9926 vdd.n9883 18.133
R35108 vdd.n12695 vdd.n9926 18.133
R35109 vdd.n12695 vdd.n12694 18.133
R35110 vdd.n12694 vdd.n12693 18.133
R35111 vdd.n12693 vdd.n9927 18.133
R35112 vdd.n9978 vdd.n9927 18.133
R35113 vdd.n12669 vdd.n9978 18.133
R35114 vdd.n12669 vdd.n12668 18.133
R35115 vdd.n12668 vdd.n12667 18.133
R35116 vdd.n12667 vdd.n9979 18.133
R35117 vdd.n10043 vdd.n9979 18.133
R35118 vdd.n10044 vdd.n10043 18.133
R35119 vdd.n12631 vdd.n10044 18.133
R35120 vdd.n12631 vdd.n12630 18.133
R35121 vdd.n12630 vdd.n12629 18.133
R35122 vdd.n12629 vdd.n10045 18.133
R35123 vdd.n12611 vdd.n10045 18.133
R35124 vdd.n12611 vdd.n12610 18.133
R35125 vdd.n12610 vdd.n12609 18.133
R35126 vdd.n12609 vdd.n10059 18.133
R35127 vdd.n10115 vdd.n10059 18.133
R35128 vdd.n12592 vdd.n10115 18.133
R35129 vdd.n12592 vdd.n12591 18.133
R35130 vdd.n12591 vdd.n12590 18.133
R35131 vdd.n12590 vdd.n10116 18.133
R35132 vdd.n10497 vdd.n10116 18.133
R35133 vdd.n12564 vdd.n10497 18.133
R35134 vdd.n12564 vdd.n12563 18.133
R35135 vdd.n12563 vdd.n12562 18.133
R35136 vdd.n12562 vdd.n10498 18.133
R35137 vdd.n12556 vdd.n10498 18.133
R35138 vdd.n12556 vdd.n12555 18.133
R35139 vdd.n12555 vdd.n12554 18.133
R35140 vdd.n12554 vdd.n10503 18.133
R35141 vdd.n12548 vdd.n10503 18.133
R35142 vdd.n12548 vdd.n12547 18.133
R35143 vdd.n12547 vdd.n12546 18.133
R35144 vdd.n12546 vdd.n10507 18.133
R35145 vdd.n12540 vdd.n10507 18.133
R35146 vdd.n12540 vdd.n12539 18.133
R35147 vdd.n12539 vdd.n12538 18.133
R35148 vdd.n12538 vdd.n10510 18.133
R35149 vdd.n12532 vdd.n10510 18.133
R35150 vdd.n12532 vdd.n12531 18.133
R35151 vdd.n12531 vdd.n12530 18.133
R35152 vdd.n12530 vdd.n10515 18.133
R35153 vdd.n12517 vdd.n10515 18.133
R35154 vdd.n12517 vdd.n12516 18.133
R35155 vdd.n12516 vdd.n12515 18.133
R35156 vdd.n12515 vdd.n10526 18.133
R35157 vdd.n10580 vdd.n10526 18.133
R35158 vdd.n12486 vdd.n10580 18.133
R35159 vdd.n12486 vdd.n12485 18.133
R35160 vdd.n12485 vdd.n12484 18.133
R35161 vdd.n12484 vdd.n10581 18.133
R35162 vdd.n10619 vdd.n10581 18.133
R35163 vdd.n12457 vdd.n10619 18.133
R35164 vdd.n12457 vdd.n12456 18.133
R35165 vdd.n12456 vdd.n12455 18.133
R35166 vdd.n12455 vdd.n10620 18.133
R35167 vdd.n10668 vdd.n10620 18.133
R35168 vdd.n12429 vdd.n10668 18.133
R35169 vdd.n12429 vdd.n12428 18.133
R35170 vdd.n12428 vdd.n12427 18.133
R35171 vdd.n12427 vdd.n10669 18.133
R35172 vdd.n10716 vdd.n10669 18.133
R35173 vdd.n12398 vdd.n10716 18.133
R35174 vdd.n12398 vdd.n12397 18.133
R35175 vdd.n12397 vdd.n12396 18.133
R35176 vdd.n12396 vdd.n10717 18.133
R35177 vdd.n10769 vdd.n10717 18.133
R35178 vdd.n10770 vdd.n10769 18.133
R35179 vdd.n12368 vdd.n10770 18.133
R35180 vdd.n12368 vdd.n12367 18.133
R35181 vdd.n12367 vdd.n12366 18.133
R35182 vdd.n12366 vdd.n10771 18.133
R35183 vdd.n10821 vdd.n10771 18.133
R35184 vdd.n12339 vdd.n10821 18.133
R35185 vdd.n12339 vdd.n12338 18.133
R35186 vdd.n12338 vdd.n12337 18.133
R35187 vdd.n12337 vdd.n10822 18.133
R35188 vdd.n12321 vdd.n10822 18.133
R35189 vdd.n12321 vdd.n12320 18.133
R35190 vdd.n12320 vdd.n12319 18.133
R35191 vdd.n12319 vdd.n10864 18.133
R35192 vdd.n10912 vdd.n10864 18.133
R35193 vdd.n12290 vdd.n10912 18.133
R35194 vdd.n12290 vdd.n12289 18.133
R35195 vdd.n12289 vdd.n12288 18.133
R35196 vdd.n12288 vdd.n10913 18.133
R35197 vdd.n10956 vdd.n10913 18.133
R35198 vdd.n12267 vdd.n10956 18.133
R35199 vdd.n12267 vdd.n12266 18.133
R35200 vdd.n12266 vdd.n12265 18.133
R35201 vdd.n12265 vdd.n10957 18.133
R35202 vdd.n11008 vdd.n10957 18.133
R35203 vdd.n12238 vdd.n11008 18.133
R35204 vdd.n12238 vdd.n12237 18.133
R35205 vdd.n12237 vdd.n12236 18.133
R35206 vdd.n12236 vdd.n11009 18.133
R35207 vdd.n11053 vdd.n11009 18.133
R35208 vdd.n12207 vdd.n11053 18.133
R35209 vdd.n12207 vdd.n12206 18.133
R35210 vdd.n12206 vdd.n12205 18.133
R35211 vdd.n12205 vdd.n11054 18.133
R35212 vdd.n11102 vdd.n11054 18.133
R35213 vdd.n12177 vdd.n11102 18.133
R35214 vdd.n12177 vdd.n12176 18.133
R35215 vdd.n12176 vdd.n12175 18.133
R35216 vdd.n12175 vdd.n11103 18.133
R35217 vdd.n11142 vdd.n11103 18.133
R35218 vdd.n12148 vdd.n11142 18.133
R35219 vdd.n12148 vdd.n12147 18.133
R35220 vdd.n12147 vdd.n12146 18.133
R35221 vdd.n12146 vdd.n11143 18.133
R35222 vdd.n11188 vdd.n11143 18.133
R35223 vdd.n12119 vdd.n11188 18.133
R35224 vdd.n12119 vdd.n12118 18.133
R35225 vdd.n12118 vdd.n12117 18.133
R35226 vdd.n12117 vdd.n11189 18.133
R35227 vdd.n11237 vdd.n11189 18.133
R35228 vdd.n12088 vdd.n11237 18.133
R35229 vdd.n12088 vdd.n12087 18.133
R35230 vdd.n12087 vdd.n12086 18.133
R35231 vdd.n12086 vdd.n11238 18.133
R35232 vdd.n11278 vdd.n11238 18.133
R35233 vdd.n12062 vdd.n11278 18.133
R35234 vdd.n12062 vdd.n12061 18.133
R35235 vdd.n12061 vdd.n12060 18.133
R35236 vdd.n12060 vdd.n11279 18.133
R35237 vdd.n11330 vdd.n11279 18.133
R35238 vdd.n12033 vdd.n11330 18.133
R35239 vdd.n12033 vdd.n12032 18.133
R35240 vdd.n12032 vdd.n12031 18.133
R35241 vdd.n12031 vdd.n11331 18.133
R35242 vdd.n12015 vdd.n11331 18.133
R35243 vdd.n12015 vdd.n12014 18.133
R35244 vdd.n12014 vdd.n12013 18.133
R35245 vdd.n12013 vdd.n11373 18.133
R35246 vdd.n11421 vdd.n11373 18.133
R35247 vdd.n11984 vdd.n11421 18.133
R35248 vdd.n11984 vdd.n11983 18.133
R35249 vdd.n11983 vdd.n11982 18.133
R35250 vdd.n11982 vdd.n11422 18.133
R35251 vdd.n11441 vdd.n11422 18.133
R35252 vdd.n11961 vdd.n11441 18.133
R35253 vdd.n11961 vdd.n11960 18.133
R35254 vdd.n11960 vdd.n11959 18.133
R35255 vdd.n11959 vdd.n11442 18.133
R35256 vdd.n11931 vdd.n11442 18.133
R35257 vdd.n11931 vdd.n11930 18.133
R35258 vdd.n11930 vdd.n11929 18.133
R35259 vdd.n11929 vdd.n11562 18.133
R35260 vdd.n11923 vdd.n11562 18.133
R35261 vdd.n15553 vdd.n15552 18.133
R35262 vdd.n15809 vdd.n15808 18.133
R35263 vdd.n16065 vdd.n16064 18.133
R35264 vdd.n16321 vdd.n16320 18.133
R35265 vdd.n16568 vdd.n16567 18.133
R35266 vdd.n16567 vdd.n16566 18.133
R35267 vdd.n16566 vdd.n16565 18.133
R35268 vdd.n16635 vdd.n16634 18.133
R35269 vdd.n16636 vdd.n16635 18.133
R35270 vdd.n16637 vdd.n16636 18.133
R35271 vdd.n16638 vdd.n16637 18.133
R35272 vdd.n15081 vdd.n15080 18.133
R35273 vdd.n15113 vdd.n15112 18.133
R35274 vdd.n15112 vdd.n15111 18.133
R35275 vdd.n15111 vdd.n15110 18.133
R35276 vdd.n15110 vdd.n15109 18.133
R35277 vdd.n15109 vdd.n15108 18.133
R35278 vdd.n15108 vdd.n15107 18.133
R35279 vdd.n15107 vdd.n15106 18.133
R35280 vdd.n15106 vdd.n15105 18.133
R35281 vdd.n15105 vdd.n15104 18.133
R35282 vdd.n16855 vdd.n16854 18.133
R35283 vdd.n16856 vdd.n16855 18.133
R35284 vdd.n16857 vdd.n16856 18.133
R35285 vdd.n16858 vdd.n16857 18.133
R35286 vdd.n16859 vdd.n16858 18.133
R35287 vdd.n16860 vdd.n16859 18.133
R35288 vdd.n16861 vdd.n16860 18.133
R35289 vdd.n16862 vdd.n16861 18.133
R35290 vdd.n14978 vdd.n14977 18.133
R35291 vdd.n14979 vdd.n14978 18.133
R35292 vdd.n14980 vdd.n14979 18.133
R35293 vdd.n14981 vdd.n14980 18.133
R35294 vdd.n14982 vdd.n14981 18.133
R35295 vdd.n14983 vdd.n14982 18.133
R35296 vdd.n14984 vdd.n14983 18.133
R35297 vdd.n14985 vdd.n14984 18.133
R35298 vdd.n14986 vdd.n14985 18.133
R35299 vdd.n14988 vdd.n14986 18.133
R35300 vdd.n14990 vdd.n14988 18.133
R35301 vdd.n14992 vdd.n14990 18.133
R35302 vdd.n14994 vdd.n14992 18.133
R35303 vdd.n14996 vdd.n14994 18.133
R35304 vdd.n14998 vdd.n14996 18.133
R35305 vdd.n15000 vdd.n14998 18.133
R35306 vdd.n15001 vdd.n15000 18.133
R35307 vdd.n11927 vdd.t186 17.972
R35308 vdd.t177 vdd.n21705 17.972
R35309 vdd.n35852 vdd.n35851 17.689
R35310 vdd.n35985 vdd.n35984 17.689
R35311 vdd.n36083 vdd.n36082 17.689
R35312 vdd.n36216 vdd.n36215 17.689
R35313 vdd.n36314 vdd.n36313 17.689
R35314 vdd.n36447 vdd.n36446 17.689
R35315 vdd.n36545 vdd.n36544 17.689
R35316 vdd.n36678 vdd.n36677 17.689
R35317 vdd.n36776 vdd.n36775 17.689
R35318 vdd.n36909 vdd.n36908 17.689
R35319 vdd.n37019 vdd.n37018 17.689
R35320 vdd.n33192 vdd.n33191 17.689
R35321 vdd.n37201 vdd.n37200 17.689
R35322 vdd.n33011 vdd.n33010 17.689
R35323 vdd.n32956 vdd.n32955 17.689
R35324 vdd.n37507 vdd.n37506 17.689
R35325 vdd.n38194 vdd.n38193 17.689
R35326 vdd.n38062 vdd.n38061 17.689
R35327 vdd.n37964 vdd.n37963 17.689
R35328 vdd.n37831 vdd.n37830 17.689
R35329 vdd.n37733 vdd.n37732 17.689
R35330 vdd.n37600 vdd.n37599 17.689
R35331 vdd.n28273 vdd.n28272 17.689
R35332 vdd.n28406 vdd.n28405 17.689
R35333 vdd.n28504 vdd.n28503 17.689
R35334 vdd.n28637 vdd.n28636 17.689
R35335 vdd.n28735 vdd.n28734 17.689
R35336 vdd.n28808 vdd.n28807 17.689
R35337 vdd.n28060 vdd.n28059 17.689
R35338 vdd.n31656 vdd.n31655 17.689
R35339 vdd.n27931 vdd.n27930 17.689
R35340 vdd.n29760 vdd.n29759 17.689
R35341 vdd.n30232 vdd.n30231 17.689
R35342 vdd.n30336 vdd.n30335 17.689
R35343 vdd.n2747 vdd.n2746 17.689
R35344 vdd.n2852 vdd.n2851 17.689
R35345 vdd.n2928 vdd.n2927 17.689
R35346 vdd.n3033 vdd.n3032 17.689
R35347 vdd.n3109 vdd.n3108 17.689
R35348 vdd.n3214 vdd.n3213 17.689
R35349 vdd.n3290 vdd.n3289 17.689
R35350 vdd.n3395 vdd.n3394 17.689
R35351 vdd.n3471 vdd.n3470 17.689
R35352 vdd.n3576 vdd.n3575 17.689
R35353 vdd.n3630 vdd.n3629 17.689
R35354 vdd.n3952 vdd.n3951 17.689
R35355 vdd.n2238 vdd.n2237 17.689
R35356 vdd.n2375 vdd.n2374 17.689
R35357 vdd.n2621 vdd.n2620 17.689
R35358 vdd.n1903 vdd.n1902 17.689
R35359 vdd.n1268 vdd.n1267 17.689
R35360 vdd.n1690 vdd.n1689 17.689
R35361 vdd.n1614 vdd.n1613 17.689
R35362 vdd.n1509 vdd.n1508 17.689
R35363 vdd.n1433 vdd.n1432 17.689
R35364 vdd.n1328 vdd.n1327 17.689
R35365 vdd.n26794 vdd.n26793 17.689
R35366 vdd.n26899 vdd.n26898 17.689
R35367 vdd.n26975 vdd.n26974 17.689
R35368 vdd.n27080 vdd.n27079 17.689
R35369 vdd.n27156 vdd.n27155 17.689
R35370 vdd.n26175 vdd.n26174 17.689
R35371 vdd.n31772 vdd.n31771 17.689
R35372 vdd.n31652 vdd.n31651 17.689
R35373 vdd.n32119 vdd.n32118 17.689
R35374 vdd.n31498 vdd.n31497 17.689
R35375 vdd.n32430 vdd.n32429 17.689
R35376 vdd.n31154 vdd.n31153 17.689
R35377 vdd.n13131 vdd.n9266 17.689
R35378 vdd.n13337 vdd.n9102 17.689
R35379 vdd.n13425 vdd.n9035 17.689
R35380 vdd.n13629 vdd.n8881 17.689
R35381 vdd.n13717 vdd.n8814 17.689
R35382 vdd.n8692 vdd.n8676 17.689
R35383 vdd.n14061 vdd.n8566 17.689
R35384 vdd.n8469 vdd.n8452 17.689
R35385 vdd.n14336 vdd.n8348 17.689
R35386 vdd.n14489 vdd.n8221 17.689
R35387 vdd.n14663 vdd.n8135 17.689
R35388 vdd.n14749 vdd.n8099 17.689
R35389 vdd.n14835 vdd.n8045 17.689
R35390 vdd.n14925 vdd.n8011 17.689
R35391 vdd.n13176 vdd.n9226 17.689
R35392 vdd.n13334 vdd.n9107 17.689
R35393 vdd.n13464 vdd.n9005 17.689
R35394 vdd.n13626 vdd.n8886 17.689
R35395 vdd.n13802 vdd.n8756 17.689
R35396 vdd.n13926 vdd.n8647 17.689
R35397 vdd.n14089 vdd.n8543 17.689
R35398 vdd.n14216 vdd.n8427 17.689
R35399 vdd.n8332 vdd.n8326 17.689
R35400 vdd.n14486 vdd.n8226 17.689
R35401 vdd.n19346 vdd.n19345 17.689
R35402 vdd.n19491 vdd.n19490 17.689
R35403 vdd.n19552 vdd.n19551 17.689
R35404 vdd.n19691 vdd.n19690 17.689
R35405 vdd.n19754 vdd.n19753 17.689
R35406 vdd.n20951 vdd.n20950 17.689
R35407 vdd.n20888 vdd.n20887 17.689
R35408 vdd.n20761 vdd.n20760 17.689
R35409 vdd.n20700 vdd.n20699 17.689
R35410 vdd.n20555 vdd.n20554 17.689
R35411 vdd.n21571 vdd.n21570 17.689
R35412 vdd.n21457 vdd.n21456 17.689
R35413 vdd.n21312 vdd.n21311 17.689
R35414 vdd.n21198 vdd.n21197 17.689
R35415 vdd.n21053 vdd.n21052 17.689
R35416 vdd.n19091 vdd.n19090 17.689
R35417 vdd.n18946 vdd.n18945 17.689
R35418 vdd.n18832 vdd.n18831 17.689
R35419 vdd.n18687 vdd.n18686 17.689
R35420 vdd.n18573 vdd.n18572 17.689
R35421 vdd.n20452 vdd.n20447 17.689
R35422 vdd.n20331 vdd.n20325 17.689
R35423 vdd.n20217 vdd.n20211 17.689
R35424 vdd.n20095 vdd.n20089 17.689
R35425 vdd.n24703 vdd.n24702 17.689
R35426 vdd.n25210 vdd.n25209 17.689
R35427 vdd.n24172 vdd.n24168 17.647
R35428 vdd.n24006 vdd.n24002 17.647
R35429 vdd.n23940 vdd.n23936 17.647
R35430 vdd.n23774 vdd.n23770 17.647
R35431 vdd.n23708 vdd.n23704 17.647
R35432 vdd.n23086 vdd.n23082 17.647
R35433 vdd.n23252 vdd.n23248 17.647
R35434 vdd.n23318 vdd.n23314 17.647
R35435 vdd.n23484 vdd.n23480 17.647
R35436 vdd.n23550 vdd.n23546 17.647
R35437 vdd.n22507 vdd.n22503 17.647
R35438 vdd.n22673 vdd.n22669 17.647
R35439 vdd.n22739 vdd.n22735 17.647
R35440 vdd.n22905 vdd.n22901 17.647
R35441 vdd.n22971 vdd.n22967 17.647
R35442 vdd.n22447 vdd.n22443 17.647
R35443 vdd.n22252 vdd.n22247 17.647
R35444 vdd.n22303 vdd.n22299 17.647
R35445 vdd.n22128 vdd.n22123 17.647
R35446 vdd.n24275 vdd.n24271 17.647
R35447 vdd.n12528 vdd.n12527 17.331
R35448 vdd.n16869 vdd.n16864 17.331
R35449 vdd.n10276 vdd.n10272 17.102
R35450 vdd.n10467 vdd.n10466 17.102
R35451 vdd.n10455 vdd.n10279 17.102
R35452 vdd.n10453 vdd.n10290 17.102
R35453 vdd.n10443 vdd.n10442 17.102
R35454 vdd.n10431 vdd.n10297 17.102
R35455 vdd.n10429 vdd.n10307 17.102
R35456 vdd.n10417 vdd.n10319 17.102
R35457 vdd.n10415 vdd.n10320 17.102
R35458 vdd.n10404 vdd.n10403 17.102
R35459 vdd.n10394 vdd.n10392 17.102
R35460 vdd.n15303 vdd.n15302 17.102
R35461 vdd.n15324 vdd.n15321 17.102
R35462 vdd.n10247 vdd.n10227 17.066
R35463 vdd.n10234 vdd.n10231 17.066
R35464 vdd.n10379 vdd.n10344 17.01
R35465 vdd.n10370 vdd.n10369 17.01
R35466 vdd.n12521 vdd.n12520 17.01
R35467 vdd.n10552 vdd.n10523 17.01
R35468 vdd.n10554 vdd.n10528 17.01
R35469 vdd.n12503 vdd.n10529 17.01
R35470 vdd.n12501 vdd.n10564 17.01
R35471 vdd.n12489 vdd.n10573 17.01
R35472 vdd.n12472 vdd.n10584 17.01
R35473 vdd.n12470 vdd.n10605 17.01
R35474 vdd.n12461 vdd.n12460 17.01
R35475 vdd.n10645 vdd.n10615 17.01
R35476 vdd.n10647 vdd.n10622 17.01
R35477 vdd.n12443 vdd.n10623 17.01
R35478 vdd.n12441 vdd.n10656 17.01
R35479 vdd.n10690 vdd.n10671 17.01
R35480 vdd.n12415 vdd.n10672 17.01
R35481 vdd.n12401 vdd.n10708 17.01
R35482 vdd.n10737 vdd.n10709 17.01
R35483 vdd.n10739 vdd.n10719 17.01
R35484 vdd.n12384 vdd.n10720 17.01
R35485 vdd.n12382 vdd.n10749 17.01
R35486 vdd.n12372 vdd.n12371 17.01
R35487 vdd.n10796 vdd.n10764 17.01
R35488 vdd.n10798 vdd.n10773 17.01
R35489 vdd.n12352 vdd.n10807 17.01
R35490 vdd.n10844 vdd.n10817 17.01
R35491 vdd.n12324 vdd.n10861 17.01
R35492 vdd.n10884 vdd.n10862 17.01
R35493 vdd.n10886 vdd.n10866 17.01
R35494 vdd.n12307 vdd.n10867 17.01
R35495 vdd.n12305 vdd.n10896 17.01
R35496 vdd.n12293 vdd.n10905 17.01
R35497 vdd.n12286 vdd.n10915 17.01
R35498 vdd.n12271 vdd.n12270 17.01
R35499 vdd.n10983 vdd.n10952 17.01
R35500 vdd.n10985 vdd.n10959 17.01
R35501 vdd.n12251 vdd.n10994 17.01
R35502 vdd.n12242 vdd.n12241 17.01
R35503 vdd.n12224 vdd.n11012 17.01
R35504 vdd.n12210 vdd.n11045 17.01
R35505 vdd.n11074 vdd.n11046 17.01
R35506 vdd.n11076 vdd.n11056 17.01
R35507 vdd.n12193 vdd.n11057 17.01
R35508 vdd.n12191 vdd.n11086 17.01
R35509 vdd.n12179 vdd.n11095 17.01
R35510 vdd.n11119 vdd.n11105 17.01
R35511 vdd.n12163 vdd.n11106 17.01
R35512 vdd.n12161 vdd.n11128 17.01
R35513 vdd.n12152 vdd.n12151 17.01
R35514 vdd.n11168 vdd.n11138 17.01
R35515 vdd.t298 vdd.n11145 17.01
R35516 vdd.n12134 vdd.n11146 17.01
R35517 vdd.n11209 vdd.n11185 17.01
R35518 vdd.n11211 vdd.n11191 17.01
R35519 vdd.n12105 vdd.n11192 17.01
R35520 vdd.n12103 vdd.n11221 17.01
R35521 vdd.n12091 vdd.n11230 17.01
R35522 vdd.n11258 vdd.n11231 17.01
R35523 vdd.n11260 vdd.n11240 17.01
R35524 vdd.n12074 vdd.n11241 17.01
R35525 vdd.n12066 vdd.n12065 17.01
R35526 vdd.n11305 vdd.n11274 17.01
R35527 vdd.n12048 vdd.n11282 17.01
R35528 vdd.n12046 vdd.n11316 17.01
R35529 vdd.n12037 vdd.n12036 17.01
R35530 vdd.n11353 vdd.n11326 17.01
R35531 vdd.n12018 vdd.n11370 17.01
R35532 vdd.n11393 vdd.n11371 17.01
R35533 vdd.n11395 vdd.n11375 17.01
R35534 vdd.n11999 vdd.n11405 17.01
R35535 vdd.n11481 vdd.n11414 17.01
R35536 vdd.n11980 vdd.n11424 17.01
R35537 vdd.n11972 vdd.n11971 17.01
R35538 vdd.n11965 vdd.n11964 17.01
R35539 vdd.n11527 vdd.n11444 17.01
R35540 vdd.n11946 vdd.n11445 17.01
R35541 vdd.n11944 vdd.n11549 17.01
R35542 vdd.n15010 vdd.n15009 17.01
R35543 vdd.n19267 vdd.t140 17.006
R35544 vdd.n19933 vdd.t150 17.006
R35545 vdd.n12526 vdd.n10519 16.978
R35546 vdd.n12440 vdd.n10655 16.978
R35547 vdd.n12424 vdd.n10673 16.978
R35548 vdd.n10842 vdd.n10818 16.978
R35549 vdd.n12325 vdd.n10857 16.978
R35550 vdd.n12243 vdd.n11001 16.978
R35551 vdd.n12225 vdd.n11036 16.978
R35552 vdd.n12143 vdd.n11148 16.978
R35553 vdd.n11208 vdd.n11199 16.978
R35554 vdd.n11351 vdd.n11327 16.978
R35555 vdd.n12019 vdd.n11366 16.978
R35556 vdd.n11934 vdd.n11559 16.978
R35557 vdd.n10391 vdd.n10390 16.978
R35558 vdd.n10355 vdd.n10345 16.978
R35559 vdd.n9443 vdd.n9432 16.978
R35560 vdd.n12983 vdd.n9420 16.978
R35561 vdd.n9606 vdd.n9573 16.978
R35562 vdd.n9636 vdd.n9631 16.978
R35563 vdd.n9802 vdd.n9792 16.978
R35564 vdd.n12775 vdd.n9781 16.978
R35565 vdd.n9966 vdd.n9932 16.978
R35566 vdd.n9996 vdd.n9991 16.978
R35567 vdd.n10245 vdd.n10237 16.978
R35568 vdd.n10488 vdd.n10481 16.978
R35569 vdd.n16870 vdd.n16837 16.978
R35570 vdd.n17088 vdd.n17082 16.978
R35571 vdd.n17140 vdd.n17134 16.978
R35572 vdd.n17360 vdd.n17354 16.978
R35573 vdd.n17412 vdd.n17406 16.978
R35574 vdd.n17618 vdd.n17612 16.978
R35575 vdd.n17670 vdd.n17664 16.978
R35576 vdd.n17889 vdd.n17883 16.978
R35577 vdd.n17941 vdd.n17935 16.978
R35578 vdd.n18161 vdd.n18155 16.978
R35579 vdd.n18213 vdd.n18207 16.978
R35580 vdd.n15014 vdd.n15013 16.978
R35581 vdd.n15406 vdd.n15405 16.978
R35582 vdd.n15424 vdd.n15423 16.978
R35583 vdd.n15654 vdd.n15653 16.978
R35584 vdd.n15674 vdd.n15673 16.978
R35585 vdd.n15910 vdd.n15909 16.978
R35586 vdd.n15930 vdd.n15929 16.978
R35587 vdd.n16166 vdd.n16165 16.978
R35588 vdd.n16186 vdd.n16185 16.978
R35589 vdd.n16422 vdd.n16421 16.978
R35590 vdd.n16442 vdd.n16441 16.978
R35591 vdd.n16607 vdd.n16606 16.978
R35592 vdd.n15077 vdd.n15076 16.978
R35593 vdd.t313 vdd.n8083 16.964
R35594 vdd.t312 vdd.n8054 16.964
R35595 vdd.n24185 vdd.n24184 16.964
R35596 vdd.n23991 vdd.n23990 16.964
R35597 vdd.n23953 vdd.n23952 16.964
R35598 vdd.n23759 vdd.n23758 16.964
R35599 vdd.n23721 vdd.n23720 16.964
R35600 vdd.n23071 vdd.n23070 16.964
R35601 vdd.n23265 vdd.n23264 16.964
R35602 vdd.n23303 vdd.n23302 16.964
R35603 vdd.n23497 vdd.n23496 16.964
R35604 vdd.n23535 vdd.n23534 16.964
R35605 vdd.n22492 vdd.n22491 16.964
R35606 vdd.n22686 vdd.n22685 16.964
R35607 vdd.n22724 vdd.n22723 16.964
R35608 vdd.n22918 vdd.n22917 16.964
R35609 vdd.n22956 vdd.n22955 16.964
R35610 vdd.n22462 vdd.n22461 16.964
R35611 vdd.n22333 vdd.n22332 16.964
R35612 vdd.n22318 vdd.n22317 16.964
R35613 vdd.n22135 vdd.n22134 16.964
R35614 vdd.n24290 vdd.n24289 16.964
R35615 vdd.n10389 vdd.n10388 16.943
R35616 vdd.n21669 vdd.t245 16.888
R35617 vdd.n12432 vdd.n12431 16.689
R35618 vdd.n12335 vdd.n10824 16.689
R35619 vdd.n12335 vdd.n10825 16.689
R35620 vdd.n11028 vdd.n11004 16.689
R35621 vdd.n11028 vdd.n11011 16.689
R35622 vdd.n12122 vdd.n11184 16.689
R35623 vdd.n12029 vdd.n11333 16.689
R35624 vdd.n12029 vdd.n11334 16.689
R35625 vdd.n17395 vdd.n17390 16.689
R35626 vdd.n17653 vdd.n17648 16.689
R35627 vdd.n17924 vdd.n17919 16.689
R35628 vdd.n18196 vdd.n18191 16.689
R35629 vdd.n9277 vdd.n9244 16.632
R35630 vdd.t306 vdd.n10906 16.368
R35631 vdd.n11927 vdd.n11564 16.368
R35632 vdd.n21705 vdd.n21704 16.368
R35633 vdd.n14549 vdd.n8188 16.21
R35634 vdd.n14646 vdd.n8146 16.21
R35635 vdd.n8160 vdd.n8140 16.21
R35636 vdd.n21414 vdd.t325 16.185
R35637 vdd.n18740 vdd.t274 16.185
R35638 vdd.n10500 vdd.t381 16.047
R35639 vdd.n10710 vdd.t357 16.047
R35640 vdd.t0 vdd.n15103 16.047
R35641 vdd.n24849 vdd.t204 15.921
R35642 vdd.n14567 vdd.n8172 15.904
R35643 vdd.n11733 vdd.n11732 15.779
R35644 vdd.n21808 vdd.n21807 15.779
R35645 vdd.n11833 vdd.n11832 15.779
R35646 vdd.n21924 vdd.n21923 15.779
R35647 vdd.n10576 vdd.n10571 15.765
R35648 vdd.n12473 vdd.n10604 15.765
R35649 vdd.n12393 vdd.n10722 15.765
R35650 vdd.n10765 vdd.n10756 15.765
R35651 vdd.n10928 vdd.n10904 15.765
R35652 vdd.n12276 vdd.n10923 15.765
R35653 vdd.n12190 vdd.n11085 15.765
R35654 vdd.n12172 vdd.n11107 15.765
R35655 vdd.n11261 vdd.n11248 15.765
R35656 vdd.n11275 vdd.n11272 15.765
R35657 vdd.n11472 vdd.n11413 15.765
R35658 vdd.n11970 vdd.n11432 15.765
R35659 vdd.n10464 vdd.n10280 15.765
R35660 vdd.n10432 vdd.n10306 15.765
R35661 vdd.n13051 vdd.n9315 15.765
R35662 vdd.n9375 vdd.n9369 15.765
R35663 vdd.n12950 vdd.n9477 15.765
R35664 vdd.n12927 vdd.n9527 15.765
R35665 vdd.n12843 vdd.n9676 15.765
R35666 vdd.n9735 vdd.n9729 15.765
R35667 vdd.n12742 vdd.n9837 15.765
R35668 vdd.n12719 vdd.n9888 15.765
R35669 vdd.n12635 vdd.n10036 15.765
R35670 vdd.n10141 vdd.n10140 15.765
R35671 vdd.n16942 vdd.n16941 15.765
R35672 vdd.n17002 vdd.n17001 15.765
R35673 vdd.n17214 vdd.n17213 15.765
R35674 vdd.n17274 vdd.n17273 15.765
R35675 vdd.n17486 vdd.n17485 15.765
R35676 vdd.n17546 vdd.n17545 15.765
R35677 vdd.n17744 vdd.n17743 15.765
R35678 vdd.n17804 vdd.n17803 15.765
R35679 vdd.n18015 vdd.n18014 15.765
R35680 vdd.n18075 vdd.n18074 15.765
R35681 vdd.n18283 vdd.n18282 15.765
R35682 vdd.n18323 vdd.n18322 15.765
R35683 vdd.n15288 vdd.n15284 15.765
R35684 vdd.n15339 vdd.n15335 15.765
R35685 vdd.n15513 vdd.n15506 15.765
R35686 vdd.n15576 vdd.n15569 15.765
R35687 vdd.n15769 vdd.n15762 15.765
R35688 vdd.n15832 vdd.n15825 15.765
R35689 vdd.n16025 vdd.n16018 15.765
R35690 vdd.n16088 vdd.n16081 15.765
R35691 vdd.n16281 vdd.n16274 15.765
R35692 vdd.n16344 vdd.n16337 15.765
R35693 vdd.n16537 vdd.n16530 15.765
R35694 vdd.n35856 vdd.n35852 15.724
R35695 vdd.n35989 vdd.n35985 15.724
R35696 vdd.n36087 vdd.n36083 15.724
R35697 vdd.n36220 vdd.n36216 15.724
R35698 vdd.n36318 vdd.n36314 15.724
R35699 vdd.n36451 vdd.n36447 15.724
R35700 vdd.n36549 vdd.n36545 15.724
R35701 vdd.n36682 vdd.n36678 15.724
R35702 vdd.n36780 vdd.n36776 15.724
R35703 vdd.n36913 vdd.n36909 15.724
R35704 vdd.n37020 vdd.n37019 15.724
R35705 vdd.n33196 vdd.n33192 15.724
R35706 vdd.n37205 vdd.n37201 15.724
R35707 vdd.n33012 vdd.n33011 15.724
R35708 vdd.n32960 vdd.n32956 15.724
R35709 vdd.n37508 vdd.n37507 15.724
R35710 vdd.n38195 vdd.n38194 15.724
R35711 vdd.n38066 vdd.n38062 15.724
R35712 vdd.n37968 vdd.n37964 15.724
R35713 vdd.n37835 vdd.n37831 15.724
R35714 vdd.n37737 vdd.n37733 15.724
R35715 vdd.n37604 vdd.n37600 15.724
R35716 vdd.n28277 vdd.n28273 15.724
R35717 vdd.n28410 vdd.n28406 15.724
R35718 vdd.n28508 vdd.n28504 15.724
R35719 vdd.n28641 vdd.n28637 15.724
R35720 vdd.n28739 vdd.n28735 15.724
R35721 vdd.n28812 vdd.n28808 15.724
R35722 vdd.n28064 vdd.n28060 15.724
R35723 vdd.n31657 vdd.n31656 15.724
R35724 vdd.n27932 vdd.n27931 15.724
R35725 vdd.n29764 vdd.n29760 15.724
R35726 vdd.n30236 vdd.n30232 15.724
R35727 vdd.n30340 vdd.n30336 15.724
R35728 vdd.n2748 vdd.n2747 15.724
R35729 vdd.n2853 vdd.n2852 15.724
R35730 vdd.n2929 vdd.n2928 15.724
R35731 vdd.n3034 vdd.n3033 15.724
R35732 vdd.n3110 vdd.n3109 15.724
R35733 vdd.n3215 vdd.n3214 15.724
R35734 vdd.n3291 vdd.n3290 15.724
R35735 vdd.n3396 vdd.n3395 15.724
R35736 vdd.n3472 vdd.n3471 15.724
R35737 vdd.n3577 vdd.n3576 15.724
R35738 vdd.n3634 vdd.n3630 15.724
R35739 vdd.n3953 vdd.n3952 15.724
R35740 vdd.n2239 vdd.n2238 15.724
R35741 vdd.n2379 vdd.n2375 15.724
R35742 vdd.n2622 vdd.n2621 15.724
R35743 vdd.n1907 vdd.n1903 15.724
R35744 vdd.n1272 vdd.n1268 15.724
R35745 vdd.n1691 vdd.n1690 15.724
R35746 vdd.n1615 vdd.n1614 15.724
R35747 vdd.n1510 vdd.n1509 15.724
R35748 vdd.n1434 vdd.n1433 15.724
R35749 vdd.n1329 vdd.n1328 15.724
R35750 vdd.n26795 vdd.n26794 15.724
R35751 vdd.n26900 vdd.n26899 15.724
R35752 vdd.n26976 vdd.n26975 15.724
R35753 vdd.n27081 vdd.n27080 15.724
R35754 vdd.n27157 vdd.n27156 15.724
R35755 vdd.n26176 vdd.n26175 15.724
R35756 vdd.n31773 vdd.n31772 15.724
R35757 vdd.n31659 vdd.n31652 15.724
R35758 vdd.n32123 vdd.n32119 15.724
R35759 vdd.n31499 vdd.n31498 15.724
R35760 vdd.n32431 vdd.n32430 15.724
R35761 vdd.n31155 vdd.n31154 15.724
R35762 vdd.n13127 vdd.n9266 15.724
R35763 vdd.n13294 vdd.n9102 15.724
R35764 vdd.n13421 vdd.n9035 15.724
R35765 vdd.n13586 vdd.n8881 15.724
R35766 vdd.n13713 vdd.n8814 15.724
R35767 vdd.n13890 vdd.n8692 15.724
R35768 vdd.n14061 vdd.n8567 15.724
R35769 vdd.n14179 vdd.n8469 15.724
R35770 vdd.n14336 vdd.n8349 15.724
R35771 vdd.n8253 vdd.n8221 15.724
R35772 vdd.n14663 vdd.n8139 15.724
R35773 vdd.n14749 vdd.n8095 15.724
R35774 vdd.n14835 vdd.n8049 15.724
R35775 vdd.n14925 vdd.n8007 15.724
R35776 vdd.n13169 vdd.n9226 15.724
R35777 vdd.n13330 vdd.n9107 15.724
R35778 vdd.n13471 vdd.n9005 15.724
R35779 vdd.n13622 vdd.n8886 15.724
R35780 vdd.n13802 vdd.n8755 15.724
R35781 vdd.n13926 vdd.n8648 15.724
R35782 vdd.n14089 vdd.n8542 15.724
R35783 vdd.n14216 vdd.n8428 15.724
R35784 vdd.n14363 vdd.n8326 15.724
R35785 vdd.n14482 vdd.n8226 15.724
R35786 vdd.n19352 vdd.n19346 15.724
R35787 vdd.n19497 vdd.n19491 15.724
R35788 vdd.n19558 vdd.n19552 15.724
R35789 vdd.n19697 vdd.n19691 15.724
R35790 vdd.n19760 vdd.n19754 15.724
R35791 vdd.n20957 vdd.n20951 15.724
R35792 vdd.n20894 vdd.n20888 15.724
R35793 vdd.n20767 vdd.n20761 15.724
R35794 vdd.n20706 vdd.n20700 15.724
R35795 vdd.n20561 vdd.n20555 15.724
R35796 vdd.n21577 vdd.n21571 15.724
R35797 vdd.n21463 vdd.n21457 15.724
R35798 vdd.n21318 vdd.n21312 15.724
R35799 vdd.n21204 vdd.n21198 15.724
R35800 vdd.n21059 vdd.n21053 15.724
R35801 vdd.n19097 vdd.n19091 15.724
R35802 vdd.n18952 vdd.n18946 15.724
R35803 vdd.n18838 vdd.n18832 15.724
R35804 vdd.n18693 vdd.n18687 15.724
R35805 vdd.n18579 vdd.n18573 15.724
R35806 vdd.n20447 vdd.n20446 15.724
R35807 vdd.n20325 vdd.n20324 15.724
R35808 vdd.n20211 vdd.n20210 15.724
R35809 vdd.n20089 vdd.n20088 15.724
R35810 vdd.n24790 vdd.n24789 15.724
R35811 vdd.n25119 vdd.n25118 15.724
R35812 vdd.n9185 vdd.n9170 15.598
R35813 vdd.n9056 vdd.n9055 15.598
R35814 vdd.n8964 vdd.n8950 15.598
R35815 vdd.n13537 vdd.n8958 15.598
R35816 vdd.n13669 vdd.n13668 15.598
R35817 vdd.n8738 vdd.n8731 15.598
R35818 vdd.n13822 vdd.n8712 15.598
R35819 vdd.n13975 vdd.n8593 15.598
R35820 vdd.n14108 vdd.n8524 15.598
R35821 vdd.n14126 vdd.n8489 15.598
R35822 vdd.n14250 vdd.n8408 15.598
R35823 vdd.n14420 vdd.n8285 15.598
R35824 vdd.n21009 vdd.n21000 15.481
R35825 vdd.n11923 vdd.n11922 15.466
R35826 vdd.n15002 vdd.n15001 15.466
R35827 vdd.n24791 vdd.n24790 15.438
R35828 vdd.n25120 vdd.n25119 15.438
R35829 vdd.n12431 vdd.t314 15.405
R35830 ldomc_0.otaldom_0.pmoslm_0.vdd vdd.n10960 15.405
R35831 vdd.t257 vdd.n17118 15.405
R35832 bandgapmd_0.otam_1.pmoslm_0.vdd vdd.n17596 15.405
R35833 vdd.n13245 vdd.t289 15.292
R35834 vdd.n14531 vdd.n14530 15.292
R35835 vdd.n10263 vdd.n10262 15.094
R35836 vdd.n14408 vdd.t317 14.987
R35837 vdd.n33533 vdd.n33532 14.919
R35838 vdd.n34272 vdd.n34271 14.919
R35839 vdd.n33925 vdd.n33924 14.919
R35840 vdd.n35416 vdd.n35415 14.919
R35841 vdd.n35538 vdd.n35537 14.919
R35842 vdd.n34927 vdd.n34926 14.919
R35843 vdd.n34820 vdd.n34819 14.919
R35844 vdd.n645 vdd.n644 14.919
R35845 vdd.n413 vdd.n412 14.919
R35846 vdd.n6199 vdd.n6198 14.919
R35847 vdd.n5970 vdd.n5969 14.919
R35848 vdd.n5674 vdd.n5673 14.919
R35849 vdd.n5567 vdd.n5566 14.919
R35850 vdd.n5000 vdd.n4999 14.919
R35851 vdd.n5111 vdd.n5110 14.919
R35852 vdd.n4501 vdd.n4500 14.919
R35853 vdd.n4393 vdd.n4392 14.919
R35854 vdd.n27417 vdd.n27416 14.919
R35855 vdd.n27523 vdd.n27522 14.919
R35856 vdd.n25863 vdd.n25862 14.919
R35857 vdd.n25960 vdd.n25959 14.919
R35858 vdd.n26748 vdd.n26747 14.772
R35859 vdd.n38126 vdd.n38116 14.771
R35860 vdd.n28156 vdd.n28155 14.771
R35861 vdd.n1740 vdd.n1733 14.771
R35862 vdd.n14611 vdd.n8169 14.682
R35863 vdd.n11579 vdd.n11576 14.682
R35864 vdd.n10524 vdd.n10522 14.553
R35865 vdd.n12452 vdd.n10625 14.553
R35866 vdd.n12416 vdd.n10699 14.553
R35867 vdd.n12344 vdd.n10814 14.553
R35868 vdd.n10883 vdd.n10874 14.553
R35869 vdd.n12250 vdd.n10993 14.553
R35870 vdd.n11049 vdd.n11037 14.553
R35871 vdd.n11170 vdd.n11154 14.553
R35872 vdd.n12114 vdd.n11193 14.553
R35873 vdd.n12038 vdd.n11323 14.553
R35874 vdd.n11392 vdd.n11383 14.553
R35875 vdd.n11943 vdd.n11548 14.553
R35876 vdd.n10336 vdd.n10327 14.553
R35877 vdd.n10367 vdd.n10356 14.553
R35878 vdd.n13003 vdd.n13002 14.553
R35879 vdd.n12975 vdd.n9453 14.553
R35880 vdd.n9597 vdd.n9572 14.553
R35881 vdd.n9650 vdd.n9629 14.553
R35882 vdd.n12795 vdd.n12794 14.553
R35883 vdd.n12767 vdd.n9812 14.553
R35884 vdd.n9957 vdd.n9931 14.553
R35885 vdd.n10010 vdd.n9989 14.553
R35886 vdd.n12596 vdd.n10101 14.553
R35887 vdd.n10492 vdd.n10270 14.553
R35888 vdd.n16884 vdd.n16878 14.553
R35889 vdd.n17072 vdd.n17066 14.553
R35890 vdd.n17156 vdd.n17150 14.553
R35891 vdd.n17344 vdd.n17338 14.553
R35892 vdd.n17428 vdd.n17422 14.553
R35893 vdd.n17602 vdd.n16823 14.553
R35894 vdd.n17686 vdd.n17680 14.553
R35895 vdd.n17873 vdd.n17868 14.553
R35896 vdd.n17957 vdd.n17951 14.553
R35897 vdd.n18145 vdd.n18139 14.553
R35898 vdd.n18228 vdd.n18223 14.553
R35899 vdd.n18398 vdd.n18397 14.553
R35900 vdd.n15392 vdd.n15391 14.553
R35901 vdd.n15438 vdd.n15437 14.553
R35902 vdd.n15637 vdd.n15636 14.553
R35903 vdd.n15691 vdd.n15690 14.553
R35904 vdd.n15893 vdd.n15892 14.553
R35905 vdd.n15947 vdd.n15946 14.553
R35906 vdd.n16149 vdd.n16148 14.553
R35907 vdd.n16203 vdd.n16202 14.553
R35908 vdd.n16405 vdd.n16404 14.553
R35909 vdd.n16459 vdd.n16458 14.553
R35910 vdd.n16630 vdd.n16629 14.553
R35911 vdd.n15071 vdd.n15070 14.553
R35912 vdd.n24981 vdd.n24980 14.493
R35913 vdd.n24980 vdd.n24979 14.493
R35914 vdd.t375 vdd.n11281 14.442
R35915 vdd.n11415 vdd.t364 14.442
R35916 vdd.t295 vdd.n10290 14.198
R35917 vdd.n24112 vdd.n24111 14.117
R35918 vdd.n24058 vdd.n24057 14.117
R35919 vdd.n23880 vdd.n23879 14.117
R35920 vdd.n23826 vdd.n23825 14.117
R35921 vdd.n23648 vdd.n23647 14.117
R35922 vdd.n23138 vdd.n23137 14.117
R35923 vdd.n23192 vdd.n23191 14.117
R35924 vdd.n23370 vdd.n23369 14.117
R35925 vdd.n23424 vdd.n23423 14.117
R35926 vdd.n23602 vdd.n23601 14.117
R35927 vdd.n22559 vdd.n22558 14.117
R35928 vdd.n22613 vdd.n22612 14.117
R35929 vdd.n22791 vdd.n22790 14.117
R35930 vdd.n22845 vdd.n22844 14.117
R35931 vdd.n23023 vdd.n23022 14.117
R35932 vdd.n22386 vdd.n22385 14.117
R35933 vdd.n22354 vdd.n22353 14.117
R35934 vdd.n24331 vdd.n24330 14.117
R35935 vdd.n22083 vdd.n22082 14.117
R35936 vdd.n24214 vdd.n24213 14.117
R35937 vdd.n8984 vdd.n8983 14.085
R35938 vdd.n13541 vdd.n13540 14.085
R35939 vdd.n13789 vdd.n8769 14.085
R35940 vdd.n13826 vdd.n13825 14.085
R35941 vdd.n8555 vdd.n8515 14.085
R35942 vdd.n8519 vdd.n8507 14.085
R35943 vdd.n20282 vdd.t255 14.074
R35944 vdd.n20264 vdd.t272 14.074
R35945 vdd.n8087 vdd.t313 14.039
R35946 vdd.n14802 vdd.t312 14.039
R35947 vdd.n14704 vdd.n8117 13.914
R35948 vdd.n14705 vdd.n8115 13.914
R35949 vdd.n14854 vdd.n8028 13.914
R35950 vdd.n14878 vdd.n8026 13.914
R35951 vdd.n11790 vdd.t373 13.847
R35952 vdd.n11790 vdd.t382 13.847
R35953 vdd.n11780 vdd.t358 13.847
R35954 vdd.n11780 vdd.t380 13.847
R35955 vdd.n11673 vdd.t384 13.847
R35956 vdd.n11673 vdd.t376 13.847
R35957 vdd.n11667 vdd.t386 13.847
R35958 vdd.n11667 vdd.t378 13.847
R35959 vdd.n11715 vdd.n11689 13.847
R35960 vdd.n11715 vdd.t187 13.847
R35961 vdd.n11688 vdd.t365 13.847
R35962 vdd.n11689 vdd.n11688 13.847
R35963 vdd.n11792 vdd.t388 13.847
R35964 vdd.n11792 vdd.t354 13.847
R35965 vdd.n11837 vdd.n11834 13.847
R35966 vdd.n11837 vdd.n11836 13.847
R35967 vdd.n11883 vdd.t367 13.847
R35968 vdd.n11883 vdd.t356 13.847
R35969 vdd.n11836 vdd.n11835 13.847
R35970 vdd.n11835 vdd.t361 13.847
R35971 vdd.n11910 vdd.t363 13.847
R35972 vdd.n11910 vdd.t369 13.847
R35973 vdd.n21881 vdd.t15 13.847
R35974 vdd.n21881 vdd.t1 13.847
R35975 vdd.n21870 vdd.t9 13.847
R35976 vdd.n21870 vdd.t26 13.847
R35977 vdd.n21849 vdd.t31 13.847
R35978 vdd.n21849 vdd.t13 13.847
R35979 vdd.n21860 vdd.t5 13.847
R35980 vdd.n21860 vdd.t11 13.847
R35981 vdd.n21764 vdd.t178 13.847
R35982 vdd.n21760 vdd.t33 13.847
R35983 vdd.n21760 vdd.n21759 13.847
R35984 vdd.n21883 vdd.t3 13.847
R35985 vdd.n21883 vdd.t17 13.847
R35986 vdd.n21928 vdd.n21925 13.847
R35987 vdd.n21928 vdd.n21927 13.847
R35988 vdd.n21974 vdd.t35 13.847
R35989 vdd.n21974 vdd.t19 13.847
R35990 vdd.n21927 vdd.n21926 13.847
R35991 vdd.n21926 vdd.t29 13.847
R35992 vdd.n21999 vdd.t7 13.847
R35993 vdd.n21999 vdd.t21 13.847
R35994 vdd.n35866 vdd.n35865 13.758
R35995 vdd.n35971 vdd.n35970 13.758
R35996 vdd.n36097 vdd.n36096 13.758
R35997 vdd.n36202 vdd.n36201 13.758
R35998 vdd.n36328 vdd.n36327 13.758
R35999 vdd.n36433 vdd.n36432 13.758
R36000 vdd.n36559 vdd.n36558 13.758
R36001 vdd.n36664 vdd.n36663 13.758
R36002 vdd.n36790 vdd.n36789 13.758
R36003 vdd.n36895 vdd.n36894 13.758
R36004 vdd.n37038 vdd.n37037 13.758
R36005 vdd.n37111 vdd.n37110 13.758
R36006 vdd.n33112 vdd.n33111 13.758
R36007 vdd.n33033 vdd.n33032 13.758
R36008 vdd.n37404 vdd.n37403 13.758
R36009 vdd.n32866 vdd.n32865 13.758
R36010 vdd.n38180 vdd.n38179 13.758
R36011 vdd.n38076 vdd.n38075 13.758
R36012 vdd.n37950 vdd.n37949 13.758
R36013 vdd.n37845 vdd.n37844 13.758
R36014 vdd.n37719 vdd.n37718 13.758
R36015 vdd.n37614 vdd.n37613 13.758
R36016 vdd.n28287 vdd.n28286 13.758
R36017 vdd.n28392 vdd.n28391 13.758
R36018 vdd.n28518 vdd.n28517 13.758
R36019 vdd.n28623 vdd.n28622 13.758
R36020 vdd.n28749 vdd.n28748 13.758
R36021 vdd.n28135 vdd.n28134 13.758
R36022 vdd.n28963 vdd.n28962 13.758
R36023 vdd.n27806 vdd.n27805 13.758
R36024 vdd.n29884 vdd.n29883 13.758
R36025 vdd.n31510 vdd.n31509 13.758
R36026 vdd.n32445 vdd.n32444 13.758
R36027 vdd.n30514 vdd.n30513 13.758
R36028 vdd.n2758 vdd.n2757 13.758
R36029 vdd.n2841 vdd.n2840 13.758
R36030 vdd.n2939 vdd.n2938 13.758
R36031 vdd.n3022 vdd.n3021 13.758
R36032 vdd.n3120 vdd.n3119 13.758
R36033 vdd.n3203 vdd.n3202 13.758
R36034 vdd.n3301 vdd.n3300 13.758
R36035 vdd.n3384 vdd.n3383 13.758
R36036 vdd.n3482 vdd.n3481 13.758
R36037 vdd.n3565 vdd.n3564 13.758
R36038 vdd.n2051 vdd.n2050 13.758
R36039 vdd.n2009 vdd.n2008 13.758
R36040 vdd.n2191 vdd.n2190 13.758
R36041 vdd.n2035 vdd.n2034 13.758
R36042 vdd.n2634 vdd.n2633 13.758
R36043 vdd.n1192 vdd.n1191 13.758
R36044 vdd.n1279 vdd.n1278 13.758
R36045 vdd.n1701 vdd.n1700 13.758
R36046 vdd.n1603 vdd.n1602 13.758
R36047 vdd.n1520 vdd.n1519 13.758
R36048 vdd.n1422 vdd.n1421 13.758
R36049 vdd.n1339 vdd.n1338 13.758
R36050 vdd.n26805 vdd.n26804 13.758
R36051 vdd.n26888 vdd.n26887 13.758
R36052 vdd.n26986 vdd.n26985 13.758
R36053 vdd.n27069 vdd.n27068 13.758
R36054 vdd.n27167 vdd.n27166 13.758
R36055 vdd.n27235 vdd.n27234 13.758
R36056 vdd.n31801 vdd.n31800 13.758
R36057 vdd.n31666 vdd.n31665 13.758
R36058 vdd.n32153 vdd.n32152 13.758
R36059 vdd.n31506 vdd.n31505 13.758
R36060 vdd.n32441 vdd.n32440 13.758
R36061 vdd.n31272 vdd.n31271 13.758
R36062 vdd.n13197 vdd.n9214 13.758
R36063 vdd.n13302 vdd.n9144 13.758
R36064 vdd.n13491 vdd.n8994 13.758
R36065 vdd.n13594 vdd.n8923 13.758
R36066 vdd.n13771 vdd.n8777 13.758
R36067 vdd.n13898 vdd.n8684 13.758
R36068 vdd.n14053 vdd.n8573 13.758
R36069 vdd.n14187 vdd.n8460 13.758
R36070 vdd.n14328 vdd.n8356 13.758
R36071 vdd.n8260 vdd.n8252 13.758
R36072 vdd.n8159 vdd.n8154 13.758
R36073 vdd.n14757 vdd.n8093 13.758
R36074 vdd.n14815 vdd.n14810 13.758
R36075 vdd.n14933 vdd.n8008 13.758
R36076 vdd.n13161 vdd.n9223 13.758
R36077 vdd.n13329 vdd.n9111 13.758
R36078 vdd.n13457 vdd.n9003 13.758
R36079 vdd.n13621 vdd.n8890 13.758
R36080 vdd.n13754 vdd.n8786 13.758
R36081 vdd.n13918 vdd.n8655 13.758
R36082 vdd.n14030 vdd.n8577 13.758
R36083 vdd.n14208 vdd.n8435 13.758
R36084 vdd.n14371 vdd.n8320 13.758
R36085 vdd.n14481 vdd.n8196 13.758
R36086 vdd.n19362 vdd.n19361 13.758
R36087 vdd.n19475 vdd.n19474 13.758
R36088 vdd.n19568 vdd.n19567 13.758
R36089 vdd.n19675 vdd.n19674 13.758
R36090 vdd.n19770 vdd.n19769 13.758
R36091 vdd.n20967 vdd.n20966 13.758
R36092 vdd.n20872 vdd.n20871 13.758
R36093 vdd.n20776 vdd.n20775 13.758
R36094 vdd.n20684 vdd.n20683 13.758
R36095 vdd.n20571 vdd.n20570 13.758
R36096 vdd.n21587 vdd.n21586 13.758
R36097 vdd.n21441 vdd.n21440 13.758
R36098 vdd.n21328 vdd.n21327 13.758
R36099 vdd.n21182 vdd.n21181 13.758
R36100 vdd.n21069 vdd.n21068 13.758
R36101 vdd.n19075 vdd.n19074 13.758
R36102 vdd.n18962 vdd.n18961 13.758
R36103 vdd.n18816 vdd.n18815 13.758
R36104 vdd.n18703 vdd.n18702 13.758
R36105 vdd.n18557 vdd.n18556 13.758
R36106 vdd.n20462 vdd.n20461 13.758
R36107 vdd.n20315 vdd.n20309 13.758
R36108 vdd.n20233 vdd.n20227 13.758
R36109 vdd.n20079 vdd.n20073 13.758
R36110 vdd.n24691 vdd.n24690 13.758
R36111 vdd.n25222 vdd.n25221 13.758
R36112 vdd.n10206 vdd.n10066 13.581
R36113 vdd.n13130 vdd.n9267 13.552
R36114 vdd.n9268 vdd.n9216 13.552
R36115 vdd.n13191 vdd.n13190 13.552
R36116 vdd.n13180 vdd.n13179 13.552
R36117 vdd.n13209 vdd.n9204 13.552
R36118 vdd.n13250 vdd.n13248 13.552
R36119 vdd.n13270 vdd.n13269 13.552
R36120 vdd.n13290 vdd.n13289 13.552
R36121 vdd.n13300 vdd.n13299 13.552
R36122 vdd.n13339 vdd.n13338 13.552
R36123 vdd.n13345 vdd.n13344 13.552
R36124 vdd.n13369 vdd.n13368 13.552
R36125 vdd.n13399 vdd.n9051 13.552
R36126 vdd.n13395 vdd.n9040 13.552
R36127 vdd.n13424 vdd.n9036 13.552
R36128 vdd.n9037 vdd.n8996 13.552
R36129 vdd.n13485 vdd.n13484 13.552
R36130 vdd.n13475 vdd.n13474 13.552
R36131 vdd.n13562 vdd.n13561 13.552
R36132 vdd.n13582 vdd.n13581 13.552
R36133 vdd.n13592 vdd.n13591 13.552
R36134 vdd.n13631 vdd.n13630 13.552
R36135 vdd.n13637 vdd.n13636 13.552
R36136 vdd.n13661 vdd.n13660 13.552
R36137 vdd.n13692 vdd.n8830 13.552
R36138 vdd.n13687 vdd.n8819 13.552
R36139 vdd.n13716 vdd.n8815 13.552
R36140 vdd.n8816 vdd.n8779 13.552
R36141 vdd.n13765 vdd.n13764 13.552
R36142 vdd.n13755 vdd.n8771 13.552
R36143 vdd.n13844 vdd.n13843 13.552
R36144 vdd.n13851 vdd.n13849 13.552
R36145 vdd.n13896 vdd.n13895 13.552
R36146 vdd.n8690 vdd.n8689 13.552
R36147 vdd.n13911 vdd.n8672 13.552
R36148 vdd.n8668 vdd.n8666 13.552
R36149 vdd.n13981 vdd.n13980 13.552
R36150 vdd.n13990 vdd.n8604 13.552
R36151 vdd.n8605 vdd.n8568 13.552
R36152 vdd.n14055 vdd.n14054 13.552
R36153 vdd.n14042 vdd.n14041 13.552
R36154 vdd.n14073 vdd.n14072 13.552
R36155 vdd.n14133 vdd.n14132 13.552
R36156 vdd.n14140 vdd.n14138 13.552
R36157 vdd.n14185 vdd.n14184 13.552
R36158 vdd.n8467 vdd.n8466 13.552
R36159 vdd.n14201 vdd.n8448 13.552
R36160 vdd.n8445 vdd.n8443 13.552
R36161 vdd.n14271 vdd.n14270 13.552
R36162 vdd.n14281 vdd.n8382 13.552
R36163 vdd.n8383 vdd.n8350 13.552
R36164 vdd.n14330 vdd.n14329 13.552
R36165 vdd.n14319 vdd.n8340 13.552
R36166 vdd.n14358 vdd.n8336 13.552
R36167 vdd.n8337 vdd.n8301 13.552
R36168 vdd.n14427 vdd.n14426 13.552
R36169 vdd.n8282 vdd.n8281 13.552
R36170 vdd.n14456 vdd.n8248 13.552
R36171 vdd.n8259 vdd.n8258 13.552
R36172 vdd.n14491 vdd.n14490 13.552
R36173 vdd.n14649 vdd.n14648 13.552
R36174 vdd.n8155 vdd.n8138 13.552
R36175 vdd.n14670 vdd.n14669 13.552
R36176 vdd.n14678 vdd.n8128 13.552
R36177 vdd.n14688 vdd.n14687 13.552
R36178 vdd.n14717 vdd.n14716 13.552
R36179 vdd.n14738 vdd.n14737 13.552
R36180 vdd.n14727 vdd.n14726 13.552
R36181 vdd.n14752 vdd.n14751 13.552
R36182 vdd.n14763 vdd.n14762 13.552
R36183 vdd.n14770 vdd.n14769 13.552
R36184 vdd.n14792 vdd.n14791 13.552
R36185 vdd.n14784 vdd.n14783 13.552
R36186 vdd.n14798 vdd.n14797 13.552
R36187 vdd.n14806 vdd.n8058 13.552
R36188 vdd.n14821 vdd.n14820 13.552
R36189 vdd.n14811 vdd.n8048 13.552
R36190 vdd.n14842 vdd.n14841 13.552
R36191 vdd.n14850 vdd.n8038 13.552
R36192 vdd.n14862 vdd.n14861 13.552
R36193 vdd.n14903 vdd.n14902 13.552
R36194 vdd.n14892 vdd.n14891 13.552
R36195 vdd.n14917 vdd.n14916 13.552
R36196 vdd.n14923 vdd.n14922 13.552
R36197 vdd.n14928 vdd.n8003 13.552
R36198 vdd.n13159 vdd.n13158 13.552
R36199 vdd.n13167 vdd.n9230 13.552
R36200 vdd.n13175 vdd.n13174 13.552
R36201 vdd.n13226 vdd.n13225 13.552
R36202 vdd.n9200 vdd.n9199 13.552
R36203 vdd.n13284 vdd.n13283 13.552
R36204 vdd.n13308 vdd.n9134 13.552
R36205 vdd.n13333 vdd.n9108 13.552
R36206 vdd.n9121 vdd.n9112 13.552
R36207 vdd.n13363 vdd.n9074 13.552
R36208 vdd.n9087 vdd.n9078 13.552
R36209 vdd.n9079 vdd.n9060 13.552
R36210 vdd.n13435 vdd.n13434 13.552
R36211 vdd.n9029 vdd.n9028 13.552
R36212 vdd.n13453 vdd.n13452 13.552
R36213 vdd.n13460 vdd.n13459 13.552
R36214 vdd.n13467 vdd.n13465 13.552
R36215 vdd.n13518 vdd.n13517 13.552
R36216 vdd.n8978 vdd.n8977 13.552
R36217 vdd.n13576 vdd.n13575 13.552
R36218 vdd.n13600 vdd.n8912 13.552
R36219 vdd.n13625 vdd.n8887 13.552
R36220 vdd.n8900 vdd.n8891 13.552
R36221 vdd.n13655 vdd.n8854 13.552
R36222 vdd.n8867 vdd.n8858 13.552
R36223 vdd.n8859 vdd.n8840 13.552
R36224 vdd.n13727 vdd.n13726 13.552
R36225 vdd.n8809 vdd.n8808 13.552
R36226 vdd.n13743 vdd.n13742 13.552
R36227 vdd.n13753 vdd.n13752 13.552
R36228 vdd.n13800 vdd.n13799 13.552
R36229 vdd.n8762 vdd.n8761 13.552
R36230 vdd.n8746 vdd.n8741 13.552
R36231 vdd.n13874 vdd.n13873 13.552
R36232 vdd.n13882 vdd.n13881 13.552
R36233 vdd.n8698 vdd.n8649 13.552
R36234 vdd.n13920 vdd.n13919 13.552
R36235 vdd.n13938 vdd.n13937 13.552
R36236 vdd.n13946 vdd.n13945 13.552
R36237 vdd.n13954 vdd.n13953 13.552
R36238 vdd.n13997 vdd.n13996 13.552
R36239 vdd.n14019 vdd.n14018 13.552
R36240 vdd.n14026 vdd.n14025 13.552
R36241 vdd.n14033 vdd.n14031 13.552
R36242 vdd.n14087 vdd.n14086 13.552
R36243 vdd.n8549 vdd.n8548 13.552
R36244 vdd.n8531 vdd.n8528 13.552
R36245 vdd.n14163 vdd.n14162 13.552
R36246 vdd.n14171 vdd.n14170 13.552
R36247 vdd.n8475 vdd.n8429 13.552
R36248 vdd.n14210 vdd.n14209 13.552
R36249 vdd.n14228 vdd.n14227 13.552
R36250 vdd.n14236 vdd.n14235 13.552
R36251 vdd.n14244 vdd.n14243 13.552
R36252 vdd.n14288 vdd.n14287 13.552
R36253 vdd.n14308 vdd.n14307 13.552
R36254 vdd.n14317 vdd.n14316 13.552
R36255 vdd.n14369 vdd.n14368 13.552
R36256 vdd.n8331 vdd.n8330 13.552
R36257 vdd.n14385 vdd.n14384 13.552
R36258 vdd.n14389 vdd.n14388 13.552
R36259 vdd.n14443 vdd.n14442 13.552
R36260 vdd.n14445 vdd.n8230 13.552
R36261 vdd.n14485 vdd.n8227 13.552
R36262 vdd.n14479 vdd.n14478 13.552
R36263 vdd.n14535 vdd.n8191 13.552
R36264 vdd.n14552 vdd.n14551 13.552
R36265 vdd.n14542 vdd.n14541 13.552
R36266 vdd.n11742 vdd.n11741 13.552
R36267 vdd.n11732 vdd.n11731 13.552
R36268 vdd.n11714 vdd.n11694 13.552
R36269 vdd.n11710 vdd.n11693 13.552
R36270 vdd.n11826 vdd.n11825 13.552
R36271 vdd.n11832 vdd.n11831 13.552
R36272 vdd.n11840 vdd.n11838 13.552
R36273 vdd.n11854 vdd.n11853 13.552
R36274 vdd.n23049 vdd.n23048 13.552
R36275 vdd.n21091 vdd.n21090 13.552
R36276 vdd.n19984 vdd.n19983 13.552
R36277 vdd.n21917 vdd.n21916 13.552
R36278 vdd.n21923 vdd.n21922 13.552
R36279 vdd.n21931 vdd.n21929 13.552
R36280 vdd.n21945 vdd.n21944 13.552
R36281 vdd.n13043 vdd.n9328 13.479
R36282 vdd.n13042 vdd.n9329 13.479
R36283 vdd.n12936 vdd.n12935 13.479
R36284 vdd.n9538 vdd.n9519 13.479
R36285 vdd.n12835 vdd.n9688 13.479
R36286 vdd.n12834 vdd.n9689 13.479
R36287 vdd.n12728 vdd.n12727 13.479
R36288 vdd.n9899 vdd.n9879 13.479
R36289 vdd.n12626 vdd.n10047 13.479
R36290 vdd.n15555 vdd.n15551 13.479
R36291 vdd.n15811 vdd.n15807 13.479
R36292 vdd.n16067 vdd.n16063 13.479
R36293 vdd.n16323 vdd.n16319 13.479
R36294 vdd.n16561 vdd.n16560 13.479
R36295 vdd.n27769 vdd.n27758 13.452
R36296 vdd.n33384 vdd.n33383 13.423
R36297 vdd.n34075 vdd.n34074 13.423
R36298 vdd.n33970 vdd.n33969 13.423
R36299 vdd.n34238 vdd.n34236 13.423
R36300 vdd.n35132 vdd.n35131 13.423
R36301 vdd.n35363 vdd.n35362 13.423
R36302 vdd.n35278 vdd.n35277 13.423
R36303 vdd.n34694 vdd.n34693 13.423
R36304 vdd.n34542 vdd.n34541 13.423
R36305 vdd.n34880 vdd.n34878 13.423
R36306 vdd.n699 vdd.n698 13.423
R36307 vdd.n498 vdd.n497 13.423
R36308 vdd.n6255 vdd.n6254 13.423
R36309 vdd.n6049 vdd.n6048 13.423
R36310 vdd.n5844 vdd.n5843 13.423
R36311 vdd.n5441 vdd.n5440 13.423
R36312 vdd.n5294 vdd.n5293 13.423
R36313 vdd.n5627 vdd.n5625 13.423
R36314 vdd.n4613 vdd.n4612 13.423
R36315 vdd.n5063 vdd.n5062 13.423
R36316 vdd.n4874 vdd.n4873 13.423
R36317 vdd.n4268 vdd.n4267 13.423
R36318 vdd.n4119 vdd.n4118 13.423
R36319 vdd.n4454 vdd.n4452 13.423
R36320 vdd.n27305 vdd.n27303 13.423
R36321 vdd.n27284 vdd.n27282 13.423
R36322 vdd.n27265 vdd.n27263 13.423
R36323 vdd.n25757 vdd.n25755 13.423
R36324 vdd.n25730 vdd.n25728 13.423
R36325 vdd.n25680 vdd.n25678 13.423
R36326 vdd.n25429 vdd.n25427 13.423
R36327 vdd.n21139 vdd.t351 13.37
R36328 vdd.n19015 vdd.t273 13.37
R36329 vdd.n3779 vdd.n3778 13.361
R36330 vdd.n2102 vdd.n2101 13.361
R36331 vdd.n1214 vdd.n1213 13.361
R36332 vdd.n3781 vdd.n3780 13.361
R36333 vdd.n2104 vdd.n2103 13.361
R36334 vdd.n1216 vdd.n1215 13.361
R36335 vdd.n33166 vdd.n33165 13.361
R36336 vdd.n37298 vdd.n37297 13.361
R36337 vdd.n37501 vdd.n37500 13.361
R36338 vdd.n33164 vdd.n33163 13.361
R36339 vdd.n37305 vdd.n37304 13.361
R36340 vdd.n37499 vdd.n37498 13.361
R36341 vdd.n31733 vdd.n31732 13.361
R36342 vdd.n31579 vdd.n31578 13.361
R36343 vdd.n32418 vdd.n32417 13.361
R36344 vdd.n31735 vdd.n31734 13.361
R36345 vdd.n31581 vdd.n31580 13.361
R36346 vdd.n32420 vdd.n32419 13.361
R36347 vdd.n28076 vdd.n28075 13.361
R36348 vdd.n27902 vdd.n27901 13.361
R36349 vdd.n30213 vdd.n30212 13.361
R36350 vdd.n28078 vdd.n28077 13.361
R36351 vdd.n27904 vdd.n27903 13.361
R36352 vdd.n30215 vdd.n30214 13.361
R36353 vdd.n33228 vdd.n33227 13.361
R36354 vdd.n37242 vdd.n37241 13.361
R36355 vdd.n32897 vdd.n32896 13.361
R36356 vdd.n13255 vdd.n9173 13.361
R36357 vdd.n13255 vdd.n13254 13.361
R36358 vdd.n13546 vdd.n8953 13.361
R36359 vdd.n13546 vdd.n13545 13.361
R36360 vdd.n13831 vdd.n8734 13.361
R36361 vdd.n13831 vdd.n13830 13.361
R36362 vdd.n8522 vdd.n8516 13.361
R36363 vdd.n8522 vdd.n8518 13.361
R36364 vdd.n14404 vdd.n8299 13.361
R36365 vdd.n14404 vdd.n14403 13.361
R36366 vdd.n13387 vdd.n9058 13.361
R36367 vdd.n13387 vdd.n13386 13.361
R36368 vdd.n13679 vdd.n8838 13.361
R36369 vdd.n13679 vdd.n13678 13.361
R36370 vdd.n14002 vdd.n8597 13.361
R36371 vdd.n14002 vdd.n14001 13.361
R36372 vdd.n14293 vdd.n8375 13.361
R36373 vdd.n14293 vdd.n14292 13.361
R36374 vdd.n8181 vdd.n8177 13.361
R36375 vdd.n8181 vdd.n8176 13.361
R36376 vdd.n19288 vdd.n19287 13.361
R36377 vdd.n19232 vdd.n19231 13.361
R36378 vdd.n19176 vdd.n19175 13.361
R36379 vdd.n19175 vdd.n19173 13.361
R36380 vdd.n19896 vdd.n19895 13.361
R36381 vdd.n19953 vdd.n19952 13.361
R36382 vdd.n18434 vdd.n18433 13.361
R36383 vdd.n18438 vdd.n18437 13.361
R36384 vdd.n18442 vdd.n18441 13.361
R36385 vdd.n18446 vdd.n18445 13.361
R36386 vdd.n18450 vdd.n18449 13.361
R36387 vdd.n12500 vdd.n10563 13.34
R36388 vdd.n10612 vdd.n10606 13.34
R36389 vdd.n10740 vdd.n10727 13.34
R36390 vdd.n10795 vdd.n10782 13.34
R36391 vdd.n10908 vdd.n10903 13.34
R36392 vdd.n10953 vdd.n10951 13.34
R36393 vdd.n12202 vdd.n11059 13.34
R36394 vdd.n12164 vdd.n11127 13.34
R36395 vdd.n11249 vdd.n11229 13.34
R36396 vdd.n11304 vdd.n11290 13.34
R36397 vdd.n11417 vdd.n11412 13.34
R36398 vdd.n11438 vdd.n11436 13.34
R36399 vdd.n10469 vdd.n10468 13.34
R36400 vdd.n10317 vdd.n10308 13.34
R36401 vdd.n13058 vdd.n9307 13.34
R36402 vdd.n9387 vdd.n9367 13.34
R36403 vdd.n9500 vdd.n9476 13.34
R36404 vdd.n12920 vdd.n9553 13.34
R36405 vdd.n12850 vdd.n9667 13.34
R36406 vdd.n9747 vdd.n9727 13.34
R36407 vdd.n9860 vdd.n9836 13.34
R36408 vdd.n12712 vdd.n9913 13.34
R36409 vdd.n12642 vdd.n10027 13.34
R36410 vdd.n10192 vdd.n10138 13.34
R36411 vdd.n16926 vdd.n16925 13.34
R36412 vdd.n17018 vdd.n17017 13.34
R36413 vdd.n17198 vdd.n17197 13.34
R36414 vdd.n17290 vdd.n17289 13.34
R36415 vdd.n17470 vdd.n17469 13.34
R36416 vdd.n17562 vdd.n17561 13.34
R36417 vdd.n17728 vdd.n17727 13.34
R36418 vdd.n17820 vdd.n17819 13.34
R36419 vdd.n17999 vdd.n17998 13.34
R36420 vdd.n18091 vdd.n18090 13.34
R36421 vdd.n18268 vdd.n18267 13.34
R36422 vdd.n18340 vdd.n18339 13.34
R36423 vdd.n15274 vdd.n15270 13.34
R36424 vdd.n15354 vdd.n15349 13.34
R36425 vdd.n15496 vdd.n15489 13.34
R36426 vdd.n15593 vdd.n15586 13.34
R36427 vdd.n15752 vdd.n15745 13.34
R36428 vdd.n15849 vdd.n15842 13.34
R36429 vdd.n16008 vdd.n16001 13.34
R36430 vdd.n16105 vdd.n16098 13.34
R36431 vdd.n16264 vdd.n16257 13.34
R36432 vdd.n16361 vdd.n16354 13.34
R36433 vdd.n16520 vdd.n16513 13.34
R36434 vdd.n16727 vdd.n16725 13.34
R36435 vdd.n203 vdd.n202 13.176
R36436 vdd.n35921 vdd.n35920 13.176
R36437 vdd.n36152 vdd.n36151 13.176
R36438 vdd.n36383 vdd.n36382 13.176
R36439 vdd.n36614 vdd.n36613 13.176
R36440 vdd.n36845 vdd.n36844 13.176
R36441 vdd.n37900 vdd.n37899 13.176
R36442 vdd.n37669 vdd.n37668 13.176
R36443 vdd.n28342 vdd.n28341 13.176
R36444 vdd.n28573 vdd.n28572 13.176
R36445 vdd.n1563 vdd.n1562 13.176
R36446 vdd.n1382 vdd.n1381 13.176
R36447 vdd.n26848 vdd.n26847 13.176
R36448 vdd.n27029 vdd.n27028 13.176
R36449 vdd.n2801 vdd.n2800 13.176
R36450 vdd.n2982 vdd.n2981 13.176
R36451 vdd.n3163 vdd.n3162 13.176
R36452 vdd.n3344 vdd.n3343 13.176
R36453 vdd.n3525 vdd.n3524 13.176
R36454 vdd.n12987 vdd.n12986 13.158
R36455 vdd.n12880 vdd.n12879 13.158
R36456 vdd.n12779 vdd.n12778 13.158
R36457 vdd.n12672 vdd.n12671 13.158
R36458 vdd.n10485 vdd.n10484 13.158
R36459 vdd.n33574 vdd.n33573 12.92
R36460 vdd.n1050 vdd.n1049 12.92
R36461 vdd.n29684 vdd.n29682 12.92
R36462 vdd.n13031 vdd.n13030 12.837
R36463 vdd.n12823 vdd.n12822 12.837
R36464 vdd.n12721 vdd.n9885 12.837
R36465 vdd.n12614 vdd.n12613 12.837
R36466 vdd.n11599 vdd.t370 12.837
R36467 vdd.n16555 vdd.n16554 12.837
R36468 vdd.n15016 vdd.t27 12.837
R36469 vdd.n25245 vdd.n25244 12.807
R36470 vdd.n25244 vdd.n25243 12.807
R36471 vdd.n14706 vdd.n14704 12.8
R36472 vdd.n14706 vdd.n14705 12.8
R36473 vdd.n14879 vdd.n8028 12.8
R36474 vdd.n14879 vdd.n14878 12.8
R36475 vdd.n11714 vdd.n11713 12.8
R36476 vdd.n11713 vdd.n11693 12.8
R36477 vdd.n11855 vdd.n11840 12.8
R36478 vdd.n11855 vdd.n11854 12.8
R36479 vdd.n24089 vdd.n24085 12.8
R36480 vdd.n24089 vdd.n24088 12.8
R36481 vdd.n23857 vdd.n23853 12.8
R36482 vdd.n23857 vdd.n23856 12.8
R36483 vdd.n23169 vdd.n23165 12.8
R36484 vdd.n23169 vdd.n23168 12.8
R36485 vdd.n23401 vdd.n23397 12.8
R36486 vdd.n23401 vdd.n23400 12.8
R36487 vdd.n22590 vdd.n22586 12.8
R36488 vdd.n22590 vdd.n22589 12.8
R36489 vdd.n22822 vdd.n22818 12.8
R36490 vdd.n22822 vdd.n22821 12.8
R36491 vdd.n22373 vdd.n22369 12.8
R36492 vdd.n22373 vdd.n22372 12.8
R36493 vdd.n24318 vdd.n24314 12.8
R36494 vdd.n24318 vdd.n24317 12.8
R36495 vdd.n20390 vdd.n20387 12.8
R36496 vdd.n20390 vdd.n20389 12.8
R36497 vdd.n20154 vdd.n20151 12.8
R36498 vdd.n20154 vdd.n20153 12.8
R36499 vdd.n21788 vdd.n21786 12.8
R36500 vdd.n21788 vdd.n21787 12.8
R36501 vdd.n21946 vdd.n21931 12.8
R36502 vdd.n21946 vdd.n21945 12.8
R36503 vdd.n24748 vdd.n24746 12.8
R36504 vdd.n24748 vdd.n24747 12.8
R36505 vdd.n25164 vdd.n25162 12.8
R36506 vdd.n25164 vdd.n25163 12.8
R36507 vdd.n9454 vdd.n9421 12.516
R36508 vdd.n9647 vdd.n9646 12.516
R36509 vdd.n9814 vdd.n9813 12.516
R36510 vdd.n10007 vdd.n10006 12.516
R36511 vdd.n10494 vdd.n10480 12.516
R36512 vdd.n12354 vdd.t310 12.516
R36513 vdd.n15083 vdd.n15079 12.516
R36514 vdd.n14603 vdd.n14602 12.234
R36515 vdd.n24803 vdd.n24802 12.234
R36516 vdd.n25108 vdd.n25107 12.234
R36517 vdd.n9384 vdd.n9383 12.195
R36518 vdd.n9555 vdd.n9554 12.195
R36519 vdd.n9744 vdd.n9743 12.195
R36520 vdd.n9915 vdd.n9914 12.195
R36521 vdd.n10189 vdd.n10188 12.195
R36522 vdd.n12343 vdd.t379 12.195
R36523 vdd.n10551 vdd.n10536 12.127
R36524 vdd.n10648 vdd.n10631 12.127
R36525 vdd.n10712 vdd.n10700 12.127
R36526 vdd.n12351 vdd.n10806 12.127
R36527 vdd.n12316 vdd.n10868 12.127
R36528 vdd.n12262 vdd.n10962 12.127
R36529 vdd.n12211 vdd.n11044 12.127
R36530 vdd.n11155 vdd.n11139 12.127
R36531 vdd.n12106 vdd.n11220 12.127
R36532 vdd.n12045 vdd.n11315 12.127
R36533 vdd.n12010 vdd.n11377 12.127
R36534 vdd.n11956 vdd.n11447 12.127
R36535 vdd.n10406 vdd.n10325 12.127
R36536 vdd.n13079 vdd.n9292 12.127
R36537 vdd.n13011 vdd.n9398 12.127
R36538 vdd.n9462 vdd.n9456 12.127
R36539 vdd.n9592 vdd.n9580 12.127
R36540 vdd.n12871 vdd.n9624 12.127
R36541 vdd.n12803 vdd.n9758 12.127
R36542 vdd.n9822 vdd.n9816 12.127
R36543 vdd.n9952 vdd.n9940 12.127
R36544 vdd.n12663 vdd.n9984 12.127
R36545 vdd.n10110 vdd.n10109 12.127
R36546 vdd.n16900 vdd.n16894 12.127
R36547 vdd.n17056 vdd.n17050 12.127
R36548 vdd.n17172 vdd.n17166 12.127
R36549 vdd.n17328 vdd.n17322 12.127
R36550 vdd.n17444 vdd.n17438 12.127
R36551 vdd.n17595 vdd.n16829 12.127
R36552 vdd.n17702 vdd.n17696 12.127
R36553 vdd.n17858 vdd.n17852 12.127
R36554 vdd.n17973 vdd.n17967 12.127
R36555 vdd.n18129 vdd.n18123 12.127
R36556 vdd.n18243 vdd.n18238 12.127
R36557 vdd.n15024 vdd.n15020 12.127
R36558 vdd.n15378 vdd.n15377 12.127
R36559 vdd.n15452 vdd.n15451 12.127
R36560 vdd.n15620 vdd.n15619 12.127
R36561 vdd.n15708 vdd.n15707 12.127
R36562 vdd.n15876 vdd.n15875 12.127
R36563 vdd.n15964 vdd.n15963 12.127
R36564 vdd.n16132 vdd.n16131 12.127
R36565 vdd.n16220 vdd.n16219 12.127
R36566 vdd.n16388 vdd.n16387 12.127
R36567 vdd.n16476 vdd.n16475 12.127
R36568 vdd.n16622 vdd.n16621 12.127
R36569 vdd.n31689 vdd.n31688 12.047
R36570 vdd.n13081 vdd.n9289 11.875
R36571 vdd.n12972 vdd.n9455 11.875
R36572 vdd.n12873 vdd.n9621 11.875
R36573 vdd.n12764 vdd.n9815 11.875
R36574 vdd.n12665 vdd.n9981 11.875
R36575 vdd.n12567 vdd.n12566 11.875
R36576 vdd.n15116 vdd.n15115 11.875
R36577 vdd.n35845 vdd.n35710 11.793
R36578 vdd.n36003 vdd.n35999 11.793
R36579 vdd.n36073 vdd.n36069 11.793
R36580 vdd.n36234 vdd.n36230 11.793
R36581 vdd.n36304 vdd.n36300 11.793
R36582 vdd.n36465 vdd.n36461 11.793
R36583 vdd.n36535 vdd.n36531 11.793
R36584 vdd.n36696 vdd.n36692 11.793
R36585 vdd.n36766 vdd.n36762 11.793
R36586 vdd.n36927 vdd.n36923 11.793
R36587 vdd.n37005 vdd.n37004 11.793
R36588 vdd.n33174 vdd.n33170 11.793
R36589 vdd.n33136 vdd.n33132 11.793
R36590 vdd.n37312 vdd.n37311 11.793
R36591 vdd.n37387 vdd.n37383 11.793
R36592 vdd.n32848 vdd.n32844 11.793
R36593 vdd.n38212 vdd.n38208 11.793
R36594 vdd.n38052 vdd.n38048 11.793
R36595 vdd.n37982 vdd.n37978 11.793
R36596 vdd.n37821 vdd.n37817 11.793
R36597 vdd.n37751 vdd.n37747 11.793
R36598 vdd.n28193 vdd.n28189 11.793
R36599 vdd.n28263 vdd.n28259 11.793
R36600 vdd.n28424 vdd.n28420 11.793
R36601 vdd.n28494 vdd.n28490 11.793
R36602 vdd.n28655 vdd.n28651 11.793
R36603 vdd.n28725 vdd.n28721 11.793
R36604 vdd.n26209 vdd.n26208 11.793
R36605 vdd.n31754 vdd.n31753 11.793
R36606 vdd.n27838 vdd.n27834 11.793
R36607 vdd.n27914 vdd.n27910 11.793
R36608 vdd.n31487 vdd.n31486 11.793
R36609 vdd.n30221 vdd.n30217 11.793
R36610 vdd.n30504 vdd.n30346 11.793
R36611 vdd.n2740 vdd.n2739 11.793
R36612 vdd.n2864 vdd.n2863 11.793
R36613 vdd.n2918 vdd.n2917 11.793
R36614 vdd.n3045 vdd.n3044 11.793
R36615 vdd.n3099 vdd.n3098 11.793
R36616 vdd.n3226 vdd.n3225 11.793
R36617 vdd.n3280 vdd.n3279 11.793
R36618 vdd.n3407 vdd.n3406 11.793
R36619 vdd.n3461 vdd.n3460 11.793
R36620 vdd.n3588 vdd.n3587 11.793
R36621 vdd.n3654 vdd.n3650 11.793
R36622 vdd.n3936 vdd.n3935 11.793
R36623 vdd.n2217 vdd.n2216 11.793
R36624 vdd.n2403 vdd.n2399 11.793
R36625 vdd.n2600 vdd.n2599 11.793
R36626 vdd.n1224 vdd.n1223 11.793
R36627 vdd.n1781 vdd.n1780 11.793
R36628 vdd.n1680 vdd.n1679 11.793
R36629 vdd.n1626 vdd.n1625 11.793
R36630 vdd.n1499 vdd.n1498 11.793
R36631 vdd.n1445 vdd.n1444 11.793
R36632 vdd.n1318 vdd.n1317 11.793
R36633 vdd.n26784 vdd.n26783 11.793
R36634 vdd.n26911 vdd.n26910 11.793
R36635 vdd.n26965 vdd.n26964 11.793
R36636 vdd.n27092 vdd.n27091 11.793
R36637 vdd.n27146 vdd.n27145 11.793
R36638 vdd.n26211 vdd.n26204 11.793
R36639 vdd.n31756 vdd.n31749 11.793
R36640 vdd.n31641 vdd.n31640 11.793
R36641 vdd.n32097 vdd.n32096 11.793
R36642 vdd.n31489 vdd.n31482 11.793
R36643 vdd.n32484 vdd.n32483 11.793
R36644 vdd.n31146 vdd.n31145 11.793
R36645 vdd.n13119 vdd.n9265 11.793
R36646 vdd.n13347 vdd.n9095 11.793
R36647 vdd.n13411 vdd.n9034 11.793
R36648 vdd.n13639 vdd.n8875 11.793
R36649 vdd.n13705 vdd.n8813 11.793
R36650 vdd.n13907 vdd.n13906 11.793
R36651 vdd.n13987 vdd.n8603 11.793
R36652 vdd.n14197 vdd.n14196 11.793
R36653 vdd.n14278 vdd.n8381 11.793
R36654 vdd.n14499 vdd.n8217 11.793
R36655 vdd.n14671 vdd.n8133 11.793
R36656 vdd.n14728 vdd.n14723 11.793
R36657 vdd.n14843 vdd.n8043 11.793
R36658 vdd.n14915 vdd.n8015 11.793
R36659 vdd.n13228 vdd.n9192 11.793
R36660 vdd.n13315 vdd.n9106 11.793
R36661 vdd.n13520 vdd.n8970 11.793
R36662 vdd.n13607 vdd.n8885 11.793
R36663 vdd.n13794 vdd.n8764 11.793
R36664 vdd.n13887 vdd.n8696 11.793
R36665 vdd.n14081 vdd.n8551 11.793
R36666 vdd.n14176 vdd.n8473 11.793
R36667 vdd.n14382 vdd.n8311 11.793
R36668 vdd.n14469 vdd.n8225 11.793
R36669 vdd.n19336 vdd.n19303 11.793
R36670 vdd.n19512 vdd.n19506 11.793
R36671 vdd.n19542 vdd.n19536 11.793
R36672 vdd.n19713 vdd.n19707 11.793
R36673 vdd.n19744 vdd.n19738 11.793
R36674 vdd.n20941 vdd.n20935 11.793
R36675 vdd.n20910 vdd.n20904 11.793
R36676 vdd.n20751 vdd.n20745 11.793
R36677 vdd.n20721 vdd.n20715 11.793
R36678 vdd.n20545 vdd.n19973 11.793
R36679 vdd.n21561 vdd.n21555 11.793
R36680 vdd.n21479 vdd.n21473 11.793
R36681 vdd.n21302 vdd.n21296 11.793
R36682 vdd.n21220 vdd.n21214 11.793
R36683 vdd.n21043 vdd.n21037 11.793
R36684 vdd.n19113 vdd.n19107 11.793
R36685 vdd.n18936 vdd.n18930 11.793
R36686 vdd.n18854 vdd.n18848 11.793
R36687 vdd.n18677 vdd.n18671 11.793
R36688 vdd.n18595 vdd.n18589 11.793
R36689 vdd.n20431 vdd.n20430 11.793
R36690 vdd.n20341 vdd.n20340 11.793
R36691 vdd.n20195 vdd.n20194 11.793
R36692 vdd.n20105 vdd.n20104 11.793
R36693 vdd.n24778 vdd.n24777 11.793
R36694 vdd.n25131 vdd.n25130 11.793
R36695 vdd.n21000 vdd.n20999 11.728
R36696 vdd.n315 vdd.n313 11.67
R36697 vdd.n2003 vdd.n2002 11.67
R36698 vdd.n11617 vdd.n11582 11.67
R36699 vdd.n35932 vdd.n35929 11.623
R36700 vdd.n36163 vdd.n36160 11.623
R36701 vdd.n36394 vdd.n36391 11.623
R36702 vdd.n36625 vdd.n36622 11.623
R36703 vdd.n36856 vdd.n36853 11.623
R36704 vdd.n33248 vdd.n33245 11.623
R36705 vdd.n37258 vdd.n37255 11.623
R36706 vdd.n37444 vdd.n37443 11.623
R36707 vdd.n38134 vdd.n38131 11.623
R36708 vdd.n37911 vdd.n37910 11.623
R36709 vdd.n37680 vdd.n37679 11.623
R36710 vdd.n28353 vdd.n28350 11.623
R36711 vdd.n28584 vdd.n28581 11.623
R36712 vdd.n28151 vdd.n28148 11.623
R36713 vdd.n27766 vdd.n27765 11.623
R36714 vdd.n29692 vdd.n29689 11.623
R36715 vdd.n30298 vdd.n30297 11.623
R36716 vdd.n13265 vdd.n9157 11.622
R36717 vdd.n13287 vdd.n13286 11.622
R36718 vdd.n9142 vdd.n9130 11.622
R36719 vdd.n13328 vdd.n9094 11.622
R36720 vdd.n13355 vdd.n13354 11.622
R36721 vdd.n13557 vdd.n13556 11.622
R36722 vdd.n13579 vdd.n13578 11.622
R36723 vdd.n8921 vdd.n8920 11.622
R36724 vdd.n13628 vdd.n13627 11.622
R36725 vdd.n13658 vdd.n13657 11.622
R36726 vdd.n13839 vdd.n8718 11.622
R36727 vdd.n13871 vdd.n8707 11.622
R36728 vdd.n13879 vdd.n8682 11.622
R36729 vdd.n8694 vdd.t110 11.622
R36730 vdd.n13917 vdd.n8656 11.622
R36731 vdd.n13943 vdd.n8621 11.622
R36732 vdd.n8498 vdd.n8496 11.622
R36733 vdd.n14160 vdd.n8484 11.622
R36734 vdd.n14168 vdd.n8458 11.622
R36735 vdd.n8471 vdd.n8425 11.622
R36736 vdd.n14225 vdd.n8420 11.622
R36737 vdd.n8286 vdd.n8239 11.622
R36738 vdd.n14440 vdd.n14438 11.622
R36739 vdd.n8261 vdd.n8232 11.622
R36740 vdd.n14480 vdd.n8216 11.622
R36741 vdd.n33476 vdd.n33475 11.609
R36742 vdd.n33384 vdd.n33382 11.609
R36743 vdd.n33386 vdd.n33385 11.609
R36744 vdd.n34075 vdd.n34073 11.609
R36745 vdd.n34235 vdd.n34234 11.609
R36746 vdd.n33970 vdd.n33968 11.609
R36747 vdd.n33967 vdd.n33966 11.609
R36748 vdd.n34238 vdd.n34237 11.609
R36749 vdd.n35134 vdd.n35133 11.609
R36750 vdd.n35132 vdd.n35130 11.609
R36751 vdd.n35360 vdd.n35359 11.609
R36752 vdd.n35363 vdd.n35361 11.609
R36753 vdd.n35278 vdd.n35276 11.609
R36754 vdd.n34694 vdd.n34692 11.609
R36755 vdd.n34877 vdd.n34876 11.609
R36756 vdd.n34547 vdd.n34546 11.609
R36757 vdd.n34542 vdd.n34540 11.609
R36758 vdd.n34880 vdd.n34879 11.609
R36759 vdd.n1048 vdd.n1047 11.609
R36760 vdd.n696 vdd.n695 11.609
R36761 vdd.n699 vdd.n697 11.609
R36762 vdd.n88 vdd.n87 11.609
R36763 vdd.n495 vdd.n494 11.609
R36764 vdd.n498 vdd.n496 11.609
R36765 vdd.n6255 vdd.n6253 11.609
R36766 vdd.n6252 vdd.n6251 11.609
R36767 vdd.n6049 vdd.n6047 11.609
R36768 vdd.n6051 vdd.n6050 11.609
R36769 vdd.n5844 vdd.n5842 11.609
R36770 vdd.n5441 vdd.n5439 11.609
R36771 vdd.n5624 vdd.n5623 11.609
R36772 vdd.n5294 vdd.n5292 11.609
R36773 vdd.n5288 vdd.n5287 11.609
R36774 vdd.n5627 vdd.n5626 11.609
R36775 vdd.n4610 vdd.n4609 11.609
R36776 vdd.n4613 vdd.n4611 11.609
R36777 vdd.n5065 vdd.n5064 11.609
R36778 vdd.n5063 vdd.n5061 11.609
R36779 vdd.n4874 vdd.n4872 11.609
R36780 vdd.n4268 vdd.n4266 11.609
R36781 vdd.n4451 vdd.n4450 11.609
R36782 vdd.n4124 vdd.n4123 11.609
R36783 vdd.n4119 vdd.n4117 11.609
R36784 vdd.n4454 vdd.n4453 11.609
R36785 vdd.n27305 vdd.n27304 11.609
R36786 vdd.n27281 vdd.n27280 11.609
R36787 vdd.n27284 vdd.n27283 11.609
R36788 vdd.n27262 vdd.n27261 11.609
R36789 vdd.n27265 vdd.n27264 11.609
R36790 vdd.n25757 vdd.n25756 11.609
R36791 vdd.n25727 vdd.n25726 11.609
R36792 vdd.n25730 vdd.n25729 11.609
R36793 vdd.n25680 vdd.n25679 11.609
R36794 vdd.n25682 vdd.n25681 11.609
R36795 vdd.n25429 vdd.n25428 11.609
R36796 vdd.n24528 vdd.n24527 11.572
R36797 vdd.n10381 vdd.n10339 11.554
R36798 vdd.n13024 vdd.n9359 11.554
R36799 vdd.n12917 vdd.n9556 11.554
R36800 vdd.n12816 vdd.n9719 11.554
R36801 vdd.n12607 vdd.n10061 11.554
R36802 vdd.n10597 vdd.n10583 11.554
R36803 vdd.n10762 vdd.n10757 11.554
R36804 vdd.n12285 vdd.n10917 11.554
R36805 vdd.n11117 vdd.n11096 11.554
R36806 vdd.n12073 vdd.n12072 11.554
R36807 vdd.n11979 vdd.n11426 11.554
R36808 vdd.t374 vdd.n11437 11.554
R36809 vdd.n16614 vdd.n16612 11.554
R36810 vdd.n13110 vdd.n9277 11.515
R36811 vdd.n13153 vdd.n9239 11.515
R36812 vdd.n13186 vdd.n9224 11.515
R36813 vdd.n13205 vdd.n9190 11.515
R36814 vdd.n13219 vdd.n13217 11.515
R36815 vdd.n11661 vdd.n11566 11.515
R36816 vdd.n15006 vdd.n15005 11.515
R36817 vdd.n34206 vdd.n34202 11.482
R36818 vdd.n35290 vdd.n35286 11.482
R36819 vdd.n34706 vdd.n34702 11.482
R36820 vdd.n5907 vdd.n5903 11.482
R36821 vdd.n5453 vdd.n5449 11.482
R36822 vdd.n4280 vdd.n4276 11.482
R36823 vdd.n27342 vdd.n27338 11.482
R36824 vdd.n25794 vdd.n25790 11.482
R36825 vdd.n11782 vdd.n11780 11.455
R36826 vdd.n24100 vdd.n24099 11.309
R36827 vdd.n24074 vdd.n24073 11.309
R36828 vdd.n23868 vdd.n23867 11.309
R36829 vdd.n23842 vdd.n23841 11.309
R36830 vdd.n23636 vdd.n23635 11.309
R36831 vdd.n23154 vdd.n23153 11.309
R36832 vdd.n23180 vdd.n23179 11.309
R36833 vdd.n23386 vdd.n23385 11.309
R36834 vdd.n23412 vdd.n23411 11.309
R36835 vdd.n23618 vdd.n23617 11.309
R36836 vdd.n22575 vdd.n22574 11.309
R36837 vdd.n22601 vdd.n22600 11.309
R36838 vdd.n22807 vdd.n22806 11.309
R36839 vdd.n22833 vdd.n22832 11.309
R36840 vdd.n23039 vdd.n23038 11.309
R36841 vdd.n22191 vdd.n22190 11.309
R36842 vdd.n22356 vdd.n22355 11.309
R36843 vdd.n22049 vdd.n22048 11.309
R36844 vdd.n22085 vdd.n22084 11.309
R36845 vdd.n22170 vdd.n22169 11.309
R36846 vdd.n33786 vdd.n33784 11.294
R36847 vdd.n862 vdd.n860 11.294
R36848 vdd.n30574 vdd.n30573 11.294
R36849 vdd.n29020 vdd.n29019 11.294
R36850 vdd.n29852 vdd.n29851 11.294
R36851 vdd.n13142 vdd.n13141 11.294
R36852 vdd.n21664 vdd.n21660 11.259
R36853 vdd.n21673 vdd.n21672 11.259
R36854 vdd.n21398 vdd.n21394 11.259
R36855 vdd.n21381 vdd.n21380 11.259
R36856 vdd.n21139 vdd.n21135 11.259
R36857 vdd.n21122 vdd.n21121 11.259
R36858 vdd.n19060 vdd.t348 11.259
R36859 vdd.n19032 vdd.n19028 11.259
R36860 vdd.n19015 vdd.n19014 11.259
R36861 vdd.n18773 vdd.n18769 11.259
R36862 vdd.n18756 vdd.n18755 11.259
R36863 vdd.n18514 vdd.n18510 11.259
R36864 vdd.n18497 vdd.n18496 11.259
R36865 vdd.n10266 vdd.n10265 11.249
R36866 vdd.n12963 vdd.n12962 11.233
R36867 vdd.n12866 vdd.n12865 11.233
R36868 vdd.n12755 vdd.n12754 11.233
R36869 vdd.n12658 vdd.n12657 11.233
R36870 vdd.n12222 vdd.t309 11.233
R36871 vdd.n15717 vdd.n15716 11.233
R36872 vdd.n15973 vdd.n15972 11.233
R36873 vdd.n16229 vdd.n16228 11.233
R36874 vdd.n16485 vdd.n16484 11.233
R36875 vdd.n13162 vdd.t324 11.195
R36876 vdd.n11626 vdd.n11625 11.18
R36877 vdd.n21636 vdd.n21632 11.18
R36878 vdd.n19243 vdd.t170 11.141
R36879 vdd.n19909 vdd.t166 11.141
R36880 vdd.n218 vdd.n216 11.112
R36881 vdd.n364 vdd.n360 11.106
R36882 vdd.n24678 vdd.n24677 11.087
R36883 vdd.n25233 vdd.n25232 11.087
R36884 vdd.n25232 vdd.n25231 11.087
R36885 vdd.n24677 vdd.n24676 11.087
R36886 vdd.n13428 vdd.n9032 11.01
R36887 vdd.n13455 vdd.n8993 11.01
R36888 vdd.n13480 vdd.n13472 11.01
R36889 vdd.n13499 vdd.n8969 11.01
R36890 vdd.n13511 vdd.n13510 11.01
R36891 vdd.n13683 vdd.n8800 11.01
R36892 vdd.n13737 vdd.n8796 11.01
R36893 vdd.n13746 vdd.n13745 11.01
R36894 vdd.n13760 vdd.n8753 11.01
R36895 vdd.n13793 vdd.n8765 11.01
R36896 vdd.n13810 vdd.n8749 11.01
R36897 vdd.n14012 vdd.n8588 11.01
R36898 vdd.n14050 vdd.n14038 11.01
R36899 vdd.n14069 vdd.n8540 11.01
R36900 vdd.n14080 vdd.n14078 11.01
R36901 vdd.n14097 vdd.n8535 11.01
R36902 vdd.n8379 vdd.n8377 11.01
R36903 vdd.n14310 vdd.n8347 11.01
R36904 vdd.n14362 vdd.n8327 11.01
R36905 vdd.n14354 vdd.n8312 11.01
R36906 vdd.n14395 vdd.n14394 11.01
R36907 vdd.n14488 vdd.t321 11.01
R36908 vdd.n25048 vdd.n24990 10.99
R36909 vdd.n31923 vdd.n31917 10.917
R36910 vdd.n30552 vdd.n30551 10.917
R36911 vdd.n12512 vdd.n10531 10.914
R36912 vdd.n10616 vdd.n10613 10.914
R36913 vdd.n10728 vdd.n10707 10.914
R36914 vdd.n12363 vdd.n10775 10.914
R36915 vdd.n12304 vdd.n10895 10.914
R36916 vdd.n10982 vdd.n10968 10.914
R36917 vdd.n11077 vdd.n11064 10.914
R36918 vdd.n11135 vdd.n11129 10.914
R36919 vdd.n11233 vdd.n11228 10.914
R36920 vdd.n12057 vdd.n11283 10.914
R36921 vdd.n11998 vdd.n11404 10.914
R36922 vdd.n11529 vdd.n11524 10.914
R36923 vdd.n10475 vdd.n10474 10.914
R36924 vdd.n10418 vdd.n10315 10.914
R36925 vdd.n13070 vdd.n9299 10.914
R36926 vdd.n13022 vdd.n9362 10.914
R36927 vdd.n9495 vdd.n9484 10.914
R36928 vdd.n12908 vdd.n9557 10.914
R36929 vdd.n12862 vdd.n9659 10.914
R36930 vdd.n12814 vdd.n9722 10.914
R36931 vdd.n9855 vdd.n9844 10.914
R36932 vdd.n12700 vdd.n9916 10.914
R36933 vdd.n12654 vdd.n10019 10.914
R36934 vdd.n12605 vdd.n12604 10.914
R36935 vdd.n16910 vdd.n16909 10.914
R36936 vdd.n17034 vdd.n17033 10.914
R36937 vdd.n17182 vdd.n17181 10.914
R36938 vdd.n17306 vdd.n17305 10.914
R36939 vdd.n17454 vdd.n17453 10.914
R36940 vdd.n17578 vdd.n17577 10.914
R36941 vdd.n17712 vdd.n17711 10.914
R36942 vdd.n17836 vdd.n17835 10.914
R36943 vdd.n17983 vdd.n17982 10.914
R36944 vdd.n18107 vdd.n18106 10.914
R36945 vdd.n18253 vdd.n18252 10.914
R36946 vdd.n18362 vdd.n18361 10.914
R36947 vdd.n15263 vdd.n15259 10.914
R36948 vdd.n15368 vdd.n15364 10.914
R36949 vdd.n15479 vdd.n15472 10.914
R36950 vdd.n15610 vdd.n15603 10.914
R36951 vdd.n15735 vdd.n15728 10.914
R36952 vdd.n15866 vdd.n15859 10.914
R36953 vdd.n15991 vdd.n15984 10.914
R36954 vdd.n16122 vdd.n16115 10.914
R36955 vdd.n16247 vdd.n16240 10.914
R36956 vdd.n16378 vdd.n16371 10.914
R36957 vdd.n16503 vdd.n16496 10.914
R36958 vdd.n9400 vdd.n9399 10.912
R36959 vdd.n12906 vdd.n12905 10.912
R36960 vdd.n9760 vdd.n9759 10.912
R36961 vdd.n12698 vdd.n12697 10.912
R36962 vdd.n10106 vdd.n10105 10.912
R36963 vdd.n10598 vdd.t368 10.912
R36964 vdd.n16620 vdd.n16618 10.912
R36965 vdd.n16976 vdd.t20 10.912
R36966 vdd.n33777 vdd.n33775 10.736
R36967 vdd.n872 vdd.n870 10.736
R36968 vdd.n33837 vdd.n33836 10.729
R36969 vdd.n798 vdd.n797 10.729
R36970 vdd.n24627 vdd.n24626 10.623
R36971 vdd.n9308 vdd.n9298 10.591
R36972 vdd.n9497 vdd.n9496 10.591
R36973 vdd.n9668 vdd.n9658 10.591
R36974 vdd.n9857 vdd.n9856 10.591
R36975 vdd.n10028 vdd.n10018 10.591
R36976 vdd.n15478 vdd.n15477 10.591
R36977 vdd.n15734 vdd.n15733 10.591
R36978 vdd.n15990 vdd.n15989 10.591
R36979 vdd.n16246 vdd.n16245 10.591
R36980 vdd.n16502 vdd.n16501 10.591
R36981 vdd.n24186 vdd.n24182 10.588
R36982 vdd.n23992 vdd.n23988 10.588
R36983 vdd.n23954 vdd.n23950 10.588
R36984 vdd.n23760 vdd.n23756 10.588
R36985 vdd.n23722 vdd.n23718 10.588
R36986 vdd.n23072 vdd.n23068 10.588
R36987 vdd.n23266 vdd.n23262 10.588
R36988 vdd.n23304 vdd.n23300 10.588
R36989 vdd.n23498 vdd.n23494 10.588
R36990 vdd.n23536 vdd.n23532 10.588
R36991 vdd.n22493 vdd.n22489 10.588
R36992 vdd.n22687 vdd.n22683 10.588
R36993 vdd.n22725 vdd.n22721 10.588
R36994 vdd.n22919 vdd.n22915 10.588
R36995 vdd.n22957 vdd.n22953 10.588
R36996 vdd.n22463 vdd.n22459 10.588
R36997 vdd.n22335 vdd.n22334 10.588
R36998 vdd.n22319 vdd.n22315 10.588
R36999 vdd.n22137 vdd.n22136 10.588
R37000 vdd.n24291 vdd.n24287 10.588
R37001 vdd.n21527 vdd.n21524 10.555
R37002 vdd.n21509 vdd.n21506 10.555
R37003 vdd.n21268 vdd.n21265 10.555
R37004 vdd.n19152 vdd.n19151 10.555
R37005 vdd.n21004 vdd.n21003 10.555
R37006 vdd.n18884 vdd.n18881 10.555
R37007 vdd.n18643 vdd.n18640 10.555
R37008 vdd.n18625 vdd.n18622 10.555
R37009 vdd.n32239 vdd.n32238 10.541
R37010 vdd.n2575 vdd.n2574 10.541
R37011 vdd.n9261 vdd.n9260 10.541
R37012 vdd.n21627 vdd.n21625 10.541
R37013 vdd.n14194 vdd.t130 10.399
R37014 vdd.n32478 vdd.n32477 10.278
R37015 vdd.n13012 vdd.n9401 10.27
R37016 vdd.n9540 vdd.t308 10.27
R37017 vdd.n9594 vdd.n9593 10.27
R37018 vdd.n12804 vdd.n9761 10.27
R37019 vdd.n9954 vdd.n9953 10.27
R37020 vdd.n10112 vdd.n10111 10.27
R37021 vdd.n12001 vdd.t291 10.27
R37022 vdd.n16628 vdd.n16626 10.27
R37023 vdd.n18257 vdd.t250 10.27
R37024 vdd.n3940 vdd.n3939 10.184
R37025 vdd.n31947 vdd.n31944 10.164
R37026 vdd.n2023 vdd.n2022 10.164
R37027 vdd.n10472 vdd.n10471 10.144
R37028 vdd.n13446 vdd.t334 10.093
R37029 vdd.n22202 vdd.n22201 10.035
R37030 vdd.n22060 vdd.n22059 10.035
R37031 vdd.n12956 vdd.n9474 9.949
R37032 vdd.n12851 vdd.n9669 9.949
R37033 vdd.n12748 vdd.n9834 9.949
R37034 vdd.n12643 vdd.n10029 9.949
R37035 vdd.t385 vdd.n12277 9.949
R37036 vdd.n15751 vdd.n15750 9.949
R37037 vdd.n16007 vdd.n16006 9.949
R37038 vdd.n16263 vdd.n16262 9.949
R37039 vdd.n16519 vdd.n16518 9.949
R37040 vdd.n21609 vdd.n21607 9.851
R37041 vdd.n21414 vdd.n21413 9.851
R37042 vdd.n21365 vdd.n21364 9.851
R37043 vdd.n21155 vdd.n21154 9.851
R37044 vdd.n21106 vdd.n21105 9.851
R37045 vdd.n19048 vdd.n19047 9.851
R37046 vdd.n18999 vdd.n18998 9.851
R37047 vdd.n18789 vdd.n18788 9.851
R37048 vdd.n18740 vdd.n18739 9.851
R37049 vdd.n18530 vdd.n18529 9.851
R37050 vdd.n35880 vdd.n35879 9.827
R37051 vdd.n35957 vdd.n35956 9.827
R37052 vdd.n36111 vdd.n36110 9.827
R37053 vdd.n36188 vdd.n36187 9.827
R37054 vdd.n36342 vdd.n36341 9.827
R37055 vdd.n36419 vdd.n36418 9.827
R37056 vdd.n36573 vdd.n36572 9.827
R37057 vdd.n36650 vdd.n36649 9.827
R37058 vdd.n36804 vdd.n36803 9.827
R37059 vdd.n36881 vdd.n36880 9.827
R37060 vdd.n33281 vdd.n33280 9.827
R37061 vdd.n33215 vdd.n33214 9.827
R37062 vdd.n37217 vdd.n37216 9.827
R37063 vdd.n37274 vdd.n37273 9.827
R37064 vdd.n37415 vdd.n37414 9.827
R37065 vdd.n37477 vdd.n37476 9.827
R37066 vdd.n38163 vdd.n38162 9.827
R37067 vdd.n38090 vdd.n38089 9.827
R37068 vdd.n37936 vdd.n37935 9.827
R37069 vdd.n37859 vdd.n37858 9.827
R37070 vdd.n37705 vdd.n37704 9.827
R37071 vdd.n37628 vdd.n37627 9.827
R37072 vdd.n28301 vdd.n28300 9.827
R37073 vdd.n28378 vdd.n28377 9.827
R37074 vdd.n28532 vdd.n28531 9.827
R37075 vdd.n28609 vdd.n28608 9.827
R37076 vdd.n28763 vdd.n28762 9.827
R37077 vdd.n28170 vdd.n28169 9.827
R37078 vdd.n28985 vdd.n28984 9.827
R37079 vdd.n27789 vdd.n27788 9.827
R37080 vdd.n31570 vdd.n31569 9.827
R37081 vdd.n29814 vdd.n29813 9.827
R37082 vdd.n30269 vdd.n30268 9.827
R37083 vdd.n30528 vdd.n30527 9.827
R37084 vdd.n2769 vdd.n2768 9.827
R37085 vdd.n2830 vdd.n2829 9.827
R37086 vdd.n2950 vdd.n2949 9.827
R37087 vdd.n3011 vdd.n3010 9.827
R37088 vdd.n3131 vdd.n3130 9.827
R37089 vdd.n3192 vdd.n3191 9.827
R37090 vdd.n3312 vdd.n3311 9.827
R37091 vdd.n3373 vdd.n3372 9.827
R37092 vdd.n3493 vdd.n3492 9.827
R37093 vdd.n3554 vdd.n3553 9.827
R37094 vdd.n2717 vdd.n2716 9.827
R37095 vdd.n3979 vdd.n3978 9.827
R37096 vdd.n2174 vdd.n2173 9.827
R37097 vdd.n2338 vdd.n2337 9.827
R37098 vdd.n2653 vdd.n2652 9.827
R37099 vdd.n1936 vdd.n1935 9.827
R37100 vdd.n1767 vdd.n1766 9.827
R37101 vdd.n1712 vdd.n1711 9.827
R37102 vdd.n1592 vdd.n1591 9.827
R37103 vdd.n1531 vdd.n1530 9.827
R37104 vdd.n1411 vdd.n1410 9.827
R37105 vdd.n1350 vdd.n1349 9.827
R37106 vdd.n26816 vdd.n26815 9.827
R37107 vdd.n26877 vdd.n26876 9.827
R37108 vdd.n26997 vdd.n26996 9.827
R37109 vdd.n27058 vdd.n27057 9.827
R37110 vdd.n27178 vdd.n27177 9.827
R37111 vdd.n26752 vdd.n26751 9.827
R37112 vdd.n31821 vdd.n31820 9.827
R37113 vdd.n31672 vdd.n31671 9.827
R37114 vdd.n31566 vdd.n31565 9.827
R37115 vdd.n31522 vdd.n31521 9.827
R37116 vdd.n31046 vdd.n31045 9.827
R37117 vdd.n31255 vdd.n31254 9.827
R37118 vdd.n13189 vdd.n9221 9.827
R37119 vdd.n13288 vdd.n9149 9.827
R37120 vdd.n13483 vdd.n9001 9.827
R37121 vdd.n13580 vdd.n8928 9.827
R37122 vdd.n13763 vdd.n8784 9.827
R37123 vdd.n13848 vdd.n8722 9.827
R37124 vdd.n14039 vdd.n8558 9.827
R37125 vdd.n14137 vdd.n8501 9.827
R37126 vdd.n14346 vdd.n8341 9.827
R37127 vdd.n8251 vdd.n8243 9.827
R37128 vdd.n14655 vdd.n8148 9.827
R37129 vdd.n14772 vdd.n8084 9.827
R37130 vdd.n14827 vdd.n8057 9.827
R37131 vdd.n14941 vdd.n8002 9.827
R37132 vdd.n13160 vdd.n9234 9.827
R37133 vdd.n13364 vdd.n9073 9.827
R37134 vdd.n13454 vdd.n9010 9.827
R37135 vdd.n13656 vdd.n8853 9.827
R37136 vdd.n13744 vdd.n8791 9.827
R37137 vdd.n13936 vdd.n8641 9.827
R37138 vdd.n14023 vdd.n8575 9.827
R37139 vdd.n14226 vdd.n8419 9.827
R37140 vdd.n14318 vdd.n8358 9.827
R37141 vdd.n14558 vdd.n8189 9.827
R37142 vdd.n19378 vdd.n19377 9.827
R37143 vdd.n19459 vdd.n19458 9.827
R37144 vdd.n19584 vdd.n19583 9.827
R37145 vdd.n19659 vdd.n19658 9.827
R37146 vdd.n19786 vdd.n19785 9.827
R37147 vdd.n20983 vdd.n20982 9.827
R37148 vdd.n19885 vdd.n19884 9.827
R37149 vdd.n20792 vdd.n20791 9.827
R37150 vdd.n20668 vdd.n20667 9.827
R37151 vdd.n20587 vdd.n20586 9.827
R37152 vdd.n21603 vdd.n21602 9.827
R37153 vdd.n21425 vdd.n21424 9.827
R37154 vdd.n21344 vdd.n21343 9.827
R37155 vdd.n21166 vdd.n21165 9.827
R37156 vdd.n21081 vdd.n21080 9.827
R37157 vdd.n19059 vdd.n19058 9.827
R37158 vdd.n18978 vdd.n18977 9.827
R37159 vdd.n18800 vdd.n18799 9.827
R37160 vdd.n18719 vdd.n18718 9.827
R37161 vdd.n18541 vdd.n18540 9.827
R37162 vdd.n20469 vdd.n19980 9.827
R37163 vdd.n20299 vdd.n20293 9.827
R37164 vdd.n20249 vdd.n20243 9.827
R37165 vdd.n20063 vdd.n20030 9.827
R37166 vdd.n24679 vdd.n24678 9.827
R37167 vdd.n25234 vdd.n25233 9.827
R37168 vdd.t327 vdd.n8835 9.787
R37169 vdd.n12512 vdd.n10530 9.702
R37170 vdd.n10632 vdd.n10616 9.702
R37171 vdd.n12402 vdd.n10707 9.702
R37172 vdd.n12363 vdd.n10776 9.702
R37173 vdd.n12308 vdd.n10895 9.702
R37174 vdd.n10986 vdd.n10968 9.702
R37175 vdd.n11073 vdd.n11064 9.702
R37176 vdd.n12153 vdd.n11135 9.702
R37177 vdd.n11233 vdd.n11222 9.702
R37178 vdd.n12057 vdd.n11284 9.702
R37179 vdd.n12002 vdd.n11404 9.702
R37180 vdd.n11529 vdd.n11525 9.702
R37181 vdd.n10414 vdd.n10315 9.702
R37182 vdd.n13070 vdd.n9296 9.702
R37183 vdd.n9397 vdd.n9362 9.702
R37184 vdd.n9484 vdd.n9463 9.702
R37185 vdd.n12908 vdd.n12907 9.702
R37186 vdd.n12862 vdd.n9657 9.702
R37187 vdd.n9757 vdd.n9722 9.702
R37188 vdd.n9844 vdd.n9823 9.702
R37189 vdd.n12700 vdd.n12699 9.702
R37190 vdd.n12654 vdd.n10017 9.702
R37191 vdd.n12604 vdd.n10064 9.702
R37192 vdd.n16916 vdd.n16910 9.702
R37193 vdd.n17040 vdd.n17034 9.702
R37194 vdd.n17188 vdd.n17182 9.702
R37195 vdd.n17312 vdd.n17306 9.702
R37196 vdd.n17460 vdd.n17454 9.702
R37197 vdd.n17584 vdd.n17578 9.702
R37198 vdd.n17718 vdd.n17712 9.702
R37199 vdd.n17842 vdd.n17836 9.702
R37200 vdd.n17989 vdd.n17983 9.702
R37201 vdd.n18113 vdd.n18107 9.702
R37202 vdd.n18258 vdd.n18253 9.702
R37203 vdd.n18366 vdd.n18362 9.702
R37204 vdd.n15364 vdd.n15363 9.702
R37205 vdd.n15472 vdd.n15471 9.702
R37206 vdd.n15603 vdd.n15602 9.702
R37207 vdd.n15728 vdd.n15727 9.702
R37208 vdd.n15859 vdd.n15858 9.702
R37209 vdd.n15984 vdd.n15983 9.702
R37210 vdd.n16115 vdd.n16114 9.702
R37211 vdd.n16240 vdd.n16239 9.702
R37212 vdd.n16371 vdd.n16370 9.702
R37213 vdd.n16496 vdd.n16495 9.702
R37214 vdd.n16699 vdd.n16698 9.702
R37215 vdd.n2497 vdd.n2450 9.669
R37216 vdd.n9320 vdd.t212 9.628
R37217 vdd.n13001 vdd.n13000 9.628
R37218 vdd.n12899 vdd.n9570 9.628
R37219 vdd.n12793 vdd.n12792 9.628
R37220 vdd.n12691 vdd.n9929 9.628
R37221 vdd.t83 vdd.n12594 9.628
R37222 vdd.t181 vdd.n15494 9.628
R37223 vdd.n16640 vdd.t337 9.628
R37224 vdd.n2582 vdd.n2581 9.565
R37225 vdd.n2446 vdd.n2445 9.554
R37226 vdd.n2588 vdd.n2587 9.552
R37227 vdd.n3829 vdd.n3828 9.544
R37228 vdd.n3796 vdd.n3795 9.543
R37229 vdd.n3788 vdd.n3787 9.525
R37230 vdd.n13960 vdd.t108 9.481
R37231 vdd.n12598 vdd.n10067 9.459
R37232 vdd.n16682 vdd.n16681 9.459
R37233 vdd.n11882 vdd.n11799 9.43
R37234 vdd.n21973 vdd.n21890 9.43
R37235 vdd.n11729 vdd.n11728 9.413
R37236 vdd.n21802 vdd.n21801 9.413
R37237 vdd.n26184 vdd.n26183 9.403
R37238 vdd.n31647 vdd.n31646 9.399
R37239 vdd.n32491 vdd.n32490 9.386
R37240 vdd.n19418 vdd.n19414 9.382
R37241 vdd.n19432 vdd.n19431 9.382
R37242 vdd.n19621 vdd.n19617 9.382
R37243 vdd.n19823 vdd.n19819 9.382
R37244 vdd.n19170 vdd.n19169 9.382
R37245 vdd.n20826 vdd.n20825 9.382
R37246 vdd.n20641 vdd.n20637 9.382
R37247 vdd.n20624 vdd.n20623 9.382
R37248 vdd.n19997 vdd.n19996 9.382
R37249 vdd.n20009 vdd.n20006 9.382
R37250 vdd.n14787 vdd.n8073 9.359
R37251 vdd.n14781 vdd.n14780 9.359
R37252 vdd.n24690 vdd.n24689 9.332
R37253 vdd.n25221 vdd.n25220 9.332
R37254 vdd.n24689 vdd.n24688 9.332
R37255 vdd.n25220 vdd.n25219 9.332
R37256 vdd.n13050 vdd.n13049 9.307
R37257 vdd.n12949 vdd.n12948 9.307
R37258 vdd.n12741 vdd.n12740 9.307
R37259 vdd.n12634 vdd.n12633 9.307
R37260 vdd.n15512 vdd.n15511 9.307
R37261 vdd.n15768 vdd.n15767 9.307
R37262 vdd.n16280 vdd.n16279 9.307
R37263 vdd.n16536 vdd.n16535 9.307
R37264 vdd.n25666 vdd.n25665 9.306
R37265 vdd.n25601 vdd.n25426 9.306
R37266 vdd.n24519 vdd.n24518 9.303
R37267 vdd.n1886 vdd.n1225 9.301
R37268 vdd.n33802 vdd.n33801 9.3
R37269 vdd.n33814 vdd.n33813 9.3
R37270 vdd.n33812 vdd.n33811 9.3
R37271 vdd.n33826 vdd.n33825 9.3
R37272 vdd.n33824 vdd.n33823 9.3
R37273 vdd.n33846 vdd.n33845 9.3
R37274 vdd.n33791 vdd.n33790 9.3
R37275 vdd.n33782 vdd.n33781 9.3
R37276 vdd.n33794 vdd.n33793 9.3
R37277 vdd.n33601 vdd.n33600 9.3
R37278 vdd.n33598 vdd.n33597 9.3
R37279 vdd.n33610 vdd.n33609 9.3
R37280 vdd.n33622 vdd.n33621 9.3
R37281 vdd.n33633 vdd.n33632 9.3
R37282 vdd.n33646 vdd.n33645 9.3
R37283 vdd.n33644 vdd.n33643 9.3
R37284 vdd.n33658 vdd.n33657 9.3
R37285 vdd.n33656 vdd.n33655 9.3
R37286 vdd.n33680 vdd.n33679 9.3
R37287 vdd.n33691 vdd.n33690 9.3
R37288 vdd.n33689 vdd.n33688 9.3
R37289 vdd.n33495 vdd.n33494 9.3
R37290 vdd.n33507 vdd.n33506 9.3
R37291 vdd.n33528 vdd.n33527 9.3
R37292 vdd.n33530 vdd.n33529 9.3
R37293 vdd.n33309 vdd.n33308 9.3
R37294 vdd.n33322 vdd.n33321 9.3
R37295 vdd.n33320 vdd.n33319 9.3
R37296 vdd.n33334 vdd.n33333 9.3
R37297 vdd.n33332 vdd.n33331 9.3
R37298 vdd.n33356 vdd.n33355 9.3
R37299 vdd.n33465 vdd.n33464 9.3
R37300 vdd.n33447 vdd.n33446 9.3
R37301 vdd.n33445 vdd.n33444 9.3
R37302 vdd.n33412 vdd.n33411 9.3
R37303 vdd.n33410 vdd.n33409 9.3
R37304 vdd.n33416 vdd.n33415 9.3
R37305 vdd.n34166 vdd.n34165 9.3
R37306 vdd.n34178 vdd.n34177 9.3
R37307 vdd.n34176 vdd.n34175 9.3
R37308 vdd.n34215 vdd.n34214 9.3
R37309 vdd.n34226 vdd.n34225 9.3
R37310 vdd.n34256 vdd.n34255 9.3
R37311 vdd.n34254 vdd.n34253 9.3
R37312 vdd.n34273 vdd.n34272 9.3
R37313 vdd.n34284 vdd.n34283 9.3
R37314 vdd.n34297 vdd.n34296 9.3
R37315 vdd.n34295 vdd.n34294 9.3
R37316 vdd.n34333 vdd.n34332 9.3
R37317 vdd.n33952 vdd.n33951 9.3
R37318 vdd.n33878 vdd.n33877 9.3
R37319 vdd.n33919 vdd.n33918 9.3
R37320 vdd.n33917 vdd.n33916 9.3
R37321 vdd.n33926 vdd.n33925 9.3
R37322 vdd.n34402 vdd.n34401 9.3
R37323 vdd.n34357 vdd.n34356 9.3
R37324 vdd.n34056 vdd.n34055 9.3
R37325 vdd.n33998 vdd.n33997 9.3
R37326 vdd.n33996 vdd.n33995 9.3
R37327 vdd.n34224 vdd.n34223 9.3
R37328 vdd.n34112 vdd.n34111 9.3
R37329 vdd.n34331 vdd.n34330 9.3
R37330 vdd.n34427 vdd.n34426 9.3
R37331 vdd.n33950 vdd.n33949 9.3
R37332 vdd.n33880 vdd.n33879 9.3
R37333 vdd.n34054 vdd.n34053 9.3
R37334 vdd.n34003 vdd.n34002 9.3
R37335 vdd.n34007 vdd.n34006 9.3
R37336 vdd.n35308 vdd.n35307 9.3
R37337 vdd.n35169 vdd.n35168 9.3
R37338 vdd.n35165 vdd.n35164 9.3
R37339 vdd.n35160 vdd.n35159 9.3
R37340 vdd.n35158 vdd.n35157 9.3
R37341 vdd.n35217 vdd.n35216 9.3
R37342 vdd.n35215 vdd.n35214 9.3
R37343 vdd.n35038 vdd.n35037 9.3
R37344 vdd.n35103 vdd.n35102 9.3
R37345 vdd.n35036 vdd.n35035 9.3
R37346 vdd.n35105 vdd.n35104 9.3
R37347 vdd.n35065 vdd.n35064 9.3
R37348 vdd.n35063 vdd.n35062 9.3
R37349 vdd.n35052 vdd.n35051 9.3
R37350 vdd.n35417 vdd.n35416 9.3
R37351 vdd.n35373 vdd.n35372 9.3
R37352 vdd.n35385 vdd.n35384 9.3
R37353 vdd.n35599 vdd.n35598 9.3
R37354 vdd.n35597 vdd.n35596 9.3
R37355 vdd.n35563 vdd.n35562 9.3
R37356 vdd.n35561 vdd.n35560 9.3
R37357 vdd.n35550 vdd.n35549 9.3
R37358 vdd.n35539 vdd.n35538 9.3
R37359 vdd.n35522 vdd.n35521 9.3
R37360 vdd.n35520 vdd.n35519 9.3
R37361 vdd.n35497 vdd.n35496 9.3
R37362 vdd.n35335 vdd.n35334 9.3
R37363 vdd.n35347 vdd.n35346 9.3
R37364 vdd.n35345 vdd.n35344 9.3
R37365 vdd.n35323 vdd.n35322 9.3
R37366 vdd.n35321 vdd.n35320 9.3
R37367 vdd.n34732 vdd.n34731 9.3
R37368 vdd.n34728 vdd.n34727 9.3
R37369 vdd.n34726 vdd.n34725 9.3
R37370 vdd.n34751 vdd.n34750 9.3
R37371 vdd.n34763 vdd.n34762 9.3
R37372 vdd.n34937 vdd.n34936 9.3
R37373 vdd.n34935 vdd.n34934 9.3
R37374 vdd.n34928 vdd.n34927 9.3
R37375 vdd.n34920 vdd.n34919 9.3
R37376 vdd.n34913 vdd.n34912 9.3
R37377 vdd.n34911 vdd.n34910 9.3
R37378 vdd.n35011 vdd.n35010 9.3
R37379 vdd.n34454 vdd.n34453 9.3
R37380 vdd.n34516 vdd.n34515 9.3
R37381 vdd.n34478 vdd.n34477 9.3
R37382 vdd.n34476 vdd.n34475 9.3
R37383 vdd.n34465 vdd.n34464 9.3
R37384 vdd.n34821 vdd.n34820 9.3
R37385 vdd.n34783 vdd.n34782 9.3
R37386 vdd.n34630 vdd.n34629 9.3
R37387 vdd.n34578 vdd.n34577 9.3
R37388 vdd.n34576 vdd.n34575 9.3
R37389 vdd.n34761 vdd.n34760 9.3
R37390 vdd.n34945 vdd.n34944 9.3
R37391 vdd.n35009 vdd.n35008 9.3
R37392 vdd.n34857 vdd.n34856 9.3
R37393 vdd.n34452 vdd.n34451 9.3
R37394 vdd.n34518 vdd.n34517 9.3
R37395 vdd.n34628 vdd.n34627 9.3
R37396 vdd.n34585 vdd.n34584 9.3
R37397 vdd.n34591 vdd.n34590 9.3
R37398 vdd.n826 vdd.n825 9.3
R37399 vdd.n822 vdd.n821 9.3
R37400 vdd.n820 vdd.n819 9.3
R37401 vdd.n837 vdd.n836 9.3
R37402 vdd.n840 vdd.n839 9.3
R37403 vdd.n847 vdd.n846 9.3
R37404 vdd.n858 vdd.n857 9.3
R37405 vdd.n868 vdd.n867 9.3
R37406 vdd.n856 vdd.n855 9.3
R37407 vdd.n1112 vdd.n1111 9.3
R37408 vdd.n1109 vdd.n1108 9.3
R37409 vdd.n1103 vdd.n1102 9.3
R37410 vdd.n1098 vdd.n1097 9.3
R37411 vdd.n1090 vdd.n1089 9.3
R37412 vdd.n1083 vdd.n1082 9.3
R37413 vdd.n1081 vdd.n1080 9.3
R37414 vdd.n1074 vdd.n1073 9.3
R37415 vdd.n1072 vdd.n1071 9.3
R37416 vdd.n1145 vdd.n1144 9.3
R37417 vdd.n1157 vdd.n1156 9.3
R37418 vdd.n1155 vdd.n1154 9.3
R37419 vdd.n985 vdd.n984 9.3
R37420 vdd.n1031 vdd.n1030 9.3
R37421 vdd.n1011 vdd.n1010 9.3
R37422 vdd.n1013 vdd.n1012 9.3
R37423 vdd.n638 vdd.n637 9.3
R37424 vdd.n632 vdd.n631 9.3
R37425 vdd.n630 vdd.n629 9.3
R37426 vdd.n623 vdd.n622 9.3
R37427 vdd.n621 vdd.n620 9.3
R37428 vdd.n674 vdd.n673 9.3
R37429 vdd.n784 vdd.n783 9.3
R37430 vdd.n766 vdd.n765 9.3
R37431 vdd.n764 vdd.n763 9.3
R37432 vdd.n736 vdd.n735 9.3
R37433 vdd.n734 vdd.n733 9.3
R37434 vdd.n742 vdd.n741 9.3
R37435 vdd.n327 vdd.n326 9.3
R37436 vdd.n339 vdd.n338 9.3
R37437 vdd.n337 vdd.n336 9.3
R37438 vdd.n351 vdd.n350 9.3
R37439 vdd.n349 vdd.n348 9.3
R37440 vdd.n373 vdd.n372 9.3
R37441 vdd.n311 vdd.n310 9.3
R37442 vdd.n214 vdd.n213 9.3
R37443 vdd.n309 vdd.n308 9.3
R37444 vdd.n100 vdd.n99 9.3
R37445 vdd.n97 vdd.n96 9.3
R37446 vdd.n109 vdd.n108 9.3
R37447 vdd.n121 vdd.n120 9.3
R37448 vdd.n132 vdd.n131 9.3
R37449 vdd.n145 vdd.n144 9.3
R37450 vdd.n143 vdd.n142 9.3
R37451 vdd.n157 vdd.n156 9.3
R37452 vdd.n155 vdd.n154 9.3
R37453 vdd.n179 vdd.n178 9.3
R37454 vdd.n191 vdd.n190 9.3
R37455 vdd.n189 vdd.n188 9.3
R37456 vdd.n18 vdd.n17 9.3
R37457 vdd.n32 vdd.n31 9.3
R37458 vdd.n20 vdd.n19 9.3
R37459 vdd.n30 vdd.n29 9.3
R37460 vdd.n52 vdd.n51 9.3
R37461 vdd.n54 vdd.n53 9.3
R37462 vdd.n394 vdd.n393 9.3
R37463 vdd.n396 vdd.n395 9.3
R37464 vdd.n414 vdd.n413 9.3
R37465 vdd.n427 vdd.n426 9.3
R37466 vdd.n425 vdd.n424 9.3
R37467 vdd.n461 vdd.n460 9.3
R37468 vdd.n479 vdd.n478 9.3
R37469 vdd.n459 vdd.n458 9.3
R37470 vdd.n566 vdd.n565 9.3
R37471 vdd.n525 vdd.n524 9.3
R37472 vdd.n523 vdd.n522 9.3
R37473 vdd.n532 vdd.n531 9.3
R37474 vdd.n530 vdd.n529 9.3
R37475 vdd.n536 vdd.n535 9.3
R37476 vdd.n5867 vdd.n5866 9.3
R37477 vdd.n6302 vdd.n6301 9.3
R37478 vdd.n6296 vdd.n6295 9.3
R37479 vdd.n6289 vdd.n6288 9.3
R37480 vdd.n6287 vdd.n6286 9.3
R37481 vdd.n6341 vdd.n6340 9.3
R37482 vdd.n6339 vdd.n6338 9.3
R37483 vdd.n6236 vdd.n6235 9.3
R37484 vdd.n6152 vdd.n6151 9.3
R37485 vdd.n6234 vdd.n6233 9.3
R37486 vdd.n6154 vdd.n6153 9.3
R37487 vdd.n6193 vdd.n6192 9.3
R37488 vdd.n6191 vdd.n6190 9.3
R37489 vdd.n6200 vdd.n6199 9.3
R37490 vdd.n6207 vdd.n6206 9.3
R37491 vdd.n6063 vdd.n6062 9.3
R37492 vdd.n6078 vdd.n6077 9.3
R37493 vdd.n6034 vdd.n6033 9.3
R37494 vdd.n6032 vdd.n6031 9.3
R37495 vdd.n5956 vdd.n5955 9.3
R37496 vdd.n5954 vdd.n5953 9.3
R37497 vdd.n5963 vdd.n5962 9.3
R37498 vdd.n5971 vdd.n5970 9.3
R37499 vdd.n5980 vdd.n5979 9.3
R37500 vdd.n5978 vdd.n5977 9.3
R37501 vdd.n5998 vdd.n5997 9.3
R37502 vdd.n5916 vdd.n5915 9.3
R37503 vdd.n5853 vdd.n5852 9.3
R37504 vdd.n5851 vdd.n5850 9.3
R37505 vdd.n5881 vdd.n5880 9.3
R37506 vdd.n5879 vdd.n5878 9.3
R37507 vdd.n5479 vdd.n5478 9.3
R37508 vdd.n5475 vdd.n5474 9.3
R37509 vdd.n5473 vdd.n5472 9.3
R37510 vdd.n5498 vdd.n5497 9.3
R37511 vdd.n5510 vdd.n5509 9.3
R37512 vdd.n5684 vdd.n5683 9.3
R37513 vdd.n5682 vdd.n5681 9.3
R37514 vdd.n5675 vdd.n5674 9.3
R37515 vdd.n5667 vdd.n5666 9.3
R37516 vdd.n5660 vdd.n5659 9.3
R37517 vdd.n5658 vdd.n5657 9.3
R37518 vdd.n5758 vdd.n5757 9.3
R37519 vdd.n5201 vdd.n5200 9.3
R37520 vdd.n5263 vdd.n5262 9.3
R37521 vdd.n5225 vdd.n5224 9.3
R37522 vdd.n5223 vdd.n5222 9.3
R37523 vdd.n5212 vdd.n5211 9.3
R37524 vdd.n5568 vdd.n5567 9.3
R37525 vdd.n5530 vdd.n5529 9.3
R37526 vdd.n5377 vdd.n5376 9.3
R37527 vdd.n5325 vdd.n5324 9.3
R37528 vdd.n5323 vdd.n5322 9.3
R37529 vdd.n5508 vdd.n5507 9.3
R37530 vdd.n5692 vdd.n5691 9.3
R37531 vdd.n5756 vdd.n5755 9.3
R37532 vdd.n5604 vdd.n5603 9.3
R37533 vdd.n5199 vdd.n5198 9.3
R37534 vdd.n5265 vdd.n5264 9.3
R37535 vdd.n5375 vdd.n5374 9.3
R37536 vdd.n5332 vdd.n5331 9.3
R37537 vdd.n5338 vdd.n5337 9.3
R37538 vdd.n4903 vdd.n4902 9.3
R37539 vdd.n4652 vdd.n4651 9.3
R37540 vdd.n4647 vdd.n4646 9.3
R37541 vdd.n4642 vdd.n4641 9.3
R37542 vdd.n4640 vdd.n4639 9.3
R37543 vdd.n4698 vdd.n4697 9.3
R37544 vdd.n4696 vdd.n4695 9.3
R37545 vdd.n4776 vdd.n4775 9.3
R37546 vdd.n4719 vdd.n4718 9.3
R37547 vdd.n4731 vdd.n4730 9.3
R37548 vdd.n5001 vdd.n5000 9.3
R37549 vdd.n4996 vdd.n4995 9.3
R37550 vdd.n4994 vdd.n4993 9.3
R37551 vdd.n4961 vdd.n4960 9.3
R37552 vdd.n5042 vdd.n5041 9.3
R37553 vdd.n4963 vdd.n4962 9.3
R37554 vdd.n5040 vdd.n5039 9.3
R37555 vdd.n5171 vdd.n5170 9.3
R37556 vdd.n5169 vdd.n5168 9.3
R37557 vdd.n5134 vdd.n5133 9.3
R37558 vdd.n5132 vdd.n5131 9.3
R37559 vdd.n5123 vdd.n5122 9.3
R37560 vdd.n5112 vdd.n5111 9.3
R37561 vdd.n5094 vdd.n5093 9.3
R37562 vdd.n5092 vdd.n5091 9.3
R37563 vdd.n4929 vdd.n4928 9.3
R37564 vdd.n4941 vdd.n4940 9.3
R37565 vdd.n4927 vdd.n4876 9.3
R37566 vdd.n4939 vdd.n4938 9.3
R37567 vdd.n4917 vdd.n4916 9.3
R37568 vdd.n4915 vdd.n4914 9.3
R37569 vdd.n4306 vdd.n4305 9.3
R37570 vdd.n4302 vdd.n4301 9.3
R37571 vdd.n4300 vdd.n4299 9.3
R37572 vdd.n4325 vdd.n4324 9.3
R37573 vdd.n4337 vdd.n4336 9.3
R37574 vdd.n4511 vdd.n4510 9.3
R37575 vdd.n4509 vdd.n4508 9.3
R37576 vdd.n4502 vdd.n4501 9.3
R37577 vdd.n4494 vdd.n4493 9.3
R37578 vdd.n4487 vdd.n4486 9.3
R37579 vdd.n4485 vdd.n4484 9.3
R37580 vdd.n4588 vdd.n4587 9.3
R37581 vdd.n4031 vdd.n4030 9.3
R37582 vdd.n4093 vdd.n4092 9.3
R37583 vdd.n4055 vdd.n4054 9.3
R37584 vdd.n4053 vdd.n4052 9.3
R37585 vdd.n4042 vdd.n4041 9.3
R37586 vdd.n4394 vdd.n4393 9.3
R37587 vdd.n4357 vdd.n4356 9.3
R37588 vdd.n4207 vdd.n4206 9.3
R37589 vdd.n4156 vdd.n4155 9.3
R37590 vdd.n4154 vdd.n4153 9.3
R37591 vdd.n4335 vdd.n4334 9.3
R37592 vdd.n4519 vdd.n4518 9.3
R37593 vdd.n4586 vdd.n4585 9.3
R37594 vdd.n4431 vdd.n4430 9.3
R37595 vdd.n4029 vdd.n4028 9.3
R37596 vdd.n4095 vdd.n4094 9.3
R37597 vdd.n4205 vdd.n4204 9.3
R37598 vdd.n4163 vdd.n4162 9.3
R37599 vdd.n4169 vdd.n4168 9.3
R37600 vdd.n37582 vdd.n37580 9.3
R37601 vdd.n37557 vdd.n37555 9.3
R37602 vdd.n32817 vdd.n32815 9.3
R37603 vdd.n35658 vdd.n35656 9.3
R37604 vdd.n37491 vdd.n37489 9.3
R37605 vdd.n32886 vdd.n32884 9.3
R37606 vdd.n32902 vdd.n32900 9.3
R37607 vdd.n37453 vdd.n37451 9.3
R37608 vdd.n37370 vdd.n37368 9.3
R37609 vdd.n37359 vdd.n37357 9.3
R37610 vdd.n35648 vdd.n35646 9.3
R37611 vdd.n37337 vdd.n37330 9.3
R37612 vdd.n33026 vdd.n33024 9.3
R37613 vdd.n33047 vdd.n33045 9.3
R37614 vdd.n37247 vdd.n37245 9.3
R37615 vdd.n33084 vdd.n33079 9.3
R37616 vdd.n37183 vdd.n37181 9.3
R37617 vdd.n35629 vdd.n35622 9.3
R37618 vdd.n37166 vdd.n37159 9.3
R37619 vdd.n33159 vdd.n33152 9.3
R37620 vdd.n33208 vdd.n33206 9.3
R37621 vdd.n37085 vdd.n37080 9.3
R37622 vdd.n33237 vdd.n33232 9.3
R37623 vdd.n37072 vdd.n37067 9.3
R37624 vdd.n36995 vdd.n36993 9.3
R37625 vdd.n36981 vdd.n36979 9.3
R37626 vdd.n36978 vdd.n36976 9.3
R37627 vdd.n36986 vdd.n36983 9.3
R37628 vdd.n36992 vdd.n36990 9.3
R37629 vdd.n37000 vdd.n36997 9.3
R37630 vdd.n37014 vdd.n37012 9.3
R37631 vdd.n37029 vdd.n37027 9.3
R37632 vdd.n37061 vdd.n37049 9.3
R37633 vdd.n33271 vdd.n33259 9.3
R37634 vdd.n37075 vdd.n37066 9.3
R37635 vdd.n37070 vdd.n37068 9.3
R37636 vdd.n33240 vdd.n33231 9.3
R37637 vdd.n33235 vdd.n33233 9.3
R37638 vdd.n37088 vdd.n37079 9.3
R37639 vdd.n37083 vdd.n37081 9.3
R37640 vdd.n33211 vdd.n33205 9.3
R37641 vdd.n37102 vdd.n37100 9.3
R37642 vdd.n37107 vdd.n37104 9.3
R37643 vdd.n37126 vdd.n37123 9.3
R37644 vdd.n33184 vdd.n33179 9.3
R37645 vdd.n37140 vdd.n37135 9.3
R37646 vdd.n33161 vdd.n33151 9.3
R37647 vdd.n33157 vdd.n33154 9.3
R37648 vdd.n37168 vdd.n37158 9.3
R37649 vdd.n37164 vdd.n37161 9.3
R37650 vdd.n35631 vdd.n35621 9.3
R37651 vdd.n35627 vdd.n35624 9.3
R37652 vdd.n37185 vdd.n37180 9.3
R37653 vdd.n33121 vdd.n33118 9.3
R37654 vdd.n33124 vdd.n33122 9.3
R37655 vdd.n33105 vdd.n33103 9.3
R37656 vdd.n33093 vdd.n33091 9.3
R37657 vdd.n37235 vdd.n37233 9.3
R37658 vdd.n33087 vdd.n33078 9.3
R37659 vdd.n33082 vdd.n33080 9.3
R37660 vdd.n37250 vdd.n37244 9.3
R37661 vdd.n33063 vdd.n33061 9.3
R37662 vdd.n33050 vdd.n33044 9.3
R37663 vdd.n37265 vdd.n37263 9.3
R37664 vdd.n37270 vdd.n37267 9.3
R37665 vdd.n33029 vdd.n33027 9.3
R37666 vdd.n37292 vdd.n37289 9.3
R37667 vdd.n33019 vdd.n33016 9.3
R37668 vdd.n37303 vdd.n37300 9.3
R37669 vdd.n33001 vdd.n32998 9.3
R37670 vdd.n37339 vdd.n37329 9.3
R37671 vdd.n37335 vdd.n37332 9.3
R37672 vdd.n35650 vdd.n35645 9.3
R37673 vdd.n37345 vdd.n37342 9.3
R37674 vdd.n37361 vdd.n37356 9.3
R37675 vdd.n32968 vdd.n32965 9.3
R37676 vdd.n37367 vdd.n37365 9.3
R37677 vdd.n37375 vdd.n37372 9.3
R37678 vdd.n32951 vdd.n32949 9.3
R37679 vdd.n37398 vdd.n37396 9.3
R37680 vdd.n37429 vdd.n37427 9.3
R37681 vdd.n37436 vdd.n37434 9.3
R37682 vdd.n37456 vdd.n37450 9.3
R37683 vdd.n32918 vdd.n32916 9.3
R37684 vdd.n32905 vdd.n32899 9.3
R37685 vdd.n37460 vdd.n37458 9.3
R37686 vdd.n32883 vdd.n32880 9.3
R37687 vdd.n32889 vdd.n32887 9.3
R37688 vdd.n37488 vdd.n37485 9.3
R37689 vdd.n37494 vdd.n37492 9.3
R37690 vdd.n32874 vdd.n32871 9.3
R37691 vdd.n37515 vdd.n37512 9.3
R37692 vdd.n32856 vdd.n32853 9.3
R37693 vdd.n37535 vdd.n37532 9.3
R37694 vdd.n35660 vdd.n35655 9.3
R37695 vdd.n37543 vdd.n37540 9.3
R37696 vdd.n37546 vdd.n37544 9.3
R37697 vdd.n32822 vdd.n32819 9.3
R37698 vdd.n37554 vdd.n37552 9.3
R37699 vdd.n37562 vdd.n37559 9.3
R37700 vdd.n37579 vdd.n37577 9.3
R37701 vdd.n37587 vdd.n37584 9.3
R37702 vdd.n38200 vdd.n37588 9.3
R37703 vdd.n38186 vdd.n37593 9.3
R37704 vdd.n37582 vdd.n37581 9.3
R37705 vdd.n37557 vdd.n37556 9.3
R37706 vdd.n32817 vdd.n32816 9.3
R37707 vdd.n35658 vdd.n35657 9.3
R37708 vdd.n37491 vdd.n37490 9.3
R37709 vdd.n32886 vdd.n32885 9.3
R37710 vdd.n32902 vdd.n32901 9.3
R37711 vdd.n37453 vdd.n37452 9.3
R37712 vdd.n37370 vdd.n37369 9.3
R37713 vdd.n37359 vdd.n37358 9.3
R37714 vdd.n35648 vdd.n35647 9.3
R37715 vdd.n37337 vdd.n37336 9.3
R37716 vdd.n33026 vdd.n33025 9.3
R37717 vdd.n33047 vdd.n33046 9.3
R37718 vdd.n37247 vdd.n37246 9.3
R37719 vdd.n33084 vdd.n33083 9.3
R37720 vdd.n37183 vdd.n37182 9.3
R37721 vdd.n35629 vdd.n35628 9.3
R37722 vdd.n37166 vdd.n37165 9.3
R37723 vdd.n33159 vdd.n33158 9.3
R37724 vdd.n33208 vdd.n33207 9.3
R37725 vdd.n37085 vdd.n37084 9.3
R37726 vdd.n33237 vdd.n33236 9.3
R37727 vdd.n37072 vdd.n37071 9.3
R37728 vdd.n36995 vdd.n36994 9.3
R37729 vdd.n36981 vdd.n36980 9.3
R37730 vdd.n36978 vdd.n36977 9.3
R37731 vdd.n36986 vdd.n36985 9.3
R37732 vdd.n36992 vdd.n36991 9.3
R37733 vdd.n37000 vdd.n36999 9.3
R37734 vdd.n37014 vdd.n37013 9.3
R37735 vdd.n37029 vdd.n37028 9.3
R37736 vdd.n37061 vdd.n37060 9.3
R37737 vdd.n33271 vdd.n33270 9.3
R37738 vdd.n37075 vdd.n37074 9.3
R37739 vdd.n37070 vdd.n37069 9.3
R37740 vdd.n33240 vdd.n33239 9.3
R37741 vdd.n33235 vdd.n33234 9.3
R37742 vdd.n37088 vdd.n37087 9.3
R37743 vdd.n37083 vdd.n37082 9.3
R37744 vdd.n33211 vdd.n33210 9.3
R37745 vdd.n37102 vdd.n37101 9.3
R37746 vdd.n37107 vdd.n37106 9.3
R37747 vdd.n37126 vdd.n37125 9.3
R37748 vdd.n33184 vdd.n33183 9.3
R37749 vdd.n37140 vdd.n37139 9.3
R37750 vdd.n33161 vdd.n33160 9.3
R37751 vdd.n33157 vdd.n33156 9.3
R37752 vdd.n37168 vdd.n37167 9.3
R37753 vdd.n37164 vdd.n37163 9.3
R37754 vdd.n35631 vdd.n35630 9.3
R37755 vdd.n35627 vdd.n35626 9.3
R37756 vdd.n37185 vdd.n37184 9.3
R37757 vdd.n33121 vdd.n33120 9.3
R37758 vdd.n33124 vdd.n33123 9.3
R37759 vdd.n33105 vdd.n33104 9.3
R37760 vdd.n33093 vdd.n33092 9.3
R37761 vdd.n37235 vdd.n37234 9.3
R37762 vdd.n33087 vdd.n33086 9.3
R37763 vdd.n33082 vdd.n33081 9.3
R37764 vdd.n37250 vdd.n37249 9.3
R37765 vdd.n33063 vdd.n33062 9.3
R37766 vdd.n33050 vdd.n33049 9.3
R37767 vdd.n37265 vdd.n37264 9.3
R37768 vdd.n37270 vdd.n37269 9.3
R37769 vdd.n33029 vdd.n33028 9.3
R37770 vdd.n37292 vdd.n37291 9.3
R37771 vdd.n33019 vdd.n33018 9.3
R37772 vdd.n37303 vdd.n37302 9.3
R37773 vdd.n33001 vdd.n33000 9.3
R37774 vdd.n37339 vdd.n37338 9.3
R37775 vdd.n37335 vdd.n37334 9.3
R37776 vdd.n35650 vdd.n35649 9.3
R37777 vdd.n37345 vdd.n37344 9.3
R37778 vdd.n37361 vdd.n37360 9.3
R37779 vdd.n32968 vdd.n32967 9.3
R37780 vdd.n37367 vdd.n37366 9.3
R37781 vdd.n37375 vdd.n37374 9.3
R37782 vdd.n32951 vdd.n32950 9.3
R37783 vdd.n37398 vdd.n37397 9.3
R37784 vdd.n37429 vdd.n37428 9.3
R37785 vdd.n37436 vdd.n37435 9.3
R37786 vdd.n37456 vdd.n37455 9.3
R37787 vdd.n32918 vdd.n32917 9.3
R37788 vdd.n32905 vdd.n32904 9.3
R37789 vdd.n37460 vdd.n37459 9.3
R37790 vdd.n32883 vdd.n32882 9.3
R37791 vdd.n32889 vdd.n32888 9.3
R37792 vdd.n37488 vdd.n37487 9.3
R37793 vdd.n37494 vdd.n37493 9.3
R37794 vdd.n32874 vdd.n32873 9.3
R37795 vdd.n37515 vdd.n37514 9.3
R37796 vdd.n32856 vdd.n32855 9.3
R37797 vdd.n37535 vdd.n37534 9.3
R37798 vdd.n35660 vdd.n35659 9.3
R37799 vdd.n37543 vdd.n37542 9.3
R37800 vdd.n37546 vdd.n37545 9.3
R37801 vdd.n32822 vdd.n32821 9.3
R37802 vdd.n37554 vdd.n37553 9.3
R37803 vdd.n37562 vdd.n37561 9.3
R37804 vdd.n37579 vdd.n37578 9.3
R37805 vdd.n37587 vdd.n37586 9.3
R37806 vdd.n38200 vdd.n38199 9.3
R37807 vdd.n38186 vdd.n38185 9.3
R37808 vdd.n31160 vdd.n31159 9.3
R37809 vdd.n31167 vdd.n31166 9.3
R37810 vdd.n31175 vdd.n31174 9.3
R37811 vdd.n32106 vdd.n32093 9.3
R37812 vdd.n32305 vdd.n32304 9.3
R37813 vdd.n32511 vdd.n32510 9.3
R37814 vdd.n31035 vdd.n31034 9.3
R37815 vdd.n31288 vdd.n31287 9.3
R37816 vdd.n31251 vdd.n31250 9.3
R37817 vdd.n31279 vdd.n31262 9.3
R37818 vdd.n28787 vdd.n28786 9.3
R37819 vdd.n28759 vdd.n28758 9.3
R37820 vdd.n28731 vdd.n28730 9.3
R37821 vdd.n28703 vdd.n28702 9.3
R37822 vdd.n28673 vdd.n28672 9.3
R37823 vdd.n28659 vdd.n28658 9.3
R37824 vdd.n28645 vdd.n28644 9.3
R37825 vdd.n28631 vdd.n28630 9.3
R37826 vdd.n28617 vdd.n28616 9.3
R37827 vdd.n28603 vdd.n28602 9.3
R37828 vdd.n28589 vdd.n28588 9.3
R37829 vdd.n28574 vdd.n28573 9.3
R37830 vdd.n28542 vdd.n28541 9.3
R37831 vdd.n28514 vdd.n28513 9.3
R37832 vdd.n28486 vdd.n28485 9.3
R37833 vdd.n28442 vdd.n28441 9.3
R37834 vdd.n28428 vdd.n28427 9.3
R37835 vdd.n28414 vdd.n28413 9.3
R37836 vdd.n28400 vdd.n28399 9.3
R37837 vdd.n28386 vdd.n28385 9.3
R37838 vdd.n28372 vdd.n28371 9.3
R37839 vdd.n28358 vdd.n28357 9.3
R37840 vdd.n28343 vdd.n28342 9.3
R37841 vdd.n28325 vdd.n28324 9.3
R37842 vdd.n28297 vdd.n28296 9.3
R37843 vdd.n28269 vdd.n28268 9.3
R37844 vdd.n28241 vdd.n28240 9.3
R37845 vdd.n28211 vdd.n28210 9.3
R37846 vdd.n28197 vdd.n28196 9.3
R37847 vdd.n28183 vdd.n28182 9.3
R37848 vdd.n37610 vdd.n37609 9.3
R37849 vdd.n37624 vdd.n37623 9.3
R37850 vdd.n37638 vdd.n37637 9.3
R37851 vdd.n37652 vdd.n37651 9.3
R37852 vdd.n37666 vdd.n37665 9.3
R37853 vdd.n37699 vdd.n37698 9.3
R37854 vdd.n37727 vdd.n37726 9.3
R37855 vdd.n37755 vdd.n37754 9.3
R37856 vdd.n37799 vdd.n37798 9.3
R37857 vdd.n37813 vdd.n37812 9.3
R37858 vdd.n37827 vdd.n37826 9.3
R37859 vdd.n37841 vdd.n37840 9.3
R37860 vdd.n37855 vdd.n37854 9.3
R37861 vdd.n37869 vdd.n37868 9.3
R37862 vdd.n37883 vdd.n37882 9.3
R37863 vdd.n37897 vdd.n37896 9.3
R37864 vdd.n37916 vdd.n37915 9.3
R37865 vdd.n37944 vdd.n37943 9.3
R37866 vdd.n37972 vdd.n37971 9.3
R37867 vdd.n38000 vdd.n37999 9.3
R37868 vdd.n38030 vdd.n38029 9.3
R37869 vdd.n38044 vdd.n38043 9.3
R37870 vdd.n38058 vdd.n38057 9.3
R37871 vdd.n38072 vdd.n38071 9.3
R37872 vdd.n38086 vdd.n38085 9.3
R37873 vdd.n38100 vdd.n38099 9.3
R37874 vdd.n38114 vdd.n38113 9.3
R37875 vdd.n38157 vdd.n38156 9.3
R37876 vdd.n38188 vdd.n38187 9.3
R37877 vdd.n37576 vdd.n37575 9.3
R37878 vdd.n35672 vdd.n35671 9.3
R37879 vdd.n37528 vdd.n37527 9.3
R37880 vdd.n32838 vdd.n32837 9.3
R37881 vdd.n32877 vdd.n32876 9.3
R37882 vdd.n37496 vdd.n37495 9.3
R37883 vdd.n32893 vdd.n32892 9.3
R37884 vdd.n32943 vdd.n32942 9.3
R37885 vdd.n37377 vdd.n37376 9.3
R37886 vdd.n37363 vdd.n37362 9.3
R37887 vdd.n37327 vdd.n37326 9.3
R37888 vdd.n32994 vdd.n32993 9.3
R37889 vdd.n33022 vdd.n33021 9.3
R37890 vdd.n37295 vdd.n37294 9.3
R37891 vdd.n33040 vdd.n33039 9.3
R37892 vdd.n37284 vdd.n37283 9.3
R37893 vdd.n33098 vdd.n33097 9.3
R37894 vdd.n37195 vdd.n37194 9.3
R37895 vdd.n37187 vdd.n37186 9.3
R37896 vdd.n37137 vdd.n37136 9.3
R37897 vdd.n33181 vdd.n33180 9.3
R37898 vdd.n37131 vdd.n37130 9.3
R37899 vdd.n33202 vdd.n33201 9.3
R37900 vdd.n37118 vdd.n37117 9.3
R37901 vdd.n33225 vdd.n33224 9.3
R37902 vdd.n37032 vdd.n37031 9.3
R37903 vdd.n37011 vdd.n37010 9.3
R37904 vdd.n36975 vdd.n36974 9.3
R37905 vdd.n36945 vdd.n36944 9.3
R37906 vdd.n36931 vdd.n36930 9.3
R37907 vdd.n36917 vdd.n36916 9.3
R37908 vdd.n36903 vdd.n36902 9.3
R37909 vdd.n36889 vdd.n36888 9.3
R37910 vdd.n36875 vdd.n36874 9.3
R37911 vdd.n36861 vdd.n36860 9.3
R37912 vdd.n36846 vdd.n36845 9.3
R37913 vdd.n36814 vdd.n36813 9.3
R37914 vdd.n36786 vdd.n36785 9.3
R37915 vdd.n36758 vdd.n36757 9.3
R37916 vdd.n36714 vdd.n36713 9.3
R37917 vdd.n36700 vdd.n36699 9.3
R37918 vdd.n36686 vdd.n36685 9.3
R37919 vdd.n36672 vdd.n36671 9.3
R37920 vdd.n36658 vdd.n36657 9.3
R37921 vdd.n36644 vdd.n36643 9.3
R37922 vdd.n36630 vdd.n36629 9.3
R37923 vdd.n36615 vdd.n36614 9.3
R37924 vdd.n36597 vdd.n36596 9.3
R37925 vdd.n36569 vdd.n36568 9.3
R37926 vdd.n36541 vdd.n36540 9.3
R37927 vdd.n36513 vdd.n36512 9.3
R37928 vdd.n36483 vdd.n36482 9.3
R37929 vdd.n36469 vdd.n36468 9.3
R37930 vdd.n36455 vdd.n36454 9.3
R37931 vdd.n36441 vdd.n36440 9.3
R37932 vdd.n36427 vdd.n36426 9.3
R37933 vdd.n36413 vdd.n36412 9.3
R37934 vdd.n36399 vdd.n36398 9.3
R37935 vdd.n36384 vdd.n36383 9.3
R37936 vdd.n36352 vdd.n36351 9.3
R37937 vdd.n36324 vdd.n36323 9.3
R37938 vdd.n36296 vdd.n36295 9.3
R37939 vdd.n36252 vdd.n36251 9.3
R37940 vdd.n36238 vdd.n36237 9.3
R37941 vdd.n36224 vdd.n36223 9.3
R37942 vdd.n36210 vdd.n36209 9.3
R37943 vdd.n36196 vdd.n36195 9.3
R37944 vdd.n36182 vdd.n36181 9.3
R37945 vdd.n36168 vdd.n36167 9.3
R37946 vdd.n36153 vdd.n36152 9.3
R37947 vdd.n36135 vdd.n36134 9.3
R37948 vdd.n36107 vdd.n36106 9.3
R37949 vdd.n36079 vdd.n36078 9.3
R37950 vdd.n36051 vdd.n36050 9.3
R37951 vdd.n36021 vdd.n36020 9.3
R37952 vdd.n36007 vdd.n36006 9.3
R37953 vdd.n35993 vdd.n35992 9.3
R37954 vdd.n35979 vdd.n35978 9.3
R37955 vdd.n35965 vdd.n35964 9.3
R37956 vdd.n35951 vdd.n35950 9.3
R37957 vdd.n35937 vdd.n35936 9.3
R37958 vdd.n35922 vdd.n35921 9.3
R37959 vdd.n35890 vdd.n35889 9.3
R37960 vdd.n35862 vdd.n35861 9.3
R37961 vdd.n35860 vdd.n35859 9.3
R37962 vdd.n35876 vdd.n35875 9.3
R37963 vdd.n35874 vdd.n35873 9.3
R37964 vdd.n35888 vdd.n35887 9.3
R37965 vdd.n35904 vdd.n35903 9.3
R37966 vdd.n35902 vdd.n35901 9.3
R37967 vdd.n35916 vdd.n35915 9.3
R37968 vdd.n35918 vdd.n35917 9.3
R37969 vdd.n35924 vdd.n35923 9.3
R37970 vdd.n35939 vdd.n35938 9.3
R37971 vdd.n35953 vdd.n35952 9.3
R37972 vdd.n35967 vdd.n35966 9.3
R37973 vdd.n35981 vdd.n35980 9.3
R37974 vdd.n35995 vdd.n35994 9.3
R37975 vdd.n36009 vdd.n36008 9.3
R37976 vdd.n36023 vdd.n36022 9.3
R37977 vdd.n36049 vdd.n36048 9.3
R37978 vdd.n36065 vdd.n36064 9.3
R37979 vdd.n36063 vdd.n36062 9.3
R37980 vdd.n36077 vdd.n36076 9.3
R37981 vdd.n36093 vdd.n36092 9.3
R37982 vdd.n36091 vdd.n36090 9.3
R37983 vdd.n36105 vdd.n36104 9.3
R37984 vdd.n36121 vdd.n36120 9.3
R37985 vdd.n36119 vdd.n36118 9.3
R37986 vdd.n36133 vdd.n36132 9.3
R37987 vdd.n36149 vdd.n36148 9.3
R37988 vdd.n36147 vdd.n36146 9.3
R37989 vdd.n36155 vdd.n36154 9.3
R37990 vdd.n36170 vdd.n36169 9.3
R37991 vdd.n36184 vdd.n36183 9.3
R37992 vdd.n36198 vdd.n36197 9.3
R37993 vdd.n36212 vdd.n36211 9.3
R37994 vdd.n36226 vdd.n36225 9.3
R37995 vdd.n36240 vdd.n36239 9.3
R37996 vdd.n36254 vdd.n36253 9.3
R37997 vdd.n36282 vdd.n36281 9.3
R37998 vdd.n36280 vdd.n36279 9.3
R37999 vdd.n36294 vdd.n36293 9.3
R38000 vdd.n36310 vdd.n36309 9.3
R38001 vdd.n36308 vdd.n36307 9.3
R38002 vdd.n36322 vdd.n36321 9.3
R38003 vdd.n36338 vdd.n36337 9.3
R38004 vdd.n36336 vdd.n36335 9.3
R38005 vdd.n36350 vdd.n36349 9.3
R38006 vdd.n36366 vdd.n36365 9.3
R38007 vdd.n36364 vdd.n36363 9.3
R38008 vdd.n36378 vdd.n36377 9.3
R38009 vdd.n36380 vdd.n36379 9.3
R38010 vdd.n36386 vdd.n36385 9.3
R38011 vdd.n36401 vdd.n36400 9.3
R38012 vdd.n36415 vdd.n36414 9.3
R38013 vdd.n36429 vdd.n36428 9.3
R38014 vdd.n36443 vdd.n36442 9.3
R38015 vdd.n36457 vdd.n36456 9.3
R38016 vdd.n36471 vdd.n36470 9.3
R38017 vdd.n36485 vdd.n36484 9.3
R38018 vdd.n36511 vdd.n36510 9.3
R38019 vdd.n36527 vdd.n36526 9.3
R38020 vdd.n36525 vdd.n36524 9.3
R38021 vdd.n36539 vdd.n36538 9.3
R38022 vdd.n36555 vdd.n36554 9.3
R38023 vdd.n36553 vdd.n36552 9.3
R38024 vdd.n36567 vdd.n36566 9.3
R38025 vdd.n36583 vdd.n36582 9.3
R38026 vdd.n36581 vdd.n36580 9.3
R38027 vdd.n36595 vdd.n36594 9.3
R38028 vdd.n36611 vdd.n36610 9.3
R38029 vdd.n36609 vdd.n36608 9.3
R38030 vdd.n36617 vdd.n36616 9.3
R38031 vdd.n36632 vdd.n36631 9.3
R38032 vdd.n36646 vdd.n36645 9.3
R38033 vdd.n36660 vdd.n36659 9.3
R38034 vdd.n36674 vdd.n36673 9.3
R38035 vdd.n36688 vdd.n36687 9.3
R38036 vdd.n36702 vdd.n36701 9.3
R38037 vdd.n36716 vdd.n36715 9.3
R38038 vdd.n36744 vdd.n36743 9.3
R38039 vdd.n36742 vdd.n36741 9.3
R38040 vdd.n36756 vdd.n36755 9.3
R38041 vdd.n36772 vdd.n36771 9.3
R38042 vdd.n36770 vdd.n36769 9.3
R38043 vdd.n36784 vdd.n36783 9.3
R38044 vdd.n36800 vdd.n36799 9.3
R38045 vdd.n36798 vdd.n36797 9.3
R38046 vdd.n36812 vdd.n36811 9.3
R38047 vdd.n36828 vdd.n36827 9.3
R38048 vdd.n36826 vdd.n36825 9.3
R38049 vdd.n36840 vdd.n36839 9.3
R38050 vdd.n36842 vdd.n36841 9.3
R38051 vdd.n36848 vdd.n36847 9.3
R38052 vdd.n36863 vdd.n36862 9.3
R38053 vdd.n36877 vdd.n36876 9.3
R38054 vdd.n36891 vdd.n36890 9.3
R38055 vdd.n36905 vdd.n36904 9.3
R38056 vdd.n36919 vdd.n36918 9.3
R38057 vdd.n36933 vdd.n36932 9.3
R38058 vdd.n36947 vdd.n36946 9.3
R38059 vdd.n36973 vdd.n36972 9.3
R38060 vdd.n36989 vdd.n36988 9.3
R38061 vdd.n37009 vdd.n37008 9.3
R38062 vdd.n37026 vdd.n37025 9.3
R38063 vdd.n37024 vdd.n37023 9.3
R38064 vdd.n37034 vdd.n37033 9.3
R38065 vdd.n37047 vdd.n37046 9.3
R38066 vdd.n33277 vdd.n33276 9.3
R38067 vdd.n33223 vdd.n33222 9.3
R38068 vdd.n37116 vdd.n37115 9.3
R38069 vdd.n33200 vdd.n33199 9.3
R38070 vdd.n37129 vdd.n37128 9.3
R38071 vdd.n35633 vdd.n35632 9.3
R38072 vdd.n33126 vdd.n33125 9.3
R38073 vdd.n33128 vdd.n33127 9.3
R38074 vdd.n37197 vdd.n37196 9.3
R38075 vdd.n37210 vdd.n37209 9.3
R38076 vdd.n33108 vdd.n33107 9.3
R38077 vdd.n33096 vdd.n33095 9.3
R38078 vdd.n37282 vdd.n37281 9.3
R38079 vdd.n33038 vdd.n33037 9.3
R38080 vdd.n33007 vdd.n33006 9.3
R38081 vdd.n37307 vdd.n37306 9.3
R38082 vdd.n32980 vdd.n32979 9.3
R38083 vdd.n37379 vdd.n37378 9.3
R38084 vdd.n37395 vdd.n37394 9.3
R38085 vdd.n37393 vdd.n37392 9.3
R38086 vdd.n32941 vdd.n32940 9.3
R38087 vdd.n37425 vdd.n37424 9.3
R38088 vdd.n37423 vdd.n37422 9.3
R38089 vdd.n32891 vdd.n32890 9.3
R38090 vdd.n32862 vdd.n32861 9.3
R38091 vdd.n37503 vdd.n37502 9.3
R38092 vdd.n32840 vdd.n32839 9.3
R38093 vdd.n32834 vdd.n32833 9.3
R38094 vdd.n38202 vdd.n38201 9.3
R38095 vdd.n38204 vdd.n38203 9.3
R38096 vdd.n38190 vdd.n38189 9.3
R38097 vdd.n38174 vdd.n38173 9.3
R38098 vdd.n38176 vdd.n38175 9.3
R38099 vdd.n38159 vdd.n38158 9.3
R38100 vdd.n38141 vdd.n38140 9.3
R38101 vdd.n38143 vdd.n38142 9.3
R38102 vdd.n38112 vdd.n38111 9.3
R38103 vdd.n38098 vdd.n38097 9.3
R38104 vdd.n38084 vdd.n38083 9.3
R38105 vdd.n38070 vdd.n38069 9.3
R38106 vdd.n38056 vdd.n38055 9.3
R38107 vdd.n38042 vdd.n38041 9.3
R38108 vdd.n38028 vdd.n38027 9.3
R38109 vdd.n38002 vdd.n38001 9.3
R38110 vdd.n37986 vdd.n37985 9.3
R38111 vdd.n37988 vdd.n37987 9.3
R38112 vdd.n37974 vdd.n37973 9.3
R38113 vdd.n37958 vdd.n37957 9.3
R38114 vdd.n37960 vdd.n37959 9.3
R38115 vdd.n37946 vdd.n37945 9.3
R38116 vdd.n37930 vdd.n37929 9.3
R38117 vdd.n37932 vdd.n37931 9.3
R38118 vdd.n37918 vdd.n37917 9.3
R38119 vdd.n37901 vdd.n37900 9.3
R38120 vdd.n37903 vdd.n37902 9.3
R38121 vdd.n37895 vdd.n37894 9.3
R38122 vdd.n37881 vdd.n37880 9.3
R38123 vdd.n37867 vdd.n37866 9.3
R38124 vdd.n37853 vdd.n37852 9.3
R38125 vdd.n37839 vdd.n37838 9.3
R38126 vdd.n37825 vdd.n37824 9.3
R38127 vdd.n37811 vdd.n37810 9.3
R38128 vdd.n37797 vdd.n37796 9.3
R38129 vdd.n37769 vdd.n37768 9.3
R38130 vdd.n37771 vdd.n37770 9.3
R38131 vdd.n37757 vdd.n37756 9.3
R38132 vdd.n37741 vdd.n37740 9.3
R38133 vdd.n37743 vdd.n37742 9.3
R38134 vdd.n37729 vdd.n37728 9.3
R38135 vdd.n37713 vdd.n37712 9.3
R38136 vdd.n37715 vdd.n37714 9.3
R38137 vdd.n37701 vdd.n37700 9.3
R38138 vdd.n37685 vdd.n37684 9.3
R38139 vdd.n37687 vdd.n37686 9.3
R38140 vdd.n37672 vdd.n37671 9.3
R38141 vdd.n37670 vdd.n37669 9.3
R38142 vdd.n37664 vdd.n37663 9.3
R38143 vdd.n37650 vdd.n37649 9.3
R38144 vdd.n37636 vdd.n37635 9.3
R38145 vdd.n37622 vdd.n37621 9.3
R38146 vdd.n37608 vdd.n37607 9.3
R38147 vdd.n28185 vdd.n28184 9.3
R38148 vdd.n28199 vdd.n28198 9.3
R38149 vdd.n28213 vdd.n28212 9.3
R38150 vdd.n28239 vdd.n28238 9.3
R38151 vdd.n28255 vdd.n28254 9.3
R38152 vdd.n28253 vdd.n28252 9.3
R38153 vdd.n28267 vdd.n28266 9.3
R38154 vdd.n28283 vdd.n28282 9.3
R38155 vdd.n28281 vdd.n28280 9.3
R38156 vdd.n28295 vdd.n28294 9.3
R38157 vdd.n28311 vdd.n28310 9.3
R38158 vdd.n28309 vdd.n28308 9.3
R38159 vdd.n28323 vdd.n28322 9.3
R38160 vdd.n28339 vdd.n28338 9.3
R38161 vdd.n28337 vdd.n28336 9.3
R38162 vdd.n28345 vdd.n28344 9.3
R38163 vdd.n28360 vdd.n28359 9.3
R38164 vdd.n28374 vdd.n28373 9.3
R38165 vdd.n28388 vdd.n28387 9.3
R38166 vdd.n28402 vdd.n28401 9.3
R38167 vdd.n28416 vdd.n28415 9.3
R38168 vdd.n28430 vdd.n28429 9.3
R38169 vdd.n28444 vdd.n28443 9.3
R38170 vdd.n28472 vdd.n28471 9.3
R38171 vdd.n28470 vdd.n28469 9.3
R38172 vdd.n28484 vdd.n28483 9.3
R38173 vdd.n28500 vdd.n28499 9.3
R38174 vdd.n28498 vdd.n28497 9.3
R38175 vdd.n28512 vdd.n28511 9.3
R38176 vdd.n28528 vdd.n28527 9.3
R38177 vdd.n28526 vdd.n28525 9.3
R38178 vdd.n28540 vdd.n28539 9.3
R38179 vdd.n28556 vdd.n28555 9.3
R38180 vdd.n28554 vdd.n28553 9.3
R38181 vdd.n28568 vdd.n28567 9.3
R38182 vdd.n28570 vdd.n28569 9.3
R38183 vdd.n28576 vdd.n28575 9.3
R38184 vdd.n28591 vdd.n28590 9.3
R38185 vdd.n28605 vdd.n28604 9.3
R38186 vdd.n28619 vdd.n28618 9.3
R38187 vdd.n28633 vdd.n28632 9.3
R38188 vdd.n28647 vdd.n28646 9.3
R38189 vdd.n28661 vdd.n28660 9.3
R38190 vdd.n28675 vdd.n28674 9.3
R38191 vdd.n28701 vdd.n28700 9.3
R38192 vdd.n28717 vdd.n28716 9.3
R38193 vdd.n28715 vdd.n28714 9.3
R38194 vdd.n28729 vdd.n28728 9.3
R38195 vdd.n28745 vdd.n28744 9.3
R38196 vdd.n28743 vdd.n28742 9.3
R38197 vdd.n28757 vdd.n28756 9.3
R38198 vdd.n28773 vdd.n28772 9.3
R38199 vdd.n28771 vdd.n28770 9.3
R38200 vdd.n28785 vdd.n28784 9.3
R38201 vdd.n28801 vdd.n28800 9.3
R38202 vdd.n28799 vdd.n28798 9.3
R38203 vdd.n28097 vdd.n28096 9.3
R38204 vdd.n27749 vdd.n27748 9.3
R38205 vdd.n28971 vdd.n28970 9.3
R38206 vdd.n27849 vdd.n27848 9.3
R38207 vdd.n27847 vdd.n27846 9.3
R38208 vdd.n27890 vdd.n27889 9.3
R38209 vdd.n27886 vdd.n27885 9.3
R38210 vdd.n29904 vdd.n29876 9.3
R38211 vdd.n29841 vdd.n29840 9.3
R38212 vdd.n29749 vdd.n29748 9.3
R38213 vdd.n29747 vdd.n29746 9.3
R38214 vdd.n29755 vdd.n29754 9.3
R38215 vdd.n29753 vdd.n29752 9.3
R38216 vdd.n30697 vdd.n30696 9.3
R38217 vdd.n29711 vdd.n29710 9.3
R38218 vdd.n30686 vdd.n30685 9.3
R38219 vdd.n30682 vdd.n30681 9.3
R38220 vdd.n30678 vdd.n30677 9.3
R38221 vdd.n30230 vdd.n30229 9.3
R38222 vdd.n28846 vdd.n28844 9.3
R38223 vdd.n28861 vdd.n28859 9.3
R38224 vdd.n28873 vdd.n28871 9.3
R38225 vdd.n28885 vdd.n28883 9.3
R38226 vdd.n28900 vdd.n28898 9.3
R38227 vdd.n28913 vdd.n28911 9.3
R38228 vdd.n28941 vdd.n28939 9.3
R38229 vdd.n28953 vdd.n28951 9.3
R38230 vdd.n28998 vdd.n28996 9.3
R38231 vdd.n29011 vdd.n29009 9.3
R38232 vdd.n28046 vdd.n27771 9.3
R38233 vdd.n28037 vdd.n27775 9.3
R38234 vdd.n28010 vdd.n27829 9.3
R38235 vdd.n28001 vdd.n27856 9.3
R38236 vdd.n27992 vdd.n27861 9.3
R38237 vdd.n27970 vdd.n27866 9.3
R38238 vdd.n27961 vdd.n27871 9.3
R38239 vdd.n27953 vdd.n27897 9.3
R38240 vdd.n29898 vdd.n29896 9.3
R38241 vdd.n29911 vdd.n29909 9.3
R38242 vdd.n29924 vdd.n29922 9.3
R38243 vdd.n29939 vdd.n29931 9.3
R38244 vdd.n29793 vdd.n29791 9.3
R38245 vdd.n29805 vdd.n29803 9.3
R38246 vdd.n29738 vdd.n29704 9.3
R38247 vdd.n29729 vdd.n29708 9.3
R38248 vdd.n30661 vdd.n30659 9.3
R38249 vdd.n30673 vdd.n30671 9.3
R38250 vdd.n30649 vdd.n30177 9.3
R38251 vdd.n30640 vdd.n30181 9.3
R38252 vdd.n30617 vdd.n30256 9.3
R38253 vdd.n30608 vdd.n30260 9.3
R38254 vdd.n30599 vdd.n30279 9.3
R38255 vdd.n30597 vdd.n30281 9.3
R38256 vdd.n30601 vdd.n30278 9.3
R38257 vdd.n30615 vdd.n30258 9.3
R38258 vdd.n30619 vdd.n30255 9.3
R38259 vdd.n30647 vdd.n30178 9.3
R38260 vdd.n30664 vdd.n30662 9.3
R38261 vdd.n29736 vdd.n29705 9.3
R38262 vdd.n29785 vdd.n29696 9.3
R38263 vdd.n29798 vdd.n29795 9.3
R38264 vdd.n29790 vdd.n29788 9.3
R38265 vdd.n29929 vdd.n29926 9.3
R38266 vdd.n29921 vdd.n29919 9.3
R38267 vdd.n29903 vdd.n29900 9.3
R38268 vdd.n29895 vdd.n29893 9.3
R38269 vdd.n27959 vdd.n27872 9.3
R38270 vdd.n27990 vdd.n27862 9.3
R38271 vdd.n28008 vdd.n27830 9.3
R38272 vdd.n28031 vdd.n27778 9.3
R38273 vdd.n28044 vdd.n27773 9.3
R38274 vdd.n28048 vdd.n27770 9.3
R38275 vdd.n29003 vdd.n29000 9.3
R38276 vdd.n28995 vdd.n28993 9.3
R38277 vdd.n28946 vdd.n28943 9.3
R38278 vdd.n28938 vdd.n28936 9.3
R38279 vdd.n28903 vdd.n28901 9.3
R38280 vdd.n28876 vdd.n28874 9.3
R38281 vdd.n28849 vdd.n28847 9.3
R38282 vdd.n28836 vdd.n28834 9.3
R38283 vdd.n28843 vdd.n28840 9.3
R38284 vdd.n28858 vdd.n28855 9.3
R38285 vdd.n28864 vdd.n28862 9.3
R38286 vdd.n28870 vdd.n28867 9.3
R38287 vdd.n28882 vdd.n28879 9.3
R38288 vdd.n28888 vdd.n28886 9.3
R38289 vdd.n28897 vdd.n28894 9.3
R38290 vdd.n28910 vdd.n28907 9.3
R38291 vdd.n28916 vdd.n28914 9.3
R38292 vdd.n28924 vdd.n28921 9.3
R38293 vdd.n28933 vdd.n28930 9.3
R38294 vdd.n28950 vdd.n28948 9.3
R38295 vdd.n28958 vdd.n28955 9.3
R38296 vdd.n29008 vdd.n29006 9.3
R38297 vdd.n29016 vdd.n29013 9.3
R38298 vdd.n28039 vdd.n27774 9.3
R38299 vdd.n28035 vdd.n27777 9.3
R38300 vdd.n28019 vdd.n27826 9.3
R38301 vdd.n28013 vdd.n27828 9.3
R38302 vdd.n28004 vdd.n27855 9.3
R38303 vdd.n27999 vdd.n27857 9.3
R38304 vdd.n27995 vdd.n27860 9.3
R38305 vdd.n27973 vdd.n27865 9.3
R38306 vdd.n27968 vdd.n27867 9.3
R38307 vdd.n27964 vdd.n27870 9.3
R38308 vdd.n27956 vdd.n27896 9.3
R38309 vdd.n27951 vdd.n27898 9.3
R38310 vdd.n27947 vdd.n27900 9.3
R38311 vdd.n27924 vdd.n27920 9.3
R38312 vdd.n29908 vdd.n29906 9.3
R38313 vdd.n29916 vdd.n29913 9.3
R38314 vdd.n29941 vdd.n29930 9.3
R38315 vdd.n29937 vdd.n29933 9.3
R38316 vdd.n29802 vdd.n29800 9.3
R38317 vdd.n29810 vdd.n29807 9.3
R38318 vdd.n29770 vdd.n29701 9.3
R38319 vdd.n29741 vdd.n29703 9.3
R38320 vdd.n29732 vdd.n29707 9.3
R38321 vdd.n29727 vdd.n29709 9.3
R38322 vdd.n30658 vdd.n30655 9.3
R38323 vdd.n30670 vdd.n30667 9.3
R38324 vdd.n30676 vdd.n30674 9.3
R38325 vdd.n30652 vdd.n30176 9.3
R38326 vdd.n30643 vdd.n30180 9.3
R38327 vdd.n30638 vdd.n30182 9.3
R38328 vdd.n30634 vdd.n30211 9.3
R38329 vdd.n30624 vdd.n30226 9.3
R38330 vdd.n30610 vdd.n30259 9.3
R38331 vdd.n30606 vdd.n30262 9.3
R38332 vdd.n30599 vdd.n30598 9.3
R38333 vdd.n30608 vdd.n30607 9.3
R38334 vdd.n30617 vdd.n30616 9.3
R38335 vdd.n30640 vdd.n30639 9.3
R38336 vdd.n30649 vdd.n30648 9.3
R38337 vdd.n30673 vdd.n30672 9.3
R38338 vdd.n30661 vdd.n30660 9.3
R38339 vdd.n29729 vdd.n29728 9.3
R38340 vdd.n29738 vdd.n29737 9.3
R38341 vdd.n29805 vdd.n29804 9.3
R38342 vdd.n29793 vdd.n29792 9.3
R38343 vdd.n29939 vdd.n29938 9.3
R38344 vdd.n29924 vdd.n29923 9.3
R38345 vdd.n29911 vdd.n29910 9.3
R38346 vdd.n29898 vdd.n29897 9.3
R38347 vdd.n27953 vdd.n27952 9.3
R38348 vdd.n27961 vdd.n27960 9.3
R38349 vdd.n27970 vdd.n27969 9.3
R38350 vdd.n27992 vdd.n27991 9.3
R38351 vdd.n28001 vdd.n28000 9.3
R38352 vdd.n28010 vdd.n28009 9.3
R38353 vdd.n28037 vdd.n28036 9.3
R38354 vdd.n28046 vdd.n28045 9.3
R38355 vdd.n29011 vdd.n29010 9.3
R38356 vdd.n28998 vdd.n28997 9.3
R38357 vdd.n28953 vdd.n28952 9.3
R38358 vdd.n28941 vdd.n28940 9.3
R38359 vdd.n28913 vdd.n28912 9.3
R38360 vdd.n28900 vdd.n28899 9.3
R38361 vdd.n28885 vdd.n28884 9.3
R38362 vdd.n28873 vdd.n28872 9.3
R38363 vdd.n28861 vdd.n28860 9.3
R38364 vdd.n28846 vdd.n28845 9.3
R38365 vdd.n28836 vdd.n28835 9.3
R38366 vdd.n28843 vdd.n28842 9.3
R38367 vdd.n28849 vdd.n28848 9.3
R38368 vdd.n28858 vdd.n28857 9.3
R38369 vdd.n28864 vdd.n28863 9.3
R38370 vdd.n28870 vdd.n28869 9.3
R38371 vdd.n28876 vdd.n28875 9.3
R38372 vdd.n28882 vdd.n28881 9.3
R38373 vdd.n28888 vdd.n28887 9.3
R38374 vdd.n28897 vdd.n28896 9.3
R38375 vdd.n28903 vdd.n28902 9.3
R38376 vdd.n28910 vdd.n28909 9.3
R38377 vdd.n28916 vdd.n28915 9.3
R38378 vdd.n28924 vdd.n28923 9.3
R38379 vdd.n28933 vdd.n28932 9.3
R38380 vdd.n28938 vdd.n28937 9.3
R38381 vdd.n28946 vdd.n28945 9.3
R38382 vdd.n28950 vdd.n28949 9.3
R38383 vdd.n28958 vdd.n28957 9.3
R38384 vdd.n28995 vdd.n28994 9.3
R38385 vdd.n29003 vdd.n29002 9.3
R38386 vdd.n29008 vdd.n29007 9.3
R38387 vdd.n29016 vdd.n29015 9.3
R38388 vdd.n28048 vdd.n28047 9.3
R38389 vdd.n28044 vdd.n28043 9.3
R38390 vdd.n28039 vdd.n28038 9.3
R38391 vdd.n28035 vdd.n28034 9.3
R38392 vdd.n28031 vdd.n28030 9.3
R38393 vdd.n28019 vdd.n28018 9.3
R38394 vdd.n28013 vdd.n28012 9.3
R38395 vdd.n28008 vdd.n28007 9.3
R38396 vdd.n28004 vdd.n28003 9.3
R38397 vdd.n27999 vdd.n27998 9.3
R38398 vdd.n27995 vdd.n27994 9.3
R38399 vdd.n27990 vdd.n27989 9.3
R38400 vdd.n27973 vdd.n27972 9.3
R38401 vdd.n27968 vdd.n27967 9.3
R38402 vdd.n27964 vdd.n27963 9.3
R38403 vdd.n27959 vdd.n27958 9.3
R38404 vdd.n27956 vdd.n27955 9.3
R38405 vdd.n27951 vdd.n27950 9.3
R38406 vdd.n27947 vdd.n27946 9.3
R38407 vdd.n27924 vdd.n27923 9.3
R38408 vdd.n29895 vdd.n29894 9.3
R38409 vdd.n29903 vdd.n29902 9.3
R38410 vdd.n29908 vdd.n29907 9.3
R38411 vdd.n29916 vdd.n29915 9.3
R38412 vdd.n29921 vdd.n29920 9.3
R38413 vdd.n29929 vdd.n29928 9.3
R38414 vdd.n29941 vdd.n29940 9.3
R38415 vdd.n29937 vdd.n29936 9.3
R38416 vdd.n29790 vdd.n29789 9.3
R38417 vdd.n29798 vdd.n29797 9.3
R38418 vdd.n29802 vdd.n29801 9.3
R38419 vdd.n29810 vdd.n29809 9.3
R38420 vdd.n29785 vdd.n29784 9.3
R38421 vdd.n29770 vdd.n29769 9.3
R38422 vdd.n29741 vdd.n29740 9.3
R38423 vdd.n29736 vdd.n29735 9.3
R38424 vdd.n29732 vdd.n29731 9.3
R38425 vdd.n29727 vdd.n29726 9.3
R38426 vdd.n30658 vdd.n30657 9.3
R38427 vdd.n30664 vdd.n30663 9.3
R38428 vdd.n30670 vdd.n30669 9.3
R38429 vdd.n30676 vdd.n30675 9.3
R38430 vdd.n30652 vdd.n30651 9.3
R38431 vdd.n30647 vdd.n30646 9.3
R38432 vdd.n30643 vdd.n30642 9.3
R38433 vdd.n30638 vdd.n30637 9.3
R38434 vdd.n30634 vdd.n30633 9.3
R38435 vdd.n30624 vdd.n30623 9.3
R38436 vdd.n30619 vdd.n30618 9.3
R38437 vdd.n30615 vdd.n30614 9.3
R38438 vdd.n30610 vdd.n30609 9.3
R38439 vdd.n30606 vdd.n30605 9.3
R38440 vdd.n30601 vdd.n30600 9.3
R38441 vdd.n30597 vdd.n30596 9.3
R38442 vdd.n28852 vdd.n28851 9.3
R38443 vdd.n28017 vdd.n28016 9.3
R38444 vdd.n27966 vdd.n27965 9.3
R38445 vdd.n29778 vdd.n29777 9.3
R38446 vdd.n30588 vdd.n30288 9.3
R38447 vdd.n30578 vdd.n30305 9.3
R38448 vdd.n30538 vdd.n30317 9.3
R38449 vdd.n30576 vdd.n30309 9.3
R38450 vdd.n30580 vdd.n30303 9.3
R38451 vdd.n30590 vdd.n30286 9.3
R38452 vdd.n30587 vdd.n30290 9.3
R38453 vdd.n30560 vdd.n30312 9.3
R38454 vdd.n30578 vdd.n30304 9.3
R38455 vdd.n30588 vdd.n30287 9.3
R38456 vdd.n30590 vdd.n30589 9.3
R38457 vdd.n30587 vdd.n30586 9.3
R38458 vdd.n30580 vdd.n30579 9.3
R38459 vdd.n30576 vdd.n30307 9.3
R38460 vdd.n30560 vdd.n30559 9.3
R38461 vdd.n30538 vdd.n30537 9.3
R38462 vdd.n30521 vdd.n30520 9.3
R38463 vdd.n30535 vdd.n30534 9.3
R38464 vdd.n30533 vdd.n30532 9.3
R38465 vdd.n30519 vdd.n30518 9.3
R38466 vdd.n27311 vdd.n27310 9.3
R38467 vdd.n27320 vdd.n27319 9.3
R38468 vdd.n27318 vdd.n27317 9.3
R38469 vdd.n27347 vdd.n27346 9.3
R38470 vdd.n27406 vdd.n27405 9.3
R38471 vdd.n27408 vdd.n27407 9.3
R38472 vdd.n27418 vdd.n27417 9.3
R38473 vdd.n27425 vdd.n27424 9.3
R38474 vdd.n27434 vdd.n27433 9.3
R38475 vdd.n27432 vdd.n27431 9.3
R38476 vdd.n27459 vdd.n27458 9.3
R38477 vdd.n27480 vdd.n27479 9.3
R38478 vdd.n27514 vdd.n27513 9.3
R38479 vdd.n27524 vdd.n27523 9.3
R38480 vdd.n27533 vdd.n27532 9.3
R38481 vdd.n27531 vdd.n27530 9.3
R38482 vdd.n27573 vdd.n27572 9.3
R38483 vdd.n27575 vdd.n27574 9.3
R38484 vdd.n27561 vdd.n27560 9.3
R38485 vdd.n27563 vdd.n27562 9.3
R38486 vdd.n27603 vdd.n27602 9.3
R38487 vdd.n27606 vdd.n27605 9.3
R38488 vdd.n27629 vdd.n27628 9.3
R38489 vdd.n27626 vdd.n27625 9.3
R38490 vdd.n27636 vdd.n27635 9.3
R38491 vdd.n27254 vdd.n27253 9.3
R38492 vdd.n25763 vdd.n25762 9.3
R38493 vdd.n25772 vdd.n25771 9.3
R38494 vdd.n25770 vdd.n25769 9.3
R38495 vdd.n25799 vdd.n25798 9.3
R38496 vdd.n25852 vdd.n25851 9.3
R38497 vdd.n25854 vdd.n25853 9.3
R38498 vdd.n25864 vdd.n25863 9.3
R38499 vdd.n25871 vdd.n25870 9.3
R38500 vdd.n25880 vdd.n25879 9.3
R38501 vdd.n25878 vdd.n25877 9.3
R38502 vdd.n25905 vdd.n25904 9.3
R38503 vdd.n25718 vdd.n25717 9.3
R38504 vdd.n26077 vdd.n26066 9.3
R38505 vdd.n25951 vdd.n25950 9.3
R38506 vdd.n25961 vdd.n25960 9.3
R38507 vdd.n25970 vdd.n25969 9.3
R38508 vdd.n25968 vdd.n25967 9.3
R38509 vdd.n25686 vdd.n25685 9.3
R38510 vdd.n25688 vdd.n25687 9.3
R38511 vdd.n25697 vdd.n25696 9.3
R38512 vdd.n25699 vdd.n25698 9.3
R38513 vdd.n26019 vdd.n26018 9.3
R38514 vdd.n26022 vdd.n26021 9.3
R38515 vdd.n26050 vdd.n26049 9.3
R38516 vdd.n26047 vdd.n26046 9.3
R38517 vdd.n26057 vdd.n26056 9.3
R38518 vdd.n25676 vdd.n25675 9.3
R38519 vdd.n25396 vdd.n25389 9.3
R38520 vdd.n25492 vdd.n25491 9.3
R38521 vdd.n25525 vdd.n25524 9.3
R38522 vdd.n25436 vdd.n25435 9.3
R38523 vdd.n25434 vdd.n25433 9.3
R38524 vdd.n25592 vdd.n25591 9.3
R38525 vdd.n25590 vdd.n25589 9.3
R38526 vdd.n25609 vdd.n25608 9.3
R38527 vdd.n25422 vdd.n25421 9.3
R38528 vdd.n25640 vdd.n25638 9.3
R38529 vdd.n25407 vdd.n25406 9.3
R38530 vdd.n25657 vdd.n25656 9.3
R38531 vdd.n25654 vdd.n25653 9.3
R38532 vdd.n3703 vdd.n3701 9.3
R38533 vdd.n3720 vdd.n3718 9.3
R38534 vdd.n4004 vdd.n3733 9.3
R38535 vdd.n3989 vdd.n3750 9.3
R38536 vdd.n3974 vdd.n3765 9.3
R38537 vdd.n3963 vdd.n3771 9.3
R38538 vdd.n3914 vdd.n3912 9.3
R38539 vdd.n3889 vdd.n3801 9.3
R38540 vdd.n3875 vdd.n3810 9.3
R38541 vdd.n3861 vdd.n3824 9.3
R38542 vdd.n3841 vdd.n3839 9.3
R38543 vdd.n2228 vdd.n2226 9.3
R38544 vdd.n2276 vdd.n2274 9.3
R38545 vdd.n2293 vdd.n2291 9.3
R38546 vdd.n2311 vdd.n2309 9.3
R38547 vdd.n2330 vdd.n2328 9.3
R38548 vdd.n2349 vdd.n2347 9.3
R38549 vdd.n2364 vdd.n2362 9.3
R38550 vdd.n2542 vdd.n2426 9.3
R38551 vdd.n2516 vdd.n2434 9.3
R38552 vdd.n2503 vdd.n2441 9.3
R38553 vdd.n2486 vdd.n2452 9.3
R38554 vdd.n2467 vdd.n2465 9.3
R38555 vdd.n2611 vdd.n2609 9.3
R38556 vdd.n1970 vdd.n1968 9.3
R38557 vdd.n1995 vdd.n1983 9.3
R38558 vdd.n2092 vdd.n2090 9.3
R38559 vdd.n2077 vdd.n2075 9.3
R38560 vdd.n1946 vdd.n1941 9.3
R38561 vdd.n1919 vdd.n1207 9.3
R38562 vdd.n1856 vdd.n1230 9.3
R38563 vdd.n1841 vdd.n1244 9.3
R38564 vdd.n1829 vdd.n1253 9.3
R38565 vdd.n1807 vdd.n1257 9.3
R38566 vdd.n1786 vdd.n1264 9.3
R38567 vdd.n1788 vdd.n1262 9.3
R38568 vdd.n1825 vdd.n1822 9.3
R38569 vdd.n1831 vdd.n1252 9.3
R38570 vdd.n1851 vdd.n1232 9.3
R38571 vdd.n1858 vdd.n1229 9.3
R38572 vdd.n1944 vdd.n1942 9.3
R38573 vdd.n2095 vdd.n2093 9.3
R38574 vdd.n1973 vdd.n1971 9.3
R38575 vdd.n2630 vdd.n2628 9.3
R38576 vdd.n2463 vdd.n2460 9.3
R38577 vdd.n2469 vdd.n2458 9.3
R38578 vdd.n2500 vdd.n2448 9.3
R38579 vdd.n2505 vdd.n2440 9.3
R38580 vdd.n2539 vdd.n2430 9.3
R38581 vdd.n2544 vdd.n2425 9.3
R38582 vdd.n2352 vdd.n2350 9.3
R38583 vdd.n2314 vdd.n2312 9.3
R38584 vdd.n2279 vdd.n2277 9.3
R38585 vdd.n2247 vdd.n2245 9.3
R38586 vdd.n3837 vdd.n3834 9.3
R38587 vdd.n3843 vdd.n3832 9.3
R38588 vdd.n3873 vdd.n3870 9.3
R38589 vdd.n3877 vdd.n3809 9.3
R38590 vdd.n3909 vdd.n3799 9.3
R38591 vdd.n3916 vdd.n3797 9.3
R38592 vdd.n3972 vdd.n3766 9.3
R38593 vdd.n4002 vdd.n3734 9.3
R38594 vdd.n3706 vdd.n3704 9.3
R38595 vdd.n3687 vdd.n3685 9.3
R38596 vdd.n3700 vdd.n3697 9.3
R38597 vdd.n3717 vdd.n3714 9.3
R38598 vdd.n4015 vdd.n3721 9.3
R38599 vdd.n4007 vdd.n3732 9.3
R38600 vdd.n3992 vdd.n3749 9.3
R38601 vdd.n3987 vdd.n3751 9.3
R38602 vdd.n3977 vdd.n3764 9.3
R38603 vdd.n3966 vdd.n3770 9.3
R38604 vdd.n3961 vdd.n3772 9.3
R38605 vdd.n3947 vdd.n3777 9.3
R38606 vdd.n3929 vdd.n3793 9.3
R38607 vdd.n3891 vdd.n3800 9.3
R38608 vdd.n3885 vdd.n3882 9.3
R38609 vdd.n3863 vdd.n3823 9.3
R38610 vdd.n3858 vdd.n3831 9.3
R38611 vdd.n2225 vdd.n2223 9.3
R38612 vdd.n2233 vdd.n2230 9.3
R38613 vdd.n2264 vdd.n2262 9.3
R38614 vdd.n2273 vdd.n2270 9.3
R38615 vdd.n2290 vdd.n2287 9.3
R38616 vdd.n2297 vdd.n2295 9.3
R38617 vdd.n2308 vdd.n2305 9.3
R38618 vdd.n2327 vdd.n2324 9.3
R38619 vdd.n2333 vdd.n2331 9.3
R38620 vdd.n2346 vdd.n2343 9.3
R38621 vdd.n2361 vdd.n2358 9.3
R38622 vdd.n2367 vdd.n2365 9.3
R38623 vdd.n2392 vdd.n2389 9.3
R38624 vdd.n2553 vdd.n2412 9.3
R38625 vdd.n2518 vdd.n2433 9.3
R38626 vdd.n2514 vdd.n2438 9.3
R38627 vdd.n2488 vdd.n2451 9.3
R38628 vdd.n2483 vdd.n2456 9.3
R38629 vdd.n2608 vdd.n2606 9.3
R38630 vdd.n2616 vdd.n2613 9.3
R38631 vdd.n2664 vdd.n2662 9.3
R38632 vdd.n1967 vdd.n1964 9.3
R38633 vdd.n1998 vdd.n1982 9.3
R38634 vdd.n1993 vdd.n1984 9.3
R38635 vdd.n2089 vdd.n2086 9.3
R38636 vdd.n2080 vdd.n2074 9.3
R38637 vdd.n1955 vdd.n1953 9.3
R38638 vdd.n1949 vdd.n1940 9.3
R38639 vdd.n1922 vdd.n1206 9.3
R38640 vdd.n1917 vdd.n1208 9.3
R38641 vdd.n1896 vdd.n1212 9.3
R38642 vdd.n1882 vdd.n1875 9.3
R38643 vdd.n1843 vdd.n1243 9.3
R38644 vdd.n1249 vdd.n1246 9.3
R38645 vdd.n1809 vdd.n1256 9.3
R38646 vdd.n1802 vdd.n1259 9.3
R38647 vdd.n3703 vdd.n3702 9.3
R38648 vdd.n3720 vdd.n3719 9.3
R38649 vdd.n4004 vdd.n4003 9.3
R38650 vdd.n3989 vdd.n3988 9.3
R38651 vdd.n3974 vdd.n3973 9.3
R38652 vdd.n3963 vdd.n3962 9.3
R38653 vdd.n3914 vdd.n3913 9.3
R38654 vdd.n3889 vdd.n3888 9.3
R38655 vdd.n3875 vdd.n3874 9.3
R38656 vdd.n3861 vdd.n3860 9.3
R38657 vdd.n3841 vdd.n3840 9.3
R38658 vdd.n2228 vdd.n2227 9.3
R38659 vdd.n2276 vdd.n2275 9.3
R38660 vdd.n2293 vdd.n2292 9.3
R38661 vdd.n2311 vdd.n2310 9.3
R38662 vdd.n2330 vdd.n2329 9.3
R38663 vdd.n2349 vdd.n2348 9.3
R38664 vdd.n2364 vdd.n2363 9.3
R38665 vdd.n2542 vdd.n2541 9.3
R38666 vdd.n2516 vdd.n2515 9.3
R38667 vdd.n2503 vdd.n2502 9.3
R38668 vdd.n2486 vdd.n2485 9.3
R38669 vdd.n2467 vdd.n2466 9.3
R38670 vdd.n2611 vdd.n2610 9.3
R38671 vdd.n1970 vdd.n1969 9.3
R38672 vdd.n1995 vdd.n1994 9.3
R38673 vdd.n2092 vdd.n2091 9.3
R38674 vdd.n2077 vdd.n2076 9.3
R38675 vdd.n1946 vdd.n1945 9.3
R38676 vdd.n1919 vdd.n1918 9.3
R38677 vdd.n1856 vdd.n1855 9.3
R38678 vdd.n1841 vdd.n1840 9.3
R38679 vdd.n1829 vdd.n1828 9.3
R38680 vdd.n1807 vdd.n1806 9.3
R38681 vdd.n1786 vdd.n1263 9.3
R38682 vdd.n1788 vdd.n1787 9.3
R38683 vdd.n1825 vdd.n1824 9.3
R38684 vdd.n1831 vdd.n1830 9.3
R38685 vdd.n1851 vdd.n1850 9.3
R38686 vdd.n1858 vdd.n1857 9.3
R38687 vdd.n1944 vdd.n1943 9.3
R38688 vdd.n2095 vdd.n2094 9.3
R38689 vdd.n1973 vdd.n1972 9.3
R38690 vdd.n2630 vdd.n2629 9.3
R38691 vdd.n2463 vdd.n2462 9.3
R38692 vdd.n2469 vdd.n2468 9.3
R38693 vdd.n2500 vdd.n2499 9.3
R38694 vdd.n2505 vdd.n2504 9.3
R38695 vdd.n2539 vdd.n2538 9.3
R38696 vdd.n2544 vdd.n2543 9.3
R38697 vdd.n2352 vdd.n2351 9.3
R38698 vdd.n2314 vdd.n2313 9.3
R38699 vdd.n2279 vdd.n2278 9.3
R38700 vdd.n2247 vdd.n2246 9.3
R38701 vdd.n3837 vdd.n3836 9.3
R38702 vdd.n3843 vdd.n3842 9.3
R38703 vdd.n3873 vdd.n3872 9.3
R38704 vdd.n3877 vdd.n3876 9.3
R38705 vdd.n3909 vdd.n3908 9.3
R38706 vdd.n3916 vdd.n3915 9.3
R38707 vdd.n3972 vdd.n3971 9.3
R38708 vdd.n4002 vdd.n4001 9.3
R38709 vdd.n3706 vdd.n3705 9.3
R38710 vdd.n3687 vdd.n3686 9.3
R38711 vdd.n3700 vdd.n3699 9.3
R38712 vdd.n3717 vdd.n3716 9.3
R38713 vdd.n4015 vdd.n4014 9.3
R38714 vdd.n4007 vdd.n4006 9.3
R38715 vdd.n3992 vdd.n3991 9.3
R38716 vdd.n3987 vdd.n3986 9.3
R38717 vdd.n3977 vdd.n3976 9.3
R38718 vdd.n3966 vdd.n3965 9.3
R38719 vdd.n3961 vdd.n3960 9.3
R38720 vdd.n3947 vdd.n3946 9.3
R38721 vdd.n3929 vdd.n3928 9.3
R38722 vdd.n3891 vdd.n3890 9.3
R38723 vdd.n3885 vdd.n3884 9.3
R38724 vdd.n3863 vdd.n3862 9.3
R38725 vdd.n3858 vdd.n3857 9.3
R38726 vdd.n2225 vdd.n2224 9.3
R38727 vdd.n2233 vdd.n2232 9.3
R38728 vdd.n2264 vdd.n2263 9.3
R38729 vdd.n2273 vdd.n2272 9.3
R38730 vdd.n2290 vdd.n2289 9.3
R38731 vdd.n2297 vdd.n2296 9.3
R38732 vdd.n2308 vdd.n2307 9.3
R38733 vdd.n2327 vdd.n2326 9.3
R38734 vdd.n2333 vdd.n2332 9.3
R38735 vdd.n2346 vdd.n2345 9.3
R38736 vdd.n2361 vdd.n2360 9.3
R38737 vdd.n2367 vdd.n2366 9.3
R38738 vdd.n2392 vdd.n2391 9.3
R38739 vdd.n2553 vdd.n2552 9.3
R38740 vdd.n2518 vdd.n2517 9.3
R38741 vdd.n2514 vdd.n2513 9.3
R38742 vdd.n2488 vdd.n2487 9.3
R38743 vdd.n2483 vdd.n2482 9.3
R38744 vdd.n2608 vdd.n2607 9.3
R38745 vdd.n2616 vdd.n2615 9.3
R38746 vdd.n2664 vdd.n2663 9.3
R38747 vdd.n1967 vdd.n1966 9.3
R38748 vdd.n1998 vdd.n1997 9.3
R38749 vdd.n1993 vdd.n1992 9.3
R38750 vdd.n2089 vdd.n2088 9.3
R38751 vdd.n2080 vdd.n2079 9.3
R38752 vdd.n1955 vdd.n1954 9.3
R38753 vdd.n1949 vdd.n1948 9.3
R38754 vdd.n1922 vdd.n1921 9.3
R38755 vdd.n1917 vdd.n1916 9.3
R38756 vdd.n1896 vdd.n1895 9.3
R38757 vdd.n1882 vdd.n1228 9.3
R38758 vdd.n1843 vdd.n1842 9.3
R38759 vdd.n1249 vdd.n1248 9.3
R38760 vdd.n1809 vdd.n1808 9.3
R38761 vdd.n1802 vdd.n1801 9.3
R38762 vdd.n1288 vdd.n1287 9.3
R38763 vdd.n1763 vdd.n1762 9.3
R38764 vdd.n1752 vdd.n1751 9.3
R38765 vdd.n1728 vdd.n1727 9.3
R38766 vdd.n1717 vdd.n1716 9.3
R38767 vdd.n1706 vdd.n1705 9.3
R38768 vdd.n1695 vdd.n1694 9.3
R38769 vdd.n1684 vdd.n1683 9.3
R38770 vdd.n1673 vdd.n1672 9.3
R38771 vdd.n1662 vdd.n1661 9.3
R38772 vdd.n1643 vdd.n1642 9.3
R38773 vdd.n1632 vdd.n1631 9.3
R38774 vdd.n1621 vdd.n1620 9.3
R38775 vdd.n1610 vdd.n1609 9.3
R38776 vdd.n1599 vdd.n1598 9.3
R38777 vdd.n1588 vdd.n1587 9.3
R38778 vdd.n1577 vdd.n1576 9.3
R38779 vdd.n1566 vdd.n1565 9.3
R38780 vdd.n1558 vdd.n1557 9.3
R38781 vdd.n1547 vdd.n1546 9.3
R38782 vdd.n1536 vdd.n1535 9.3
R38783 vdd.n1525 vdd.n1524 9.3
R38784 vdd.n1514 vdd.n1513 9.3
R38785 vdd.n1503 vdd.n1502 9.3
R38786 vdd.n1492 vdd.n1491 9.3
R38787 vdd.n1481 vdd.n1480 9.3
R38788 vdd.n1462 vdd.n1461 9.3
R38789 vdd.n1451 vdd.n1450 9.3
R38790 vdd.n1440 vdd.n1439 9.3
R38791 vdd.n1429 vdd.n1428 9.3
R38792 vdd.n1418 vdd.n1417 9.3
R38793 vdd.n1407 vdd.n1406 9.3
R38794 vdd.n1396 vdd.n1395 9.3
R38795 vdd.n1385 vdd.n1384 9.3
R38796 vdd.n1377 vdd.n1376 9.3
R38797 vdd.n1366 vdd.n1365 9.3
R38798 vdd.n1355 vdd.n1354 9.3
R38799 vdd.n1344 vdd.n1343 9.3
R38800 vdd.n1333 vdd.n1332 9.3
R38801 vdd.n1322 vdd.n1321 9.3
R38802 vdd.n1311 vdd.n1310 9.3
R38803 vdd.n1300 vdd.n1299 9.3
R38804 vdd.n26766 vdd.n26765 9.3
R38805 vdd.n26777 vdd.n26776 9.3
R38806 vdd.n26788 vdd.n26787 9.3
R38807 vdd.n26799 vdd.n26798 9.3
R38808 vdd.n26810 vdd.n26809 9.3
R38809 vdd.n26821 vdd.n26820 9.3
R38810 vdd.n26832 vdd.n26831 9.3
R38811 vdd.n26843 vdd.n26842 9.3
R38812 vdd.n26851 vdd.n26850 9.3
R38813 vdd.n26862 vdd.n26861 9.3
R38814 vdd.n26873 vdd.n26872 9.3
R38815 vdd.n26884 vdd.n26883 9.3
R38816 vdd.n26895 vdd.n26894 9.3
R38817 vdd.n26906 vdd.n26905 9.3
R38818 vdd.n26917 vdd.n26916 9.3
R38819 vdd.n26928 vdd.n26927 9.3
R38820 vdd.n26947 vdd.n26946 9.3
R38821 vdd.n26958 vdd.n26957 9.3
R38822 vdd.n26969 vdd.n26968 9.3
R38823 vdd.n26980 vdd.n26979 9.3
R38824 vdd.n26991 vdd.n26990 9.3
R38825 vdd.n27002 vdd.n27001 9.3
R38826 vdd.n27013 vdd.n27012 9.3
R38827 vdd.n27024 vdd.n27023 9.3
R38828 vdd.n27032 vdd.n27031 9.3
R38829 vdd.n27043 vdd.n27042 9.3
R38830 vdd.n27054 vdd.n27053 9.3
R38831 vdd.n27065 vdd.n27064 9.3
R38832 vdd.n27076 vdd.n27075 9.3
R38833 vdd.n27087 vdd.n27086 9.3
R38834 vdd.n27098 vdd.n27097 9.3
R38835 vdd.n27109 vdd.n27108 9.3
R38836 vdd.n27128 vdd.n27127 9.3
R38837 vdd.n27139 vdd.n27138 9.3
R38838 vdd.n27150 vdd.n27149 9.3
R38839 vdd.n27161 vdd.n27160 9.3
R38840 vdd.n27172 vdd.n27171 9.3
R38841 vdd.n27183 vdd.n27182 9.3
R38842 vdd.n27194 vdd.n27193 9.3
R38843 vdd.n27205 vdd.n27204 9.3
R38844 vdd.n26757 vdd.n26756 9.3
R38845 vdd.n1286 vdd.n1275 9.3
R38846 vdd.n1761 vdd.n1760 9.3
R38847 vdd.n1750 vdd.n1749 9.3
R38848 vdd.n1730 vdd.n1729 9.3
R38849 vdd.n1719 vdd.n1718 9.3
R38850 vdd.n1708 vdd.n1707 9.3
R38851 vdd.n1697 vdd.n1696 9.3
R38852 vdd.n1686 vdd.n1685 9.3
R38853 vdd.n1675 vdd.n1674 9.3
R38854 vdd.n1664 vdd.n1663 9.3
R38855 vdd.n1641 vdd.n1640 9.3
R38856 vdd.n1630 vdd.n1629 9.3
R38857 vdd.n1619 vdd.n1618 9.3
R38858 vdd.n1608 vdd.n1607 9.3
R38859 vdd.n1597 vdd.n1596 9.3
R38860 vdd.n1586 vdd.n1585 9.3
R38861 vdd.n1575 vdd.n1574 9.3
R38862 vdd.n1564 vdd.n1563 9.3
R38863 vdd.n1560 vdd.n1559 9.3
R38864 vdd.n1549 vdd.n1548 9.3
R38865 vdd.n1538 vdd.n1537 9.3
R38866 vdd.n1527 vdd.n1526 9.3
R38867 vdd.n1516 vdd.n1515 9.3
R38868 vdd.n1505 vdd.n1504 9.3
R38869 vdd.n1494 vdd.n1493 9.3
R38870 vdd.n1483 vdd.n1482 9.3
R38871 vdd.n1460 vdd.n1459 9.3
R38872 vdd.n1449 vdd.n1448 9.3
R38873 vdd.n1438 vdd.n1437 9.3
R38874 vdd.n1427 vdd.n1426 9.3
R38875 vdd.n1416 vdd.n1415 9.3
R38876 vdd.n1405 vdd.n1404 9.3
R38877 vdd.n1394 vdd.n1393 9.3
R38878 vdd.n1383 vdd.n1382 9.3
R38879 vdd.n1379 vdd.n1378 9.3
R38880 vdd.n1368 vdd.n1367 9.3
R38881 vdd.n1357 vdd.n1356 9.3
R38882 vdd.n1346 vdd.n1345 9.3
R38883 vdd.n1335 vdd.n1334 9.3
R38884 vdd.n1324 vdd.n1323 9.3
R38885 vdd.n1313 vdd.n1312 9.3
R38886 vdd.n1302 vdd.n1301 9.3
R38887 vdd.n26768 vdd.n26767 9.3
R38888 vdd.n26779 vdd.n26778 9.3
R38889 vdd.n26790 vdd.n26789 9.3
R38890 vdd.n26801 vdd.n26800 9.3
R38891 vdd.n26812 vdd.n26811 9.3
R38892 vdd.n26823 vdd.n26822 9.3
R38893 vdd.n26834 vdd.n26833 9.3
R38894 vdd.n26845 vdd.n26844 9.3
R38895 vdd.n26849 vdd.n26848 9.3
R38896 vdd.n26860 vdd.n26859 9.3
R38897 vdd.n26871 vdd.n26870 9.3
R38898 vdd.n26882 vdd.n26881 9.3
R38899 vdd.n26893 vdd.n26892 9.3
R38900 vdd.n26904 vdd.n26903 9.3
R38901 vdd.n26915 vdd.n26914 9.3
R38902 vdd.n26926 vdd.n26925 9.3
R38903 vdd.n26949 vdd.n26948 9.3
R38904 vdd.n26960 vdd.n26959 9.3
R38905 vdd.n26971 vdd.n26970 9.3
R38906 vdd.n26982 vdd.n26981 9.3
R38907 vdd.n26993 vdd.n26992 9.3
R38908 vdd.n27004 vdd.n27003 9.3
R38909 vdd.n27015 vdd.n27014 9.3
R38910 vdd.n27026 vdd.n27025 9.3
R38911 vdd.n27030 vdd.n27029 9.3
R38912 vdd.n27041 vdd.n27040 9.3
R38913 vdd.n27052 vdd.n27051 9.3
R38914 vdd.n27063 vdd.n27062 9.3
R38915 vdd.n27074 vdd.n27073 9.3
R38916 vdd.n27085 vdd.n27084 9.3
R38917 vdd.n27096 vdd.n27095 9.3
R38918 vdd.n27107 vdd.n27106 9.3
R38919 vdd.n27130 vdd.n27129 9.3
R38920 vdd.n27141 vdd.n27140 9.3
R38921 vdd.n27152 vdd.n27151 9.3
R38922 vdd.n27163 vdd.n27162 9.3
R38923 vdd.n27174 vdd.n27173 9.3
R38924 vdd.n27185 vdd.n27184 9.3
R38925 vdd.n27196 vdd.n27195 9.3
R38926 vdd.n27207 vdd.n27206 9.3
R38927 vdd.n26755 vdd.n26739 9.3
R38928 vdd.n26731 vdd.n26730 9.3
R38929 vdd.n1790 vdd.n1789 9.3
R38930 vdd.n1848 vdd.n1847 9.3
R38931 vdd.n1872 vdd.n1871 9.3
R38932 vdd.n2063 vdd.n2062 9.3
R38933 vdd.n2669 vdd.n2668 9.3
R38934 vdd.n2658 vdd.n2657 9.3
R38935 vdd.n2642 vdd.n2641 9.3
R38936 vdd.n2644 vdd.n2643 9.3
R38937 vdd.n2627 vdd.n2626 9.3
R38938 vdd.n2605 vdd.n2604 9.3
R38939 vdd.n2471 vdd.n2470 9.3
R38940 vdd.n2490 vdd.n2489 9.3
R38941 vdd.n2121 vdd.n2120 9.3
R38942 vdd.n2168 vdd.n2167 9.3
R38943 vdd.n2186 vdd.n2185 9.3
R38944 vdd.n2244 vdd.n2243 9.3
R38945 vdd.n2222 vdd.n2221 9.3
R38946 vdd.n3845 vdd.n3844 9.3
R38947 vdd.n3906 vdd.n3905 9.3
R38948 vdd.n3924 vdd.n3923 9.3
R38949 vdd.n3926 vdd.n3925 9.3
R38950 vdd.n3942 vdd.n3941 9.3
R38951 vdd.n3958 vdd.n3957 9.3
R38952 vdd.n3753 vdd.n3752 9.3
R38953 vdd.n3738 vdd.n3737 9.3
R38954 vdd.n2694 vdd.n2693 9.3
R38955 vdd.n2710 vdd.n2709 9.3
R38956 vdd.n2752 vdd.n2751 9.3
R38957 vdd.n2763 vdd.n2762 9.3
R38958 vdd.n2774 vdd.n2773 9.3
R38959 vdd.n2785 vdd.n2784 9.3
R38960 vdd.n2796 vdd.n2795 9.3
R38961 vdd.n2804 vdd.n2803 9.3
R38962 vdd.n2815 vdd.n2814 9.3
R38963 vdd.n2826 vdd.n2825 9.3
R38964 vdd.n2837 vdd.n2836 9.3
R38965 vdd.n2848 vdd.n2847 9.3
R38966 vdd.n2859 vdd.n2858 9.3
R38967 vdd.n2870 vdd.n2869 9.3
R38968 vdd.n2881 vdd.n2880 9.3
R38969 vdd.n2900 vdd.n2899 9.3
R38970 vdd.n2911 vdd.n2910 9.3
R38971 vdd.n2922 vdd.n2921 9.3
R38972 vdd.n2933 vdd.n2932 9.3
R38973 vdd.n2944 vdd.n2943 9.3
R38974 vdd.n2955 vdd.n2954 9.3
R38975 vdd.n2966 vdd.n2965 9.3
R38976 vdd.n2977 vdd.n2976 9.3
R38977 vdd.n2985 vdd.n2984 9.3
R38978 vdd.n2996 vdd.n2995 9.3
R38979 vdd.n3007 vdd.n3006 9.3
R38980 vdd.n3018 vdd.n3017 9.3
R38981 vdd.n3029 vdd.n3028 9.3
R38982 vdd.n3040 vdd.n3039 9.3
R38983 vdd.n3051 vdd.n3050 9.3
R38984 vdd.n3062 vdd.n3061 9.3
R38985 vdd.n3081 vdd.n3080 9.3
R38986 vdd.n3092 vdd.n3091 9.3
R38987 vdd.n3103 vdd.n3102 9.3
R38988 vdd.n3114 vdd.n3113 9.3
R38989 vdd.n3125 vdd.n3124 9.3
R38990 vdd.n3136 vdd.n3135 9.3
R38991 vdd.n3147 vdd.n3146 9.3
R38992 vdd.n3158 vdd.n3157 9.3
R38993 vdd.n3166 vdd.n3165 9.3
R38994 vdd.n3177 vdd.n3176 9.3
R38995 vdd.n3188 vdd.n3187 9.3
R38996 vdd.n3199 vdd.n3198 9.3
R38997 vdd.n3210 vdd.n3209 9.3
R38998 vdd.n3221 vdd.n3220 9.3
R38999 vdd.n3232 vdd.n3231 9.3
R39000 vdd.n3243 vdd.n3242 9.3
R39001 vdd.n3262 vdd.n3261 9.3
R39002 vdd.n3273 vdd.n3272 9.3
R39003 vdd.n3284 vdd.n3283 9.3
R39004 vdd.n3295 vdd.n3294 9.3
R39005 vdd.n3306 vdd.n3305 9.3
R39006 vdd.n3317 vdd.n3316 9.3
R39007 vdd.n3328 vdd.n3327 9.3
R39008 vdd.n3339 vdd.n3338 9.3
R39009 vdd.n3347 vdd.n3346 9.3
R39010 vdd.n3358 vdd.n3357 9.3
R39011 vdd.n3369 vdd.n3368 9.3
R39012 vdd.n3380 vdd.n3379 9.3
R39013 vdd.n3391 vdd.n3390 9.3
R39014 vdd.n3402 vdd.n3401 9.3
R39015 vdd.n3413 vdd.n3412 9.3
R39016 vdd.n3424 vdd.n3423 9.3
R39017 vdd.n3443 vdd.n3442 9.3
R39018 vdd.n3454 vdd.n3453 9.3
R39019 vdd.n3465 vdd.n3464 9.3
R39020 vdd.n3476 vdd.n3475 9.3
R39021 vdd.n3487 vdd.n3486 9.3
R39022 vdd.n3498 vdd.n3497 9.3
R39023 vdd.n3509 vdd.n3508 9.3
R39024 vdd.n3520 vdd.n3519 9.3
R39025 vdd.n3528 vdd.n3527 9.3
R39026 vdd.n3539 vdd.n3538 9.3
R39027 vdd.n3550 vdd.n3549 9.3
R39028 vdd.n3561 vdd.n3560 9.3
R39029 vdd.n3572 vdd.n3571 9.3
R39030 vdd.n3583 vdd.n3582 9.3
R39031 vdd.n3594 vdd.n3593 9.3
R39032 vdd.n3605 vdd.n3604 9.3
R39033 vdd.n3624 vdd.n3623 9.3
R39034 vdd.n2754 vdd.n2753 9.3
R39035 vdd.n2765 vdd.n2764 9.3
R39036 vdd.n2776 vdd.n2775 9.3
R39037 vdd.n2787 vdd.n2786 9.3
R39038 vdd.n2798 vdd.n2797 9.3
R39039 vdd.n2802 vdd.n2801 9.3
R39040 vdd.n2813 vdd.n2812 9.3
R39041 vdd.n2824 vdd.n2823 9.3
R39042 vdd.n2835 vdd.n2834 9.3
R39043 vdd.n2846 vdd.n2845 9.3
R39044 vdd.n2857 vdd.n2856 9.3
R39045 vdd.n2868 vdd.n2867 9.3
R39046 vdd.n2879 vdd.n2878 9.3
R39047 vdd.n2902 vdd.n2901 9.3
R39048 vdd.n2913 vdd.n2912 9.3
R39049 vdd.n2924 vdd.n2923 9.3
R39050 vdd.n2935 vdd.n2934 9.3
R39051 vdd.n2946 vdd.n2945 9.3
R39052 vdd.n2957 vdd.n2956 9.3
R39053 vdd.n2968 vdd.n2967 9.3
R39054 vdd.n2979 vdd.n2978 9.3
R39055 vdd.n2983 vdd.n2982 9.3
R39056 vdd.n2994 vdd.n2993 9.3
R39057 vdd.n3005 vdd.n3004 9.3
R39058 vdd.n3016 vdd.n3015 9.3
R39059 vdd.n3027 vdd.n3026 9.3
R39060 vdd.n3038 vdd.n3037 9.3
R39061 vdd.n3049 vdd.n3048 9.3
R39062 vdd.n3060 vdd.n3059 9.3
R39063 vdd.n3083 vdd.n3082 9.3
R39064 vdd.n3094 vdd.n3093 9.3
R39065 vdd.n3105 vdd.n3104 9.3
R39066 vdd.n3116 vdd.n3115 9.3
R39067 vdd.n3127 vdd.n3126 9.3
R39068 vdd.n3138 vdd.n3137 9.3
R39069 vdd.n3149 vdd.n3148 9.3
R39070 vdd.n3160 vdd.n3159 9.3
R39071 vdd.n3164 vdd.n3163 9.3
R39072 vdd.n3175 vdd.n3174 9.3
R39073 vdd.n3186 vdd.n3185 9.3
R39074 vdd.n3197 vdd.n3196 9.3
R39075 vdd.n3208 vdd.n3207 9.3
R39076 vdd.n3219 vdd.n3218 9.3
R39077 vdd.n3230 vdd.n3229 9.3
R39078 vdd.n3241 vdd.n3240 9.3
R39079 vdd.n3264 vdd.n3263 9.3
R39080 vdd.n3275 vdd.n3274 9.3
R39081 vdd.n3286 vdd.n3285 9.3
R39082 vdd.n3297 vdd.n3296 9.3
R39083 vdd.n3308 vdd.n3307 9.3
R39084 vdd.n3319 vdd.n3318 9.3
R39085 vdd.n3330 vdd.n3329 9.3
R39086 vdd.n3341 vdd.n3340 9.3
R39087 vdd.n3345 vdd.n3344 9.3
R39088 vdd.n3356 vdd.n3355 9.3
R39089 vdd.n3367 vdd.n3366 9.3
R39090 vdd.n3378 vdd.n3377 9.3
R39091 vdd.n3389 vdd.n3388 9.3
R39092 vdd.n3400 vdd.n3399 9.3
R39093 vdd.n3411 vdd.n3410 9.3
R39094 vdd.n3422 vdd.n3421 9.3
R39095 vdd.n3445 vdd.n3444 9.3
R39096 vdd.n3456 vdd.n3455 9.3
R39097 vdd.n3467 vdd.n3466 9.3
R39098 vdd.n3478 vdd.n3477 9.3
R39099 vdd.n3489 vdd.n3488 9.3
R39100 vdd.n3500 vdd.n3499 9.3
R39101 vdd.n3511 vdd.n3510 9.3
R39102 vdd.n3522 vdd.n3521 9.3
R39103 vdd.n3526 vdd.n3525 9.3
R39104 vdd.n3537 vdd.n3536 9.3
R39105 vdd.n3548 vdd.n3547 9.3
R39106 vdd.n3559 vdd.n3558 9.3
R39107 vdd.n3570 vdd.n3569 9.3
R39108 vdd.n3581 vdd.n3580 9.3
R39109 vdd.n3592 vdd.n3591 9.3
R39110 vdd.n3603 vdd.n3602 9.3
R39111 vdd.n3626 vdd.n3625 9.3
R39112 vdd.n30300 vdd.n30299 9.3
R39113 vdd.n30299 vdd.n30298 9.3
R39114 vdd.n27768 vdd.n27767 9.3
R39115 vdd.n27767 vdd.n27766 9.3
R39116 vdd.n28566 vdd.n28565 9.3
R39117 vdd.n28565 vdd.n28564 9.3
R39118 vdd.n28564 vdd.n28563 9.3
R39119 vdd.n37683 vdd.n37682 9.3
R39120 vdd.n37682 vdd.n37681 9.3
R39121 vdd.n37681 vdd.n37680 9.3
R39122 vdd.n38125 vdd.n38124 9.3
R39123 vdd.n38124 vdd.n38123 9.3
R39124 vdd.n33075 vdd.n33074 9.3
R39125 vdd.n33074 vdd.n33073 9.3
R39126 vdd.n33073 vdd.n33072 9.3
R39127 vdd.n36838 vdd.n36837 9.3
R39128 vdd.n36837 vdd.n36836 9.3
R39129 vdd.n36836 vdd.n36835 9.3
R39130 vdd.n36376 vdd.n36375 9.3
R39131 vdd.n36375 vdd.n36374 9.3
R39132 vdd.n36374 vdd.n36373 9.3
R39133 vdd.n35914 vdd.n35913 9.3
R39134 vdd.n35913 vdd.n35912 9.3
R39135 vdd.n35912 vdd.n35911 9.3
R39136 vdd.n35846 vdd.n35845 9.3
R39137 vdd.n35845 vdd.n35844 9.3
R39138 vdd.n35858 vdd.n35857 9.3
R39139 vdd.n35857 vdd.n35856 9.3
R39140 vdd.n35856 vdd.n35855 9.3
R39141 vdd.n35872 vdd.n35871 9.3
R39142 vdd.n35871 vdd.n35870 9.3
R39143 vdd.n35870 vdd.n35869 9.3
R39144 vdd.n35886 vdd.n35885 9.3
R39145 vdd.n35885 vdd.n35884 9.3
R39146 vdd.n35884 vdd.n35883 9.3
R39147 vdd.n35900 vdd.n35899 9.3
R39148 vdd.n35899 vdd.n35898 9.3
R39149 vdd.n35898 vdd.n35897 9.3
R39150 vdd.n35935 vdd.n35934 9.3
R39151 vdd.n35934 vdd.n35933 9.3
R39152 vdd.n35933 vdd.n35932 9.3
R39153 vdd.n35949 vdd.n35948 9.3
R39154 vdd.n35948 vdd.n35947 9.3
R39155 vdd.n35947 vdd.n35946 9.3
R39156 vdd.n35963 vdd.n35962 9.3
R39157 vdd.n35962 vdd.n35961 9.3
R39158 vdd.n35961 vdd.n35960 9.3
R39159 vdd.n35977 vdd.n35976 9.3
R39160 vdd.n35976 vdd.n35975 9.3
R39161 vdd.n35975 vdd.n35974 9.3
R39162 vdd.n35991 vdd.n35990 9.3
R39163 vdd.n35990 vdd.n35989 9.3
R39164 vdd.n35989 vdd.n35988 9.3
R39165 vdd.n36005 vdd.n36004 9.3
R39166 vdd.n36004 vdd.n36003 9.3
R39167 vdd.n36003 vdd.n36002 9.3
R39168 vdd.n36019 vdd.n36018 9.3
R39169 vdd.n36018 vdd.n36017 9.3
R39170 vdd.n36017 vdd.n36016 9.3
R39171 vdd.n36033 vdd.n36032 9.3
R39172 vdd.n36032 vdd.n36031 9.3
R39173 vdd.n36031 vdd.n36030 9.3
R39174 vdd.n36047 vdd.n36046 9.3
R39175 vdd.n36046 vdd.n36045 9.3
R39176 vdd.n36045 vdd.n36044 9.3
R39177 vdd.n36061 vdd.n36060 9.3
R39178 vdd.n36060 vdd.n36059 9.3
R39179 vdd.n36059 vdd.n36058 9.3
R39180 vdd.n36075 vdd.n36074 9.3
R39181 vdd.n36074 vdd.n36073 9.3
R39182 vdd.n36073 vdd.n36072 9.3
R39183 vdd.n36089 vdd.n36088 9.3
R39184 vdd.n36088 vdd.n36087 9.3
R39185 vdd.n36087 vdd.n36086 9.3
R39186 vdd.n36103 vdd.n36102 9.3
R39187 vdd.n36102 vdd.n36101 9.3
R39188 vdd.n36101 vdd.n36100 9.3
R39189 vdd.n36117 vdd.n36116 9.3
R39190 vdd.n36116 vdd.n36115 9.3
R39191 vdd.n36115 vdd.n36114 9.3
R39192 vdd.n36131 vdd.n36130 9.3
R39193 vdd.n36130 vdd.n36129 9.3
R39194 vdd.n36129 vdd.n36128 9.3
R39195 vdd.n36145 vdd.n36144 9.3
R39196 vdd.n36144 vdd.n36143 9.3
R39197 vdd.n36143 vdd.n36142 9.3
R39198 vdd.n36166 vdd.n36165 9.3
R39199 vdd.n36165 vdd.n36164 9.3
R39200 vdd.n36164 vdd.n36163 9.3
R39201 vdd.n36180 vdd.n36179 9.3
R39202 vdd.n36179 vdd.n36178 9.3
R39203 vdd.n36178 vdd.n36177 9.3
R39204 vdd.n36194 vdd.n36193 9.3
R39205 vdd.n36193 vdd.n36192 9.3
R39206 vdd.n36192 vdd.n36191 9.3
R39207 vdd.n36208 vdd.n36207 9.3
R39208 vdd.n36207 vdd.n36206 9.3
R39209 vdd.n36206 vdd.n36205 9.3
R39210 vdd.n36222 vdd.n36221 9.3
R39211 vdd.n36221 vdd.n36220 9.3
R39212 vdd.n36220 vdd.n36219 9.3
R39213 vdd.n36236 vdd.n36235 9.3
R39214 vdd.n36235 vdd.n36234 9.3
R39215 vdd.n36234 vdd.n36233 9.3
R39216 vdd.n36250 vdd.n36249 9.3
R39217 vdd.n36249 vdd.n36248 9.3
R39218 vdd.n36248 vdd.n36247 9.3
R39219 vdd.n36264 vdd.n36263 9.3
R39220 vdd.n36263 vdd.n36262 9.3
R39221 vdd.n36262 vdd.n36261 9.3
R39222 vdd.n36278 vdd.n36277 9.3
R39223 vdd.n36277 vdd.n36276 9.3
R39224 vdd.n36276 vdd.n36275 9.3
R39225 vdd.n36292 vdd.n36291 9.3
R39226 vdd.n36291 vdd.n36290 9.3
R39227 vdd.n36290 vdd.n36289 9.3
R39228 vdd.n36306 vdd.n36305 9.3
R39229 vdd.n36305 vdd.n36304 9.3
R39230 vdd.n36304 vdd.n36303 9.3
R39231 vdd.n36320 vdd.n36319 9.3
R39232 vdd.n36319 vdd.n36318 9.3
R39233 vdd.n36318 vdd.n36317 9.3
R39234 vdd.n36334 vdd.n36333 9.3
R39235 vdd.n36333 vdd.n36332 9.3
R39236 vdd.n36332 vdd.n36331 9.3
R39237 vdd.n36348 vdd.n36347 9.3
R39238 vdd.n36347 vdd.n36346 9.3
R39239 vdd.n36346 vdd.n36345 9.3
R39240 vdd.n36362 vdd.n36361 9.3
R39241 vdd.n36361 vdd.n36360 9.3
R39242 vdd.n36360 vdd.n36359 9.3
R39243 vdd.n36397 vdd.n36396 9.3
R39244 vdd.n36396 vdd.n36395 9.3
R39245 vdd.n36395 vdd.n36394 9.3
R39246 vdd.n36411 vdd.n36410 9.3
R39247 vdd.n36410 vdd.n36409 9.3
R39248 vdd.n36409 vdd.n36408 9.3
R39249 vdd.n36425 vdd.n36424 9.3
R39250 vdd.n36424 vdd.n36423 9.3
R39251 vdd.n36423 vdd.n36422 9.3
R39252 vdd.n36439 vdd.n36438 9.3
R39253 vdd.n36438 vdd.n36437 9.3
R39254 vdd.n36437 vdd.n36436 9.3
R39255 vdd.n36453 vdd.n36452 9.3
R39256 vdd.n36452 vdd.n36451 9.3
R39257 vdd.n36451 vdd.n36450 9.3
R39258 vdd.n36467 vdd.n36466 9.3
R39259 vdd.n36466 vdd.n36465 9.3
R39260 vdd.n36465 vdd.n36464 9.3
R39261 vdd.n36481 vdd.n36480 9.3
R39262 vdd.n36480 vdd.n36479 9.3
R39263 vdd.n36479 vdd.n36478 9.3
R39264 vdd.n36495 vdd.n36494 9.3
R39265 vdd.n36494 vdd.n36493 9.3
R39266 vdd.n36493 vdd.n36492 9.3
R39267 vdd.n36509 vdd.n36508 9.3
R39268 vdd.n36508 vdd.n36507 9.3
R39269 vdd.n36507 vdd.n36506 9.3
R39270 vdd.n36523 vdd.n36522 9.3
R39271 vdd.n36522 vdd.n36521 9.3
R39272 vdd.n36521 vdd.n36520 9.3
R39273 vdd.n36537 vdd.n36536 9.3
R39274 vdd.n36536 vdd.n36535 9.3
R39275 vdd.n36535 vdd.n36534 9.3
R39276 vdd.n36551 vdd.n36550 9.3
R39277 vdd.n36550 vdd.n36549 9.3
R39278 vdd.n36549 vdd.n36548 9.3
R39279 vdd.n36565 vdd.n36564 9.3
R39280 vdd.n36564 vdd.n36563 9.3
R39281 vdd.n36563 vdd.n36562 9.3
R39282 vdd.n36579 vdd.n36578 9.3
R39283 vdd.n36578 vdd.n36577 9.3
R39284 vdd.n36577 vdd.n36576 9.3
R39285 vdd.n36593 vdd.n36592 9.3
R39286 vdd.n36592 vdd.n36591 9.3
R39287 vdd.n36591 vdd.n36590 9.3
R39288 vdd.n36607 vdd.n36606 9.3
R39289 vdd.n36606 vdd.n36605 9.3
R39290 vdd.n36605 vdd.n36604 9.3
R39291 vdd.n36628 vdd.n36627 9.3
R39292 vdd.n36627 vdd.n36626 9.3
R39293 vdd.n36626 vdd.n36625 9.3
R39294 vdd.n36642 vdd.n36641 9.3
R39295 vdd.n36641 vdd.n36640 9.3
R39296 vdd.n36640 vdd.n36639 9.3
R39297 vdd.n36656 vdd.n36655 9.3
R39298 vdd.n36655 vdd.n36654 9.3
R39299 vdd.n36654 vdd.n36653 9.3
R39300 vdd.n36670 vdd.n36669 9.3
R39301 vdd.n36669 vdd.n36668 9.3
R39302 vdd.n36668 vdd.n36667 9.3
R39303 vdd.n36684 vdd.n36683 9.3
R39304 vdd.n36683 vdd.n36682 9.3
R39305 vdd.n36682 vdd.n36681 9.3
R39306 vdd.n36698 vdd.n36697 9.3
R39307 vdd.n36697 vdd.n36696 9.3
R39308 vdd.n36696 vdd.n36695 9.3
R39309 vdd.n36712 vdd.n36711 9.3
R39310 vdd.n36711 vdd.n36710 9.3
R39311 vdd.n36710 vdd.n36709 9.3
R39312 vdd.n36726 vdd.n36725 9.3
R39313 vdd.n36725 vdd.n36724 9.3
R39314 vdd.n36724 vdd.n36723 9.3
R39315 vdd.n36740 vdd.n36739 9.3
R39316 vdd.n36739 vdd.n36738 9.3
R39317 vdd.n36738 vdd.n36737 9.3
R39318 vdd.n36754 vdd.n36753 9.3
R39319 vdd.n36753 vdd.n36752 9.3
R39320 vdd.n36752 vdd.n36751 9.3
R39321 vdd.n36768 vdd.n36767 9.3
R39322 vdd.n36767 vdd.n36766 9.3
R39323 vdd.n36766 vdd.n36765 9.3
R39324 vdd.n36782 vdd.n36781 9.3
R39325 vdd.n36781 vdd.n36780 9.3
R39326 vdd.n36780 vdd.n36779 9.3
R39327 vdd.n36796 vdd.n36795 9.3
R39328 vdd.n36795 vdd.n36794 9.3
R39329 vdd.n36794 vdd.n36793 9.3
R39330 vdd.n36810 vdd.n36809 9.3
R39331 vdd.n36809 vdd.n36808 9.3
R39332 vdd.n36808 vdd.n36807 9.3
R39333 vdd.n36824 vdd.n36823 9.3
R39334 vdd.n36823 vdd.n36822 9.3
R39335 vdd.n36822 vdd.n36821 9.3
R39336 vdd.n36859 vdd.n36858 9.3
R39337 vdd.n36858 vdd.n36857 9.3
R39338 vdd.n36857 vdd.n36856 9.3
R39339 vdd.n36873 vdd.n36872 9.3
R39340 vdd.n36872 vdd.n36871 9.3
R39341 vdd.n36871 vdd.n36870 9.3
R39342 vdd.n36887 vdd.n36886 9.3
R39343 vdd.n36886 vdd.n36885 9.3
R39344 vdd.n36885 vdd.n36884 9.3
R39345 vdd.n36901 vdd.n36900 9.3
R39346 vdd.n36900 vdd.n36899 9.3
R39347 vdd.n36899 vdd.n36898 9.3
R39348 vdd.n36915 vdd.n36914 9.3
R39349 vdd.n36914 vdd.n36913 9.3
R39350 vdd.n36913 vdd.n36912 9.3
R39351 vdd.n36929 vdd.n36928 9.3
R39352 vdd.n36928 vdd.n36927 9.3
R39353 vdd.n36927 vdd.n36926 9.3
R39354 vdd.n36943 vdd.n36942 9.3
R39355 vdd.n36942 vdd.n36941 9.3
R39356 vdd.n36941 vdd.n36940 9.3
R39357 vdd.n36957 vdd.n36956 9.3
R39358 vdd.n36956 vdd.n36955 9.3
R39359 vdd.n36955 vdd.n36954 9.3
R39360 vdd.n36971 vdd.n36970 9.3
R39361 vdd.n36970 vdd.n36969 9.3
R39362 vdd.n36969 vdd.n36968 9.3
R39363 vdd.n35686 vdd.n35685 9.3
R39364 vdd.n37007 vdd.n37006 9.3
R39365 vdd.n37006 vdd.n37005 9.3
R39366 vdd.n37022 vdd.n37021 9.3
R39367 vdd.n37021 vdd.n37020 9.3
R39368 vdd.n37041 vdd.n37040 9.3
R39369 vdd.n37040 vdd.n37039 9.3
R39370 vdd.n33284 vdd.n33283 9.3
R39371 vdd.n33283 vdd.n33282 9.3
R39372 vdd.n37059 vdd.n37058 9.3
R39373 vdd.n37058 vdd.n37057 9.3
R39374 vdd.n37057 vdd.n37056 9.3
R39375 vdd.n33269 vdd.n33268 9.3
R39376 vdd.n33268 vdd.n33267 9.3
R39377 vdd.n33267 vdd.n33266 9.3
R39378 vdd.n33251 vdd.n33250 9.3
R39379 vdd.n33250 vdd.n33249 9.3
R39380 vdd.n33249 vdd.n33248 9.3
R39381 vdd.n37098 vdd.n37097 9.3
R39382 vdd.n37097 vdd.n37096 9.3
R39383 vdd.n37096 vdd.n37095 9.3
R39384 vdd.n33221 vdd.n33220 9.3
R39385 vdd.n33220 vdd.n33219 9.3
R39386 vdd.n33219 vdd.n33218 9.3
R39387 vdd.n37114 vdd.n37113 9.3
R39388 vdd.n37113 vdd.n37112 9.3
R39389 vdd.n33198 vdd.n33197 9.3
R39390 vdd.n33197 vdd.n33196 9.3
R39391 vdd.n33196 vdd.n33195 9.3
R39392 vdd.n33176 vdd.n33175 9.3
R39393 vdd.n33175 vdd.n33174 9.3
R39394 vdd.n33174 vdd.n33173 9.3
R39395 vdd.n37150 vdd.n37149 9.3
R39396 vdd.n37149 vdd.n37148 9.3
R39397 vdd.n33148 vdd.n33147 9.3
R39398 vdd.n33147 vdd.n33146 9.3
R39399 vdd.n35642 vdd.n35641 9.3
R39400 vdd.n35641 vdd.n35640 9.3
R39401 vdd.n37178 vdd.n37177 9.3
R39402 vdd.n37177 vdd.n37176 9.3
R39403 vdd.n33138 vdd.n33137 9.3
R39404 vdd.n33137 vdd.n33136 9.3
R39405 vdd.n33136 vdd.n33135 9.3
R39406 vdd.n37207 vdd.n37206 9.3
R39407 vdd.n37206 vdd.n37205 9.3
R39408 vdd.n37205 vdd.n37204 9.3
R39409 vdd.n33115 vdd.n33114 9.3
R39410 vdd.n33114 vdd.n33113 9.3
R39411 vdd.n37220 vdd.n37219 9.3
R39412 vdd.n37219 vdd.n37218 9.3
R39413 vdd.n37229 vdd.n37228 9.3
R39414 vdd.n37228 vdd.n37227 9.3
R39415 vdd.n37261 vdd.n37260 9.3
R39416 vdd.n37260 vdd.n37259 9.3
R39417 vdd.n37259 vdd.n37258 9.3
R39418 vdd.n33060 vdd.n33059 9.3
R39419 vdd.n33059 vdd.n33058 9.3
R39420 vdd.n33058 vdd.n33057 9.3
R39421 vdd.n37280 vdd.n37279 9.3
R39422 vdd.n37279 vdd.n37278 9.3
R39423 vdd.n37278 vdd.n37277 9.3
R39424 vdd.n33036 vdd.n33035 9.3
R39425 vdd.n33035 vdd.n33034 9.3
R39426 vdd.n33014 vdd.n33013 9.3
R39427 vdd.n33013 vdd.n33012 9.3
R39428 vdd.n37314 vdd.n37313 9.3
R39429 vdd.n37313 vdd.n37312 9.3
R39430 vdd.n32991 vdd.n32990 9.3
R39431 vdd.n32990 vdd.n32989 9.3
R39432 vdd.n37324 vdd.n37323 9.3
R39433 vdd.n37323 vdd.n37322 9.3
R39434 vdd.n37354 vdd.n37353 9.3
R39435 vdd.n37353 vdd.n37352 9.3
R39436 vdd.n32977 vdd.n32976 9.3
R39437 vdd.n32976 vdd.n32975 9.3
R39438 vdd.n37389 vdd.n37388 9.3
R39439 vdd.n37388 vdd.n37387 9.3
R39440 vdd.n37387 vdd.n37386 9.3
R39441 vdd.n32962 vdd.n32961 9.3
R39442 vdd.n32961 vdd.n32960 9.3
R39443 vdd.n32960 vdd.n32959 9.3
R39444 vdd.n37410 vdd.n37409 9.3
R39445 vdd.n37409 vdd.n37408 9.3
R39446 vdd.n37408 vdd.n37407 9.3
R39447 vdd.n37421 vdd.n37420 9.3
R39448 vdd.n37420 vdd.n37419 9.3
R39449 vdd.n37419 vdd.n37418 9.3
R39450 vdd.n32930 vdd.n32929 9.3
R39451 vdd.n32929 vdd.n32928 9.3
R39452 vdd.n32928 vdd.n32927 9.3
R39453 vdd.n37447 vdd.n37446 9.3
R39454 vdd.n37446 vdd.n37445 9.3
R39455 vdd.n37445 vdd.n37444 9.3
R39456 vdd.n32915 vdd.n32914 9.3
R39457 vdd.n32914 vdd.n32913 9.3
R39458 vdd.n32913 vdd.n32912 9.3
R39459 vdd.n37471 vdd.n37470 9.3
R39460 vdd.n37470 vdd.n37469 9.3
R39461 vdd.n37469 vdd.n37468 9.3
R39462 vdd.n37483 vdd.n37482 9.3
R39463 vdd.n37482 vdd.n37481 9.3
R39464 vdd.n37481 vdd.n37480 9.3
R39465 vdd.n32869 vdd.n32868 9.3
R39466 vdd.n32868 vdd.n32867 9.3
R39467 vdd.n37510 vdd.n37509 9.3
R39468 vdd.n37509 vdd.n37508 9.3
R39469 vdd.n32850 vdd.n32849 9.3
R39470 vdd.n32849 vdd.n32848 9.3
R39471 vdd.n32848 vdd.n32847 9.3
R39472 vdd.n37525 vdd.n37524 9.3
R39473 vdd.n37524 vdd.n37523 9.3
R39474 vdd.n35669 vdd.n35668 9.3
R39475 vdd.n35668 vdd.n35667 9.3
R39476 vdd.n32831 vdd.n32830 9.3
R39477 vdd.n32830 vdd.n32829 9.3
R39478 vdd.n37571 vdd.n37570 9.3
R39479 vdd.n37570 vdd.n37569 9.3
R39480 vdd.n38214 vdd.n38213 9.3
R39481 vdd.n38213 vdd.n38212 9.3
R39482 vdd.n38212 vdd.n38211 9.3
R39483 vdd.n38197 vdd.n38196 9.3
R39484 vdd.n38196 vdd.n38195 9.3
R39485 vdd.n38183 vdd.n38182 9.3
R39486 vdd.n38182 vdd.n38181 9.3
R39487 vdd.n38169 vdd.n38168 9.3
R39488 vdd.n38168 vdd.n38167 9.3
R39489 vdd.n38167 vdd.n38166 9.3
R39490 vdd.n38153 vdd.n38152 9.3
R39491 vdd.n38152 vdd.n38151 9.3
R39492 vdd.n38151 vdd.n38150 9.3
R39493 vdd.n38136 vdd.n38135 9.3
R39494 vdd.n38135 vdd.n38134 9.3
R39495 vdd.n38110 vdd.n38109 9.3
R39496 vdd.n38109 vdd.n38108 9.3
R39497 vdd.n38108 vdd.n38107 9.3
R39498 vdd.n38096 vdd.n38095 9.3
R39499 vdd.n38095 vdd.n38094 9.3
R39500 vdd.n38094 vdd.n38093 9.3
R39501 vdd.n38082 vdd.n38081 9.3
R39502 vdd.n38081 vdd.n38080 9.3
R39503 vdd.n38080 vdd.n38079 9.3
R39504 vdd.n38068 vdd.n38067 9.3
R39505 vdd.n38067 vdd.n38066 9.3
R39506 vdd.n38066 vdd.n38065 9.3
R39507 vdd.n38054 vdd.n38053 9.3
R39508 vdd.n38053 vdd.n38052 9.3
R39509 vdd.n38052 vdd.n38051 9.3
R39510 vdd.n38040 vdd.n38039 9.3
R39511 vdd.n38039 vdd.n38038 9.3
R39512 vdd.n38038 vdd.n38037 9.3
R39513 vdd.n38026 vdd.n38025 9.3
R39514 vdd.n38025 vdd.n38024 9.3
R39515 vdd.n38024 vdd.n38023 9.3
R39516 vdd.n38012 vdd.n38011 9.3
R39517 vdd.n38011 vdd.n38010 9.3
R39518 vdd.n38010 vdd.n38009 9.3
R39519 vdd.n37998 vdd.n37997 9.3
R39520 vdd.n37997 vdd.n37996 9.3
R39521 vdd.n37996 vdd.n37995 9.3
R39522 vdd.n37984 vdd.n37983 9.3
R39523 vdd.n37983 vdd.n37982 9.3
R39524 vdd.n37982 vdd.n37981 9.3
R39525 vdd.n37970 vdd.n37969 9.3
R39526 vdd.n37969 vdd.n37968 9.3
R39527 vdd.n37968 vdd.n37967 9.3
R39528 vdd.n37956 vdd.n37955 9.3
R39529 vdd.n37955 vdd.n37954 9.3
R39530 vdd.n37954 vdd.n37953 9.3
R39531 vdd.n37942 vdd.n37941 9.3
R39532 vdd.n37941 vdd.n37940 9.3
R39533 vdd.n37940 vdd.n37939 9.3
R39534 vdd.n37928 vdd.n37927 9.3
R39535 vdd.n37927 vdd.n37926 9.3
R39536 vdd.n37926 vdd.n37925 9.3
R39537 vdd.n37914 vdd.n37913 9.3
R39538 vdd.n37913 vdd.n37912 9.3
R39539 vdd.n37912 vdd.n37911 9.3
R39540 vdd.n37893 vdd.n37892 9.3
R39541 vdd.n37892 vdd.n37891 9.3
R39542 vdd.n37891 vdd.n37890 9.3
R39543 vdd.n37879 vdd.n37878 9.3
R39544 vdd.n37878 vdd.n37877 9.3
R39545 vdd.n37877 vdd.n37876 9.3
R39546 vdd.n37865 vdd.n37864 9.3
R39547 vdd.n37864 vdd.n37863 9.3
R39548 vdd.n37863 vdd.n37862 9.3
R39549 vdd.n37851 vdd.n37850 9.3
R39550 vdd.n37850 vdd.n37849 9.3
R39551 vdd.n37849 vdd.n37848 9.3
R39552 vdd.n37837 vdd.n37836 9.3
R39553 vdd.n37836 vdd.n37835 9.3
R39554 vdd.n37835 vdd.n37834 9.3
R39555 vdd.n37823 vdd.n37822 9.3
R39556 vdd.n37822 vdd.n37821 9.3
R39557 vdd.n37821 vdd.n37820 9.3
R39558 vdd.n37809 vdd.n37808 9.3
R39559 vdd.n37808 vdd.n37807 9.3
R39560 vdd.n37807 vdd.n37806 9.3
R39561 vdd.n37795 vdd.n37794 9.3
R39562 vdd.n37794 vdd.n37793 9.3
R39563 vdd.n37793 vdd.n37792 9.3
R39564 vdd.n37781 vdd.n37780 9.3
R39565 vdd.n37780 vdd.n37779 9.3
R39566 vdd.n37779 vdd.n37778 9.3
R39567 vdd.n37767 vdd.n37766 9.3
R39568 vdd.n37766 vdd.n37765 9.3
R39569 vdd.n37765 vdd.n37764 9.3
R39570 vdd.n37753 vdd.n37752 9.3
R39571 vdd.n37752 vdd.n37751 9.3
R39572 vdd.n37751 vdd.n37750 9.3
R39573 vdd.n37739 vdd.n37738 9.3
R39574 vdd.n37738 vdd.n37737 9.3
R39575 vdd.n37737 vdd.n37736 9.3
R39576 vdd.n37725 vdd.n37724 9.3
R39577 vdd.n37724 vdd.n37723 9.3
R39578 vdd.n37723 vdd.n37722 9.3
R39579 vdd.n37711 vdd.n37710 9.3
R39580 vdd.n37710 vdd.n37709 9.3
R39581 vdd.n37709 vdd.n37708 9.3
R39582 vdd.n37697 vdd.n37696 9.3
R39583 vdd.n37696 vdd.n37695 9.3
R39584 vdd.n37695 vdd.n37694 9.3
R39585 vdd.n37662 vdd.n37661 9.3
R39586 vdd.n37661 vdd.n37660 9.3
R39587 vdd.n37660 vdd.n37659 9.3
R39588 vdd.n37648 vdd.n37647 9.3
R39589 vdd.n37647 vdd.n37646 9.3
R39590 vdd.n37646 vdd.n37645 9.3
R39591 vdd.n37634 vdd.n37633 9.3
R39592 vdd.n37633 vdd.n37632 9.3
R39593 vdd.n37632 vdd.n37631 9.3
R39594 vdd.n37620 vdd.n37619 9.3
R39595 vdd.n37619 vdd.n37618 9.3
R39596 vdd.n37618 vdd.n37617 9.3
R39597 vdd.n37606 vdd.n37605 9.3
R39598 vdd.n37605 vdd.n37604 9.3
R39599 vdd.n37604 vdd.n37603 9.3
R39600 vdd.n28195 vdd.n28194 9.3
R39601 vdd.n28194 vdd.n28193 9.3
R39602 vdd.n28193 vdd.n28192 9.3
R39603 vdd.n28209 vdd.n28208 9.3
R39604 vdd.n28208 vdd.n28207 9.3
R39605 vdd.n28207 vdd.n28206 9.3
R39606 vdd.n28223 vdd.n28222 9.3
R39607 vdd.n28222 vdd.n28221 9.3
R39608 vdd.n28221 vdd.n28220 9.3
R39609 vdd.n28237 vdd.n28236 9.3
R39610 vdd.n28236 vdd.n28235 9.3
R39611 vdd.n28235 vdd.n28234 9.3
R39612 vdd.n28251 vdd.n28250 9.3
R39613 vdd.n28250 vdd.n28249 9.3
R39614 vdd.n28249 vdd.n28248 9.3
R39615 vdd.n28265 vdd.n28264 9.3
R39616 vdd.n28264 vdd.n28263 9.3
R39617 vdd.n28263 vdd.n28262 9.3
R39618 vdd.n28279 vdd.n28278 9.3
R39619 vdd.n28278 vdd.n28277 9.3
R39620 vdd.n28277 vdd.n28276 9.3
R39621 vdd.n28293 vdd.n28292 9.3
R39622 vdd.n28292 vdd.n28291 9.3
R39623 vdd.n28291 vdd.n28290 9.3
R39624 vdd.n28307 vdd.n28306 9.3
R39625 vdd.n28306 vdd.n28305 9.3
R39626 vdd.n28305 vdd.n28304 9.3
R39627 vdd.n28321 vdd.n28320 9.3
R39628 vdd.n28320 vdd.n28319 9.3
R39629 vdd.n28319 vdd.n28318 9.3
R39630 vdd.n28335 vdd.n28334 9.3
R39631 vdd.n28334 vdd.n28333 9.3
R39632 vdd.n28333 vdd.n28332 9.3
R39633 vdd.n28356 vdd.n28355 9.3
R39634 vdd.n28355 vdd.n28354 9.3
R39635 vdd.n28354 vdd.n28353 9.3
R39636 vdd.n28370 vdd.n28369 9.3
R39637 vdd.n28369 vdd.n28368 9.3
R39638 vdd.n28368 vdd.n28367 9.3
R39639 vdd.n28384 vdd.n28383 9.3
R39640 vdd.n28383 vdd.n28382 9.3
R39641 vdd.n28382 vdd.n28381 9.3
R39642 vdd.n28398 vdd.n28397 9.3
R39643 vdd.n28397 vdd.n28396 9.3
R39644 vdd.n28396 vdd.n28395 9.3
R39645 vdd.n28412 vdd.n28411 9.3
R39646 vdd.n28411 vdd.n28410 9.3
R39647 vdd.n28410 vdd.n28409 9.3
R39648 vdd.n28426 vdd.n28425 9.3
R39649 vdd.n28425 vdd.n28424 9.3
R39650 vdd.n28424 vdd.n28423 9.3
R39651 vdd.n28440 vdd.n28439 9.3
R39652 vdd.n28439 vdd.n28438 9.3
R39653 vdd.n28438 vdd.n28437 9.3
R39654 vdd.n28454 vdd.n28453 9.3
R39655 vdd.n28453 vdd.n28452 9.3
R39656 vdd.n28452 vdd.n28451 9.3
R39657 vdd.n28468 vdd.n28467 9.3
R39658 vdd.n28467 vdd.n28466 9.3
R39659 vdd.n28466 vdd.n28465 9.3
R39660 vdd.n28482 vdd.n28481 9.3
R39661 vdd.n28481 vdd.n28480 9.3
R39662 vdd.n28480 vdd.n28479 9.3
R39663 vdd.n28496 vdd.n28495 9.3
R39664 vdd.n28495 vdd.n28494 9.3
R39665 vdd.n28494 vdd.n28493 9.3
R39666 vdd.n28510 vdd.n28509 9.3
R39667 vdd.n28509 vdd.n28508 9.3
R39668 vdd.n28508 vdd.n28507 9.3
R39669 vdd.n28524 vdd.n28523 9.3
R39670 vdd.n28523 vdd.n28522 9.3
R39671 vdd.n28522 vdd.n28521 9.3
R39672 vdd.n28538 vdd.n28537 9.3
R39673 vdd.n28537 vdd.n28536 9.3
R39674 vdd.n28536 vdd.n28535 9.3
R39675 vdd.n28552 vdd.n28551 9.3
R39676 vdd.n28551 vdd.n28550 9.3
R39677 vdd.n28550 vdd.n28549 9.3
R39678 vdd.n28587 vdd.n28586 9.3
R39679 vdd.n28586 vdd.n28585 9.3
R39680 vdd.n28585 vdd.n28584 9.3
R39681 vdd.n28601 vdd.n28600 9.3
R39682 vdd.n28600 vdd.n28599 9.3
R39683 vdd.n28599 vdd.n28598 9.3
R39684 vdd.n28615 vdd.n28614 9.3
R39685 vdd.n28614 vdd.n28613 9.3
R39686 vdd.n28613 vdd.n28612 9.3
R39687 vdd.n28629 vdd.n28628 9.3
R39688 vdd.n28628 vdd.n28627 9.3
R39689 vdd.n28627 vdd.n28626 9.3
R39690 vdd.n28643 vdd.n28642 9.3
R39691 vdd.n28642 vdd.n28641 9.3
R39692 vdd.n28641 vdd.n28640 9.3
R39693 vdd.n28657 vdd.n28656 9.3
R39694 vdd.n28656 vdd.n28655 9.3
R39695 vdd.n28655 vdd.n28654 9.3
R39696 vdd.n28671 vdd.n28670 9.3
R39697 vdd.n28670 vdd.n28669 9.3
R39698 vdd.n28669 vdd.n28668 9.3
R39699 vdd.n28685 vdd.n28684 9.3
R39700 vdd.n28684 vdd.n28683 9.3
R39701 vdd.n28683 vdd.n28682 9.3
R39702 vdd.n28699 vdd.n28698 9.3
R39703 vdd.n28698 vdd.n28697 9.3
R39704 vdd.n28697 vdd.n28696 9.3
R39705 vdd.n28713 vdd.n28712 9.3
R39706 vdd.n28712 vdd.n28711 9.3
R39707 vdd.n28711 vdd.n28710 9.3
R39708 vdd.n28727 vdd.n28726 9.3
R39709 vdd.n28726 vdd.n28725 9.3
R39710 vdd.n28725 vdd.n28724 9.3
R39711 vdd.n28741 vdd.n28740 9.3
R39712 vdd.n28740 vdd.n28739 9.3
R39713 vdd.n28739 vdd.n28738 9.3
R39714 vdd.n28755 vdd.n28754 9.3
R39715 vdd.n28754 vdd.n28753 9.3
R39716 vdd.n28753 vdd.n28752 9.3
R39717 vdd.n28769 vdd.n28768 9.3
R39718 vdd.n28768 vdd.n28767 9.3
R39719 vdd.n28767 vdd.n28766 9.3
R39720 vdd.n28783 vdd.n28782 9.3
R39721 vdd.n28782 vdd.n28781 9.3
R39722 vdd.n28781 vdd.n28780 9.3
R39723 vdd.n28797 vdd.n28796 9.3
R39724 vdd.n28796 vdd.n28795 9.3
R39725 vdd.n28795 vdd.n28794 9.3
R39726 vdd.n28153 vdd.n28152 9.3
R39727 vdd.n28152 vdd.n28151 9.3
R39728 vdd.n28165 vdd.n28164 9.3
R39729 vdd.n28164 vdd.n28163 9.3
R39730 vdd.n28175 vdd.n28174 9.3
R39731 vdd.n28174 vdd.n28173 9.3
R39732 vdd.n28140 vdd.n28139 9.3
R39733 vdd.n28139 vdd.n28138 9.3
R39734 vdd.n28813 vdd.n28812 9.3
R39735 vdd.n28812 vdd.n28811 9.3
R39736 vdd.n26210 vdd.n26209 9.3
R39737 vdd.n28115 vdd.n28114 9.3
R39738 vdd.n28114 vdd.n28113 9.3
R39739 vdd.n26701 vdd.n26700 9.3
R39740 vdd.n26310 vdd.n26309 9.3
R39741 vdd.n28089 vdd.n28088 9.3
R39742 vdd.n28088 vdd.n28087 9.3
R39743 vdd.n31755 vdd.n31754 9.3
R39744 vdd.n28065 vdd.n28064 9.3
R39745 vdd.n28064 vdd.n28063 9.3
R39746 vdd.n28969 vdd.n28968 9.3
R39747 vdd.n28968 vdd.n28967 9.3
R39748 vdd.n28967 vdd.n28966 9.3
R39749 vdd.n28990 vdd.n28989 9.3
R39750 vdd.n28989 vdd.n28988 9.3
R39751 vdd.n31846 vdd.n31845 9.3
R39752 vdd.n31891 vdd.n31890 9.3
R39753 vdd.n29030 vdd.n29029 9.3
R39754 vdd.n29029 vdd.n29028 9.3
R39755 vdd.n27794 vdd.n27793 9.3
R39756 vdd.n27793 vdd.n27792 9.3
R39757 vdd.n27811 vdd.n27810 9.3
R39758 vdd.n27810 vdd.n27809 9.3
R39759 vdd.n31658 vdd.n31657 9.3
R39760 vdd.n27839 vdd.n27838 9.3
R39761 vdd.n27838 vdd.n27837 9.3
R39762 vdd.n31629 vdd.n31628 9.3
R39763 vdd.n27986 vdd.n27985 9.3
R39764 vdd.n27985 vdd.n27984 9.3
R39765 vdd.n27883 vdd.n27882 9.3
R39766 vdd.n27882 vdd.n27881 9.3
R39767 vdd.n32067 vdd.n32066 9.3
R39768 vdd.n27915 vdd.n27914 9.3
R39769 vdd.n27914 vdd.n27913 9.3
R39770 vdd.n27934 vdd.n27933 9.3
R39771 vdd.n27933 vdd.n27932 9.3
R39772 vdd.n29887 vdd.n29886 9.3
R39773 vdd.n29886 vdd.n29885 9.3
R39774 vdd.n31572 vdd.n31571 9.3
R39775 vdd.n29873 vdd.n29872 9.3
R39776 vdd.n29872 vdd.n29871 9.3
R39777 vdd.n29871 vdd.n29870 9.3
R39778 vdd.n32229 vdd.n32228 9.3
R39779 vdd.n29694 vdd.n29693 9.3
R39780 vdd.n29693 vdd.n29692 9.3
R39781 vdd.n29839 vdd.n29838 9.3
R39782 vdd.n29838 vdd.n29837 9.3
R39783 vdd.n29837 vdd.n29836 9.3
R39784 vdd.n29819 vdd.n29818 9.3
R39785 vdd.n29818 vdd.n29817 9.3
R39786 vdd.n31512 vdd.n31511 9.3
R39787 vdd.n29765 vdd.n29764 9.3
R39788 vdd.n29764 vdd.n29763 9.3
R39789 vdd.n31488 vdd.n31487 9.3
R39790 vdd.n29723 vdd.n29722 9.3
R39791 vdd.n29722 vdd.n29721 9.3
R39792 vdd.n31460 vdd.n31459 9.3
R39793 vdd.n32403 vdd.n32402 9.3
R39794 vdd.n30191 vdd.n30190 9.3
R39795 vdd.n30190 vdd.n30189 9.3
R39796 vdd.n30223 vdd.n30222 9.3
R39797 vdd.n30222 vdd.n30221 9.3
R39798 vdd.n30221 vdd.n30220 9.3
R39799 vdd.n30238 vdd.n30237 9.3
R39800 vdd.n30237 vdd.n30236 9.3
R39801 vdd.n30236 vdd.n30235 9.3
R39802 vdd.n32447 vdd.n32446 9.3
R39803 vdd.n30274 vdd.n30273 9.3
R39804 vdd.n30273 vdd.n30272 9.3
R39805 vdd.n31094 vdd.n31093 9.3
R39806 vdd.n30569 vdd.n30568 9.3
R39807 vdd.n30568 vdd.n30567 9.3
R39808 vdd.n30567 vdd.n30566 9.3
R39809 vdd.n30548 vdd.n30547 9.3
R39810 vdd.n30547 vdd.n30546 9.3
R39811 vdd.n30546 vdd.n30545 9.3
R39812 vdd.n30531 vdd.n30530 9.3
R39813 vdd.n30530 vdd.n30529 9.3
R39814 vdd.n30517 vdd.n30516 9.3
R39815 vdd.n30516 vdd.n30515 9.3
R39816 vdd.n30341 vdd.n30340 9.3
R39817 vdd.n30340 vdd.n30339 9.3
R39818 vdd.n30505 vdd.n30504 9.3
R39819 vdd.n30504 vdd.n30503 9.3
R39820 vdd.n1817 vdd.n1816 9.3
R39821 vdd.n1980 vdd.n1979 9.3
R39822 vdd.n1979 vdd.n1978 9.3
R39823 vdd.n2624 vdd.n2623 9.3
R39824 vdd.n2623 vdd.n2622 9.3
R39825 vdd.n2480 vdd.n2479 9.3
R39826 vdd.n2479 vdd.n2478 9.3
R39827 vdd.n2196 vdd.n2195 9.3
R39828 vdd.n2195 vdd.n2194 9.3
R39829 vdd.n2219 vdd.n2218 9.3
R39830 vdd.n2218 vdd.n2217 9.3
R39831 vdd.n3815 vdd.n3814 9.3
R39832 vdd.n3711 vdd.n3710 9.3
R39833 vdd.n3710 vdd.n3709 9.3
R39834 vdd.n2722 vdd.n2721 9.3
R39835 vdd.n2721 vdd.n2720 9.3
R39836 vdd.n2750 vdd.n2749 9.3
R39837 vdd.n2749 vdd.n2748 9.3
R39838 vdd.n2761 vdd.n2760 9.3
R39839 vdd.n2760 vdd.n2759 9.3
R39840 vdd.n2772 vdd.n2771 9.3
R39841 vdd.n2771 vdd.n2770 9.3
R39842 vdd.n2783 vdd.n2782 9.3
R39843 vdd.n2782 vdd.n2781 9.3
R39844 vdd.n2794 vdd.n2793 9.3
R39845 vdd.n2793 vdd.n2792 9.3
R39846 vdd.n2811 vdd.n2810 9.3
R39847 vdd.n2810 vdd.n2809 9.3
R39848 vdd.n2822 vdd.n2821 9.3
R39849 vdd.n2821 vdd.n2820 9.3
R39850 vdd.n2833 vdd.n2832 9.3
R39851 vdd.n2832 vdd.n2831 9.3
R39852 vdd.n2844 vdd.n2843 9.3
R39853 vdd.n2843 vdd.n2842 9.3
R39854 vdd.n2855 vdd.n2854 9.3
R39855 vdd.n2854 vdd.n2853 9.3
R39856 vdd.n2866 vdd.n2865 9.3
R39857 vdd.n2865 vdd.n2864 9.3
R39858 vdd.n2877 vdd.n2876 9.3
R39859 vdd.n2876 vdd.n2875 9.3
R39860 vdd.n2888 vdd.n2887 9.3
R39861 vdd.n2887 vdd.n2886 9.3
R39862 vdd.n2898 vdd.n2897 9.3
R39863 vdd.n2897 vdd.n2896 9.3
R39864 vdd.n2909 vdd.n2908 9.3
R39865 vdd.n2908 vdd.n2907 9.3
R39866 vdd.n2920 vdd.n2919 9.3
R39867 vdd.n2919 vdd.n2918 9.3
R39868 vdd.n2931 vdd.n2930 9.3
R39869 vdd.n2930 vdd.n2929 9.3
R39870 vdd.n2942 vdd.n2941 9.3
R39871 vdd.n2941 vdd.n2940 9.3
R39872 vdd.n2953 vdd.n2952 9.3
R39873 vdd.n2952 vdd.n2951 9.3
R39874 vdd.n2964 vdd.n2963 9.3
R39875 vdd.n2963 vdd.n2962 9.3
R39876 vdd.n2975 vdd.n2974 9.3
R39877 vdd.n2974 vdd.n2973 9.3
R39878 vdd.n2992 vdd.n2991 9.3
R39879 vdd.n2991 vdd.n2990 9.3
R39880 vdd.n3003 vdd.n3002 9.3
R39881 vdd.n3002 vdd.n3001 9.3
R39882 vdd.n3014 vdd.n3013 9.3
R39883 vdd.n3013 vdd.n3012 9.3
R39884 vdd.n3025 vdd.n3024 9.3
R39885 vdd.n3024 vdd.n3023 9.3
R39886 vdd.n3036 vdd.n3035 9.3
R39887 vdd.n3035 vdd.n3034 9.3
R39888 vdd.n3047 vdd.n3046 9.3
R39889 vdd.n3046 vdd.n3045 9.3
R39890 vdd.n3058 vdd.n3057 9.3
R39891 vdd.n3057 vdd.n3056 9.3
R39892 vdd.n3069 vdd.n3068 9.3
R39893 vdd.n3068 vdd.n3067 9.3
R39894 vdd.n3079 vdd.n3078 9.3
R39895 vdd.n3078 vdd.n3077 9.3
R39896 vdd.n3090 vdd.n3089 9.3
R39897 vdd.n3089 vdd.n3088 9.3
R39898 vdd.n3101 vdd.n3100 9.3
R39899 vdd.n3100 vdd.n3099 9.3
R39900 vdd.n3112 vdd.n3111 9.3
R39901 vdd.n3111 vdd.n3110 9.3
R39902 vdd.n3123 vdd.n3122 9.3
R39903 vdd.n3122 vdd.n3121 9.3
R39904 vdd.n3134 vdd.n3133 9.3
R39905 vdd.n3133 vdd.n3132 9.3
R39906 vdd.n3145 vdd.n3144 9.3
R39907 vdd.n3144 vdd.n3143 9.3
R39908 vdd.n3156 vdd.n3155 9.3
R39909 vdd.n3155 vdd.n3154 9.3
R39910 vdd.n3173 vdd.n3172 9.3
R39911 vdd.n3172 vdd.n3171 9.3
R39912 vdd.n3184 vdd.n3183 9.3
R39913 vdd.n3183 vdd.n3182 9.3
R39914 vdd.n3195 vdd.n3194 9.3
R39915 vdd.n3194 vdd.n3193 9.3
R39916 vdd.n3206 vdd.n3205 9.3
R39917 vdd.n3205 vdd.n3204 9.3
R39918 vdd.n3217 vdd.n3216 9.3
R39919 vdd.n3216 vdd.n3215 9.3
R39920 vdd.n3228 vdd.n3227 9.3
R39921 vdd.n3227 vdd.n3226 9.3
R39922 vdd.n3239 vdd.n3238 9.3
R39923 vdd.n3238 vdd.n3237 9.3
R39924 vdd.n3250 vdd.n3249 9.3
R39925 vdd.n3249 vdd.n3248 9.3
R39926 vdd.n3260 vdd.n3259 9.3
R39927 vdd.n3259 vdd.n3258 9.3
R39928 vdd.n3271 vdd.n3270 9.3
R39929 vdd.n3270 vdd.n3269 9.3
R39930 vdd.n3282 vdd.n3281 9.3
R39931 vdd.n3281 vdd.n3280 9.3
R39932 vdd.n3293 vdd.n3292 9.3
R39933 vdd.n3292 vdd.n3291 9.3
R39934 vdd.n3304 vdd.n3303 9.3
R39935 vdd.n3303 vdd.n3302 9.3
R39936 vdd.n3315 vdd.n3314 9.3
R39937 vdd.n3314 vdd.n3313 9.3
R39938 vdd.n3326 vdd.n3325 9.3
R39939 vdd.n3325 vdd.n3324 9.3
R39940 vdd.n3337 vdd.n3336 9.3
R39941 vdd.n3336 vdd.n3335 9.3
R39942 vdd.n3354 vdd.n3353 9.3
R39943 vdd.n3353 vdd.n3352 9.3
R39944 vdd.n3365 vdd.n3364 9.3
R39945 vdd.n3364 vdd.n3363 9.3
R39946 vdd.n3376 vdd.n3375 9.3
R39947 vdd.n3375 vdd.n3374 9.3
R39948 vdd.n3387 vdd.n3386 9.3
R39949 vdd.n3386 vdd.n3385 9.3
R39950 vdd.n3398 vdd.n3397 9.3
R39951 vdd.n3397 vdd.n3396 9.3
R39952 vdd.n3409 vdd.n3408 9.3
R39953 vdd.n3408 vdd.n3407 9.3
R39954 vdd.n3420 vdd.n3419 9.3
R39955 vdd.n3419 vdd.n3418 9.3
R39956 vdd.n3431 vdd.n3430 9.3
R39957 vdd.n3430 vdd.n3429 9.3
R39958 vdd.n3441 vdd.n3440 9.3
R39959 vdd.n3440 vdd.n3439 9.3
R39960 vdd.n3452 vdd.n3451 9.3
R39961 vdd.n3451 vdd.n3450 9.3
R39962 vdd.n3463 vdd.n3462 9.3
R39963 vdd.n3462 vdd.n3461 9.3
R39964 vdd.n3474 vdd.n3473 9.3
R39965 vdd.n3473 vdd.n3472 9.3
R39966 vdd.n3485 vdd.n3484 9.3
R39967 vdd.n3484 vdd.n3483 9.3
R39968 vdd.n3496 vdd.n3495 9.3
R39969 vdd.n3495 vdd.n3494 9.3
R39970 vdd.n3507 vdd.n3506 9.3
R39971 vdd.n3506 vdd.n3505 9.3
R39972 vdd.n3518 vdd.n3517 9.3
R39973 vdd.n3517 vdd.n3516 9.3
R39974 vdd.n3535 vdd.n3534 9.3
R39975 vdd.n3534 vdd.n3533 9.3
R39976 vdd.n3546 vdd.n3545 9.3
R39977 vdd.n3545 vdd.n3544 9.3
R39978 vdd.n3557 vdd.n3556 9.3
R39979 vdd.n3556 vdd.n3555 9.3
R39980 vdd.n3568 vdd.n3567 9.3
R39981 vdd.n3567 vdd.n3566 9.3
R39982 vdd.n3579 vdd.n3578 9.3
R39983 vdd.n3578 vdd.n3577 9.3
R39984 vdd.n3590 vdd.n3589 9.3
R39985 vdd.n3589 vdd.n3588 9.3
R39986 vdd.n3601 vdd.n3600 9.3
R39987 vdd.n3600 vdd.n3599 9.3
R39988 vdd.n3612 vdd.n3611 9.3
R39989 vdd.n3611 vdd.n3610 9.3
R39990 vdd.n3622 vdd.n3621 9.3
R39991 vdd.n3621 vdd.n3620 9.3
R39992 vdd.n3645 vdd.n3644 9.3
R39993 vdd.n3644 vdd.n3643 9.3
R39994 vdd.n3655 vdd.n3654 9.3
R39995 vdd.n3654 vdd.n3653 9.3
R39996 vdd.n3635 vdd.n3634 9.3
R39997 vdd.n3634 vdd.n3633 9.3
R39998 vdd.n2056 vdd.n2055 9.3
R39999 vdd.n2055 vdd.n2054 9.3
R40000 vdd.n3692 vdd.n3691 9.3
R40001 vdd.n3691 vdd.n3690 9.3
R40002 vdd.n4012 vdd.n4011 9.3
R40003 vdd.n4011 vdd.n4010 9.3
R40004 vdd.n3997 vdd.n3996 9.3
R40005 vdd.n3996 vdd.n3995 9.3
R40006 vdd.n3982 vdd.n3981 9.3
R40007 vdd.n3981 vdd.n3980 9.3
R40008 vdd.n2014 vdd.n2013 9.3
R40009 vdd.n2013 vdd.n2012 9.3
R40010 vdd.n3955 vdd.n3954 9.3
R40011 vdd.n3954 vdd.n3953 9.3
R40012 vdd.n3938 vdd.n3937 9.3
R40013 vdd.n3937 vdd.n3936 9.3
R40014 vdd.n3921 vdd.n3920 9.3
R40015 vdd.n3920 vdd.n3919 9.3
R40016 vdd.n3898 vdd.n3897 9.3
R40017 vdd.n3855 vdd.n3854 9.3
R40018 vdd.n3854 vdd.n3853 9.3
R40019 vdd.n2241 vdd.n2240 9.3
R40020 vdd.n2240 vdd.n2239 9.3
R40021 vdd.n2179 vdd.n2178 9.3
R40022 vdd.n2178 vdd.n2177 9.3
R40023 vdd.n2158 vdd.n2157 9.3
R40024 vdd.n2157 vdd.n2156 9.3
R40025 vdd.n2284 vdd.n2283 9.3
R40026 vdd.n2283 vdd.n2282 9.3
R40027 vdd.n2303 vdd.n2302 9.3
R40028 vdd.n2302 vdd.n2301 9.3
R40029 vdd.n2322 vdd.n2321 9.3
R40030 vdd.n2321 vdd.n2320 9.3
R40031 vdd.n2341 vdd.n2340 9.3
R40032 vdd.n2340 vdd.n2339 9.3
R40033 vdd.n2040 vdd.n2039 9.3
R40034 vdd.n2039 vdd.n2038 9.3
R40035 vdd.n2380 vdd.n2379 9.3
R40036 vdd.n2379 vdd.n2378 9.3
R40037 vdd.n2404 vdd.n2403 9.3
R40038 vdd.n2403 vdd.n2402 9.3
R40039 vdd.n2420 vdd.n2419 9.3
R40040 vdd.n2526 vdd.n2525 9.3
R40041 vdd.n2497 vdd.n2496 9.3
R40042 vdd.n2496 vdd.n2495 9.3
R40043 vdd.n2602 vdd.n2601 9.3
R40044 vdd.n2601 vdd.n2600 9.3
R40045 vdd.n2637 vdd.n2636 9.3
R40046 vdd.n2636 vdd.n2635 9.3
R40047 vdd.n2656 vdd.n2655 9.3
R40048 vdd.n2655 vdd.n2654 9.3
R40049 vdd.n2665 vdd.n2567 9.3
R40050 vdd.n2567 vdd.n2566 9.3
R40051 vdd.n1990 vdd.n1989 9.3
R40052 vdd.n1989 vdd.n1988 9.3
R40053 vdd.n2082 vdd.n2072 9.3
R40054 vdd.n2072 vdd.n2071 9.3
R40055 vdd.n1950 vdd.n1938 9.3
R40056 vdd.n1938 vdd.n1937 9.3
R40057 vdd.n1197 vdd.n1196 9.3
R40058 vdd.n1196 vdd.n1195 9.3
R40059 vdd.n1908 vdd.n1907 9.3
R40060 vdd.n1907 vdd.n1906 9.3
R40061 vdd.n1225 vdd.n1224 9.3
R40062 vdd.n1866 vdd.n1865 9.3
R40063 vdd.n1865 vdd.n1864 9.3
R40064 vdd.n1241 vdd.n1240 9.3
R40065 vdd.n1799 vdd.n1798 9.3
R40066 vdd.n1798 vdd.n1797 9.3
R40067 vdd.n1783 vdd.n1782 9.3
R40068 vdd.n1782 vdd.n1781 9.3
R40069 vdd.n1273 vdd.n1272 9.3
R40070 vdd.n1272 vdd.n1271 9.3
R40071 vdd.n1284 vdd.n1283 9.3
R40072 vdd.n1283 vdd.n1282 9.3
R40073 vdd.n1770 vdd.n1769 9.3
R40074 vdd.n1769 vdd.n1768 9.3
R40075 vdd.n1759 vdd.n1758 9.3
R40076 vdd.n1758 vdd.n1757 9.3
R40077 vdd.n1739 vdd.n1738 9.3
R40078 vdd.n1746 vdd.n1745 9.3
R40079 vdd.n1726 vdd.n1725 9.3
R40080 vdd.n1725 vdd.n1724 9.3
R40081 vdd.n1715 vdd.n1714 9.3
R40082 vdd.n1714 vdd.n1713 9.3
R40083 vdd.n1704 vdd.n1703 9.3
R40084 vdd.n1703 vdd.n1702 9.3
R40085 vdd.n1693 vdd.n1692 9.3
R40086 vdd.n1692 vdd.n1691 9.3
R40087 vdd.n1682 vdd.n1681 9.3
R40088 vdd.n1681 vdd.n1680 9.3
R40089 vdd.n1671 vdd.n1670 9.3
R40090 vdd.n1670 vdd.n1669 9.3
R40091 vdd.n1660 vdd.n1659 9.3
R40092 vdd.n1659 vdd.n1658 9.3
R40093 vdd.n1650 vdd.n1649 9.3
R40094 vdd.n1649 vdd.n1648 9.3
R40095 vdd.n1639 vdd.n1638 9.3
R40096 vdd.n1638 vdd.n1637 9.3
R40097 vdd.n1628 vdd.n1627 9.3
R40098 vdd.n1627 vdd.n1626 9.3
R40099 vdd.n1617 vdd.n1616 9.3
R40100 vdd.n1616 vdd.n1615 9.3
R40101 vdd.n1606 vdd.n1605 9.3
R40102 vdd.n1605 vdd.n1604 9.3
R40103 vdd.n1595 vdd.n1594 9.3
R40104 vdd.n1594 vdd.n1593 9.3
R40105 vdd.n1584 vdd.n1583 9.3
R40106 vdd.n1583 vdd.n1582 9.3
R40107 vdd.n1573 vdd.n1572 9.3
R40108 vdd.n1572 vdd.n1571 9.3
R40109 vdd.n1556 vdd.n1555 9.3
R40110 vdd.n1555 vdd.n1554 9.3
R40111 vdd.n1545 vdd.n1544 9.3
R40112 vdd.n1544 vdd.n1543 9.3
R40113 vdd.n1534 vdd.n1533 9.3
R40114 vdd.n1533 vdd.n1532 9.3
R40115 vdd.n1523 vdd.n1522 9.3
R40116 vdd.n1522 vdd.n1521 9.3
R40117 vdd.n1512 vdd.n1511 9.3
R40118 vdd.n1511 vdd.n1510 9.3
R40119 vdd.n1501 vdd.n1500 9.3
R40120 vdd.n1500 vdd.n1499 9.3
R40121 vdd.n1490 vdd.n1489 9.3
R40122 vdd.n1489 vdd.n1488 9.3
R40123 vdd.n1479 vdd.n1478 9.3
R40124 vdd.n1478 vdd.n1477 9.3
R40125 vdd.n1469 vdd.n1468 9.3
R40126 vdd.n1468 vdd.n1467 9.3
R40127 vdd.n1458 vdd.n1457 9.3
R40128 vdd.n1457 vdd.n1456 9.3
R40129 vdd.n1447 vdd.n1446 9.3
R40130 vdd.n1446 vdd.n1445 9.3
R40131 vdd.n1436 vdd.n1435 9.3
R40132 vdd.n1435 vdd.n1434 9.3
R40133 vdd.n1425 vdd.n1424 9.3
R40134 vdd.n1424 vdd.n1423 9.3
R40135 vdd.n1414 vdd.n1413 9.3
R40136 vdd.n1413 vdd.n1412 9.3
R40137 vdd.n1403 vdd.n1402 9.3
R40138 vdd.n1402 vdd.n1401 9.3
R40139 vdd.n1392 vdd.n1391 9.3
R40140 vdd.n1391 vdd.n1390 9.3
R40141 vdd.n1375 vdd.n1374 9.3
R40142 vdd.n1374 vdd.n1373 9.3
R40143 vdd.n1364 vdd.n1363 9.3
R40144 vdd.n1363 vdd.n1362 9.3
R40145 vdd.n1353 vdd.n1352 9.3
R40146 vdd.n1352 vdd.n1351 9.3
R40147 vdd.n1342 vdd.n1341 9.3
R40148 vdd.n1341 vdd.n1340 9.3
R40149 vdd.n1331 vdd.n1330 9.3
R40150 vdd.n1330 vdd.n1329 9.3
R40151 vdd.n1320 vdd.n1319 9.3
R40152 vdd.n1319 vdd.n1318 9.3
R40153 vdd.n1309 vdd.n1308 9.3
R40154 vdd.n1308 vdd.n1307 9.3
R40155 vdd.n1298 vdd.n1297 9.3
R40156 vdd.n1297 vdd.n1296 9.3
R40157 vdd.n26764 vdd.n26763 9.3
R40158 vdd.n26763 vdd.n26762 9.3
R40159 vdd.n26775 vdd.n26774 9.3
R40160 vdd.n26774 vdd.n26773 9.3
R40161 vdd.n26786 vdd.n26785 9.3
R40162 vdd.n26785 vdd.n26784 9.3
R40163 vdd.n26797 vdd.n26796 9.3
R40164 vdd.n26796 vdd.n26795 9.3
R40165 vdd.n26808 vdd.n26807 9.3
R40166 vdd.n26807 vdd.n26806 9.3
R40167 vdd.n26819 vdd.n26818 9.3
R40168 vdd.n26818 vdd.n26817 9.3
R40169 vdd.n26830 vdd.n26829 9.3
R40170 vdd.n26829 vdd.n26828 9.3
R40171 vdd.n26841 vdd.n26840 9.3
R40172 vdd.n26840 vdd.n26839 9.3
R40173 vdd.n26858 vdd.n26857 9.3
R40174 vdd.n26857 vdd.n26856 9.3
R40175 vdd.n26869 vdd.n26868 9.3
R40176 vdd.n26868 vdd.n26867 9.3
R40177 vdd.n26880 vdd.n26879 9.3
R40178 vdd.n26879 vdd.n26878 9.3
R40179 vdd.n26891 vdd.n26890 9.3
R40180 vdd.n26890 vdd.n26889 9.3
R40181 vdd.n26902 vdd.n26901 9.3
R40182 vdd.n26901 vdd.n26900 9.3
R40183 vdd.n26913 vdd.n26912 9.3
R40184 vdd.n26912 vdd.n26911 9.3
R40185 vdd.n26924 vdd.n26923 9.3
R40186 vdd.n26923 vdd.n26922 9.3
R40187 vdd.n26935 vdd.n26934 9.3
R40188 vdd.n26934 vdd.n26933 9.3
R40189 vdd.n26945 vdd.n26944 9.3
R40190 vdd.n26944 vdd.n26943 9.3
R40191 vdd.n26956 vdd.n26955 9.3
R40192 vdd.n26955 vdd.n26954 9.3
R40193 vdd.n26967 vdd.n26966 9.3
R40194 vdd.n26966 vdd.n26965 9.3
R40195 vdd.n26978 vdd.n26977 9.3
R40196 vdd.n26977 vdd.n26976 9.3
R40197 vdd.n26989 vdd.n26988 9.3
R40198 vdd.n26988 vdd.n26987 9.3
R40199 vdd.n27000 vdd.n26999 9.3
R40200 vdd.n26999 vdd.n26998 9.3
R40201 vdd.n27011 vdd.n27010 9.3
R40202 vdd.n27010 vdd.n27009 9.3
R40203 vdd.n27022 vdd.n27021 9.3
R40204 vdd.n27021 vdd.n27020 9.3
R40205 vdd.n27039 vdd.n27038 9.3
R40206 vdd.n27038 vdd.n27037 9.3
R40207 vdd.n27050 vdd.n27049 9.3
R40208 vdd.n27049 vdd.n27048 9.3
R40209 vdd.n27061 vdd.n27060 9.3
R40210 vdd.n27060 vdd.n27059 9.3
R40211 vdd.n27072 vdd.n27071 9.3
R40212 vdd.n27071 vdd.n27070 9.3
R40213 vdd.n27083 vdd.n27082 9.3
R40214 vdd.n27082 vdd.n27081 9.3
R40215 vdd.n27094 vdd.n27093 9.3
R40216 vdd.n27093 vdd.n27092 9.3
R40217 vdd.n27105 vdd.n27104 9.3
R40218 vdd.n27104 vdd.n27103 9.3
R40219 vdd.n27116 vdd.n27115 9.3
R40220 vdd.n27115 vdd.n27114 9.3
R40221 vdd.n27126 vdd.n27125 9.3
R40222 vdd.n27125 vdd.n27124 9.3
R40223 vdd.n27137 vdd.n27136 9.3
R40224 vdd.n27136 vdd.n27135 9.3
R40225 vdd.n27148 vdd.n27147 9.3
R40226 vdd.n27147 vdd.n27146 9.3
R40227 vdd.n27159 vdd.n27158 9.3
R40228 vdd.n27158 vdd.n27157 9.3
R40229 vdd.n27170 vdd.n27169 9.3
R40230 vdd.n27169 vdd.n27168 9.3
R40231 vdd.n27181 vdd.n27180 9.3
R40232 vdd.n27180 vdd.n27179 9.3
R40233 vdd.n27192 vdd.n27191 9.3
R40234 vdd.n27191 vdd.n27190 9.3
R40235 vdd.n27203 vdd.n27202 9.3
R40236 vdd.n27202 vdd.n27201 9.3
R40237 vdd.n26745 vdd.n26744 9.3
R40238 vdd.n26737 vdd.n26736 9.3
R40239 vdd.n26755 vdd.n26754 9.3
R40240 vdd.n26754 vdd.n26753 9.3
R40241 vdd.n31279 vdd.n31268 9.3
R40242 vdd.n31268 vdd.n31267 9.3
R40243 vdd.n31260 vdd.n31259 9.3
R40244 vdd.n31259 vdd.n31258 9.3
R40245 vdd.n31277 vdd.n31276 9.3
R40246 vdd.n31276 vdd.n31275 9.3
R40247 vdd.n31156 vdd.n31155 9.3
R40248 vdd.n31147 vdd.n31146 9.3
R40249 vdd.n2741 vdd.n2740 9.3
R40250 vdd.n31693 vdd.n31692 9.3
R40251 vdd.n31933 vdd.n31932 9.3
R40252 vdd.n26193 vdd.n26191 9.3
R40253 vdd.n26595 vdd.n26593 9.3
R40254 vdd.n26608 vdd.n26606 9.3
R40255 vdd.n26682 vdd.n26677 9.3
R40256 vdd.n26296 vdd.n26294 9.3
R40257 vdd.n26336 vdd.n26331 9.3
R40258 vdd.n31794 vdd.n31792 9.3
R40259 vdd.n31814 vdd.n31812 9.3
R40260 vdd.n31833 vdd.n31831 9.3
R40261 vdd.n31858 vdd.n31856 9.3
R40262 vdd.n31875 vdd.n31873 9.3
R40263 vdd.n31900 vdd.n31898 9.3
R40264 vdd.n31973 vdd.n31645 9.3
R40265 vdd.n31988 vdd.n31633 9.3
R40266 vdd.n32007 vdd.n32005 9.3
R40267 vdd.n32019 vdd.n32017 9.3
R40268 vdd.n32037 vdd.n32035 9.3
R40269 vdd.n32050 vdd.n32048 9.3
R40270 vdd.n32144 vdd.n32142 9.3
R40271 vdd.n32172 vdd.n32170 9.3
R40272 vdd.n32194 vdd.n32192 9.3
R40273 vdd.n32216 vdd.n32214 9.3
R40274 vdd.n32248 vdd.n32246 9.3
R40275 vdd.n32265 vdd.n32263 9.3
R40276 vdd.n32331 vdd.n31493 9.3
R40277 vdd.n32348 vdd.n31477 9.3
R40278 vdd.n32362 vdd.n32360 9.3
R40279 vdd.n32378 vdd.n32376 9.3
R40280 vdd.n32533 vdd.n32391 9.3
R40281 vdd.n32517 vdd.n32411 9.3
R40282 vdd.n32459 vdd.n32435 9.3
R40283 vdd.n31058 vdd.n31056 9.3
R40284 vdd.n31081 vdd.n31079 9.3
R40285 vdd.n31110 vdd.n31108 9.3
R40286 vdd.n31186 vdd.n31125 9.3
R40287 vdd.n31184 vdd.n31127 9.3
R40288 vdd.n31124 vdd.n31122 9.3
R40289 vdd.n31086 vdd.n31083 9.3
R40290 vdd.n31078 vdd.n31076 9.3
R40291 vdd.n32457 vdd.n32437 9.3
R40292 vdd.n32461 vdd.n32434 9.3
R40293 vdd.n32531 vdd.n32392 9.3
R40294 vdd.n32365 vdd.n32363 9.3
R40295 vdd.n32334 vdd.n32332 9.3
R40296 vdd.n32287 vdd.n32285 9.3
R40297 vdd.n32253 vdd.n32250 9.3
R40298 vdd.n32236 vdd.n32234 9.3
R40299 vdd.n32199 vdd.n32196 9.3
R40300 vdd.n32191 vdd.n32189 9.3
R40301 vdd.n32149 vdd.n32146 9.3
R40302 vdd.n32141 vdd.n32139 9.3
R40303 vdd.n32040 vdd.n32038 9.3
R40304 vdd.n32010 vdd.n32008 9.3
R40305 vdd.n31976 vdd.n31974 9.3
R40306 vdd.n31915 vdd.n31913 9.3
R40307 vdd.n31880 vdd.n31877 9.3
R40308 vdd.n31872 vdd.n31870 9.3
R40309 vdd.n31838 vdd.n31835 9.3
R40310 vdd.n31830 vdd.n31828 9.3
R40311 vdd.n31799 vdd.n31796 9.3
R40312 vdd.n31791 vdd.n31789 9.3
R40313 vdd.n26316 vdd.n26314 9.3
R40314 vdd.n26690 vdd.n26688 9.3
R40315 vdd.n26196 vdd.n26194 9.3
R40316 vdd.n26168 vdd.n26166 9.3
R40317 vdd.n26190 vdd.n26187 9.3
R40318 vdd.n26591 vdd.n26588 9.3
R40319 vdd.n26598 vdd.n26596 9.3
R40320 vdd.n26612 vdd.n26603 9.3
R40321 vdd.n26686 vdd.n26675 9.3
R40322 vdd.n26680 vdd.n26678 9.3
R40323 vdd.n26291 vdd.n26288 9.3
R40324 vdd.n26330 vdd.n26327 9.3
R40325 vdd.n26334 vdd.n26332 9.3
R40326 vdd.n26402 vdd.n26399 9.3
R40327 vdd.n31767 vdd.n31764 9.3
R40328 vdd.n31811 vdd.n31809 9.3
R40329 vdd.n31819 vdd.n31816 9.3
R40330 vdd.n31855 vdd.n31853 9.3
R40331 vdd.n31863 vdd.n31860 9.3
R40332 vdd.n31897 vdd.n31895 9.3
R40333 vdd.n31905 vdd.n31902 9.3
R40334 vdd.n31962 vdd.n31960 9.3
R40335 vdd.n31972 vdd.n31969 9.3
R40336 vdd.n31986 vdd.n31983 9.3
R40337 vdd.n31991 vdd.n31989 9.3
R40338 vdd.n32001 vdd.n31998 9.3
R40339 vdd.n31609 vdd.n31606 9.3
R40340 vdd.n32022 vdd.n32020 9.3
R40341 vdd.n32034 vdd.n31604 9.3
R40342 vdd.n32047 vdd.n31591 9.3
R40343 vdd.n32053 vdd.n32051 9.3
R40344 vdd.n32084 vdd.n32081 9.3
R40345 vdd.n32116 vdd.n32113 9.3
R40346 vdd.n32169 vdd.n32167 9.3
R40347 vdd.n32177 vdd.n32174 9.3
R40348 vdd.n32213 vdd.n32211 9.3
R40349 vdd.n32221 vdd.n32218 9.3
R40350 vdd.n32262 vdd.n32260 9.3
R40351 vdd.n32270 vdd.n32267 9.3
R40352 vdd.n32318 vdd.n32316 9.3
R40353 vdd.n32328 vdd.n32325 9.3
R40354 vdd.n32345 vdd.n32342 9.3
R40355 vdd.n32351 vdd.n32349 9.3
R40356 vdd.n31468 vdd.n31465 9.3
R40357 vdd.n32375 vdd.n32373 9.3
R40358 vdd.n32381 vdd.n32379 9.3
R40359 vdd.n31446 vdd.n31443 9.3
R40360 vdd.n32523 vdd.n32410 9.3
R40361 vdd.n32515 vdd.n32412 9.3
R40362 vdd.n32495 vdd.n32415 9.3
R40363 vdd.n32471 vdd.n32424 9.3
R40364 vdd.n31055 vdd.n31053 9.3
R40365 vdd.n31063 vdd.n31060 9.3
R40366 vdd.n31107 vdd.n31105 9.3
R40367 vdd.n31115 vdd.n31112 9.3
R40368 vdd.n26193 vdd.n26192 9.3
R40369 vdd.n26595 vdd.n26594 9.3
R40370 vdd.n26608 vdd.n26607 9.3
R40371 vdd.n26682 vdd.n26681 9.3
R40372 vdd.n26296 vdd.n26295 9.3
R40373 vdd.n26336 vdd.n26335 9.3
R40374 vdd.n31794 vdd.n31793 9.3
R40375 vdd.n31814 vdd.n31813 9.3
R40376 vdd.n31833 vdd.n31832 9.3
R40377 vdd.n31858 vdd.n31857 9.3
R40378 vdd.n31875 vdd.n31874 9.3
R40379 vdd.n31900 vdd.n31899 9.3
R40380 vdd.n31973 vdd.n31644 9.3
R40381 vdd.n31988 vdd.n31632 9.3
R40382 vdd.n32007 vdd.n32006 9.3
R40383 vdd.n32019 vdd.n32018 9.3
R40384 vdd.n32037 vdd.n32036 9.3
R40385 vdd.n32050 vdd.n32049 9.3
R40386 vdd.n32144 vdd.n32143 9.3
R40387 vdd.n32172 vdd.n32171 9.3
R40388 vdd.n32194 vdd.n32193 9.3
R40389 vdd.n32216 vdd.n32215 9.3
R40390 vdd.n32248 vdd.n32247 9.3
R40391 vdd.n32265 vdd.n32264 9.3
R40392 vdd.n32331 vdd.n31492 9.3
R40393 vdd.n32348 vdd.n31476 9.3
R40394 vdd.n32362 vdd.n32361 9.3
R40395 vdd.n32378 vdd.n32377 9.3
R40396 vdd.n32533 vdd.n32532 9.3
R40397 vdd.n32517 vdd.n32516 9.3
R40398 vdd.n32459 vdd.n32458 9.3
R40399 vdd.n31058 vdd.n31057 9.3
R40400 vdd.n31081 vdd.n31080 9.3
R40401 vdd.n31110 vdd.n31109 9.3
R40402 vdd.n31186 vdd.n31185 9.3
R40403 vdd.n31184 vdd.n31183 9.3
R40404 vdd.n31124 vdd.n31123 9.3
R40405 vdd.n31086 vdd.n31085 9.3
R40406 vdd.n31078 vdd.n31077 9.3
R40407 vdd.n32457 vdd.n32456 9.3
R40408 vdd.n32461 vdd.n32460 9.3
R40409 vdd.n32531 vdd.n32530 9.3
R40410 vdd.n32365 vdd.n32364 9.3
R40411 vdd.n32334 vdd.n32333 9.3
R40412 vdd.n32287 vdd.n32286 9.3
R40413 vdd.n32253 vdd.n32252 9.3
R40414 vdd.n32236 vdd.n32235 9.3
R40415 vdd.n32199 vdd.n32198 9.3
R40416 vdd.n32191 vdd.n32190 9.3
R40417 vdd.n32149 vdd.n32148 9.3
R40418 vdd.n32141 vdd.n32140 9.3
R40419 vdd.n32040 vdd.n32039 9.3
R40420 vdd.n32010 vdd.n32009 9.3
R40421 vdd.n31976 vdd.n31975 9.3
R40422 vdd.n31915 vdd.n31914 9.3
R40423 vdd.n31880 vdd.n31879 9.3
R40424 vdd.n31872 vdd.n31871 9.3
R40425 vdd.n31838 vdd.n31837 9.3
R40426 vdd.n31830 vdd.n31829 9.3
R40427 vdd.n31799 vdd.n31798 9.3
R40428 vdd.n31791 vdd.n31790 9.3
R40429 vdd.n26316 vdd.n26315 9.3
R40430 vdd.n26690 vdd.n26689 9.3
R40431 vdd.n26196 vdd.n26195 9.3
R40432 vdd.n26168 vdd.n26167 9.3
R40433 vdd.n26190 vdd.n26189 9.3
R40434 vdd.n26591 vdd.n26590 9.3
R40435 vdd.n26598 vdd.n26597 9.3
R40436 vdd.n26612 vdd.n26611 9.3
R40437 vdd.n26686 vdd.n26685 9.3
R40438 vdd.n26680 vdd.n26679 9.3
R40439 vdd.n26291 vdd.n26290 9.3
R40440 vdd.n26330 vdd.n26329 9.3
R40441 vdd.n26334 vdd.n26333 9.3
R40442 vdd.n26402 vdd.n26401 9.3
R40443 vdd.n31767 vdd.n31766 9.3
R40444 vdd.n31811 vdd.n31810 9.3
R40445 vdd.n31819 vdd.n31818 9.3
R40446 vdd.n31855 vdd.n31854 9.3
R40447 vdd.n31863 vdd.n31862 9.3
R40448 vdd.n31897 vdd.n31896 9.3
R40449 vdd.n31905 vdd.n31904 9.3
R40450 vdd.n31962 vdd.n31961 9.3
R40451 vdd.n31972 vdd.n31971 9.3
R40452 vdd.n31986 vdd.n31985 9.3
R40453 vdd.n31991 vdd.n31990 9.3
R40454 vdd.n32001 vdd.n32000 9.3
R40455 vdd.n31609 vdd.n31608 9.3
R40456 vdd.n32022 vdd.n32021 9.3
R40457 vdd.n32034 vdd.n31602 9.3
R40458 vdd.n32047 vdd.n31589 9.3
R40459 vdd.n32053 vdd.n32052 9.3
R40460 vdd.n32084 vdd.n32083 9.3
R40461 vdd.n32116 vdd.n32115 9.3
R40462 vdd.n32169 vdd.n32168 9.3
R40463 vdd.n32177 vdd.n32176 9.3
R40464 vdd.n32213 vdd.n32212 9.3
R40465 vdd.n32221 vdd.n32220 9.3
R40466 vdd.n32262 vdd.n32261 9.3
R40467 vdd.n32270 vdd.n32269 9.3
R40468 vdd.n32318 vdd.n32317 9.3
R40469 vdd.n32328 vdd.n32327 9.3
R40470 vdd.n32345 vdd.n32344 9.3
R40471 vdd.n32351 vdd.n32350 9.3
R40472 vdd.n31468 vdd.n31467 9.3
R40473 vdd.n32375 vdd.n32371 9.3
R40474 vdd.n32381 vdd.n32380 9.3
R40475 vdd.n31446 vdd.n31445 9.3
R40476 vdd.n32523 vdd.n32522 9.3
R40477 vdd.n32515 vdd.n32514 9.3
R40478 vdd.n32495 vdd.n32494 9.3
R40479 vdd.n32471 vdd.n32470 9.3
R40480 vdd.n31055 vdd.n31054 9.3
R40481 vdd.n31063 vdd.n31062 9.3
R40482 vdd.n31107 vdd.n31106 9.3
R40483 vdd.n31115 vdd.n31114 9.3
R40484 vdd.n31071 vdd.n31048 9.3
R40485 vdd.n31048 vdd.n31047 9.3
R40486 vdd.n32468 vdd.n32432 9.3
R40487 vdd.n32432 vdd.n32431 9.3
R40488 vdd.n32507 vdd.n32506 9.3
R40489 vdd.n32506 vdd.n32505 9.3
R40490 vdd.n32502 vdd.n32501 9.3
R40491 vdd.n32353 vdd.n32352 9.3
R40492 vdd.n32320 vdd.n32319 9.3
R40493 vdd.n32204 vdd.n32203 9.3
R40494 vdd.n32203 vdd.n32202 9.3
R40495 vdd.n32158 vdd.n32157 9.3
R40496 vdd.n32157 vdd.n32156 9.3
R40497 vdd.n32098 vdd.n32097 9.3
R40498 vdd.n31599 vdd.n31598 9.3
R40499 vdd.n31978 vdd.n31977 9.3
R40500 vdd.n31953 vdd.n31952 9.3
R40501 vdd.n31868 vdd.n31867 9.3
R40502 vdd.n31867 vdd.n31866 9.3
R40503 vdd.n31824 vdd.n31823 9.3
R40504 vdd.n31823 vdd.n31822 9.3
R40505 vdd.n31774 vdd.n31773 9.3
R40506 vdd.n26348 vdd.n26347 9.3
R40507 vdd.n26347 vdd.n26346 9.3
R40508 vdd.n26343 vdd.n26342 9.3
R40509 vdd.n26600 vdd.n26599 9.3
R40510 vdd.n27238 vdd.n27237 9.3
R40511 vdd.n27237 vdd.n27236 9.3
R40512 vdd.n26178 vdd.n26177 9.3
R40513 vdd.n26177 vdd.n26176 9.3
R40514 vdd.n26198 vdd.n26197 9.3
R40515 vdd.n26213 vdd.n26212 9.3
R40516 vdd.n26212 vdd.n26211 9.3
R40517 vdd.n26211 vdd.n26210 9.3
R40518 vdd.n26620 vdd.n26619 9.3
R40519 vdd.n26619 vdd.n26618 9.3
R40520 vdd.n26703 vdd.n26702 9.3
R40521 vdd.n26702 vdd.n26701 9.3
R40522 vdd.n26312 vdd.n26311 9.3
R40523 vdd.n26311 vdd.n26310 9.3
R40524 vdd.n31758 vdd.n31757 9.3
R40525 vdd.n31757 vdd.n31756 9.3
R40526 vdd.n31756 vdd.n31755 9.3
R40527 vdd.n31804 vdd.n31803 9.3
R40528 vdd.n31803 vdd.n31802 9.3
R40529 vdd.n31849 vdd.n31848 9.3
R40530 vdd.n31848 vdd.n31847 9.3
R40531 vdd.n31847 vdd.n31846 9.3
R40532 vdd.n31894 vdd.n31893 9.3
R40533 vdd.n31893 vdd.n31892 9.3
R40534 vdd.n31892 vdd.n31891 9.3
R40535 vdd.n31912 vdd.n31911 9.3
R40536 vdd.n31911 vdd.n31910 9.3
R40537 vdd.n31939 vdd.n31674 9.3
R40538 vdd.n31674 vdd.n31673 9.3
R40539 vdd.n31954 vdd.n31668 9.3
R40540 vdd.n31668 vdd.n31667 9.3
R40541 vdd.n31964 vdd.n31963 9.3
R40542 vdd.n31967 vdd.n31660 9.3
R40543 vdd.n31660 vdd.n31659 9.3
R40544 vdd.n31659 vdd.n31658 9.3
R40545 vdd.n31981 vdd.n31642 9.3
R40546 vdd.n31642 vdd.n31641 9.3
R40547 vdd.n31993 vdd.n31992 9.3
R40548 vdd.n31996 vdd.n31631 9.3
R40549 vdd.n31631 vdd.n31630 9.3
R40550 vdd.n31630 vdd.n31629 9.3
R40551 vdd.n31615 vdd.n31614 9.3
R40552 vdd.n32069 vdd.n32068 9.3
R40553 vdd.n32068 vdd.n32067 9.3
R40554 vdd.n32124 vdd.n32123 9.3
R40555 vdd.n32123 vdd.n32122 9.3
R40556 vdd.n32185 vdd.n31574 9.3
R40557 vdd.n31574 vdd.n31573 9.3
R40558 vdd.n31573 vdd.n31572 9.3
R40559 vdd.n32232 vdd.n32231 9.3
R40560 vdd.n32231 vdd.n32230 9.3
R40561 vdd.n32230 vdd.n32229 9.3
R40562 vdd.n32259 vdd.n32258 9.3
R40563 vdd.n32258 vdd.n32257 9.3
R40564 vdd.n32284 vdd.n32283 9.3
R40565 vdd.n32283 vdd.n32282 9.3
R40566 vdd.n31524 vdd.n31523 9.3
R40567 vdd.n31514 vdd.n31513 9.3
R40568 vdd.n31513 vdd.n31512 9.3
R40569 vdd.n32323 vdd.n31500 9.3
R40570 vdd.n31500 vdd.n31499 9.3
R40571 vdd.n32336 vdd.n32335 9.3
R40572 vdd.n32340 vdd.n31490 9.3
R40573 vdd.n31490 vdd.n31489 9.3
R40574 vdd.n31489 vdd.n31488 9.3
R40575 vdd.n32356 vdd.n31475 9.3
R40576 vdd.n31475 vdd.n31474 9.3
R40577 vdd.n31462 vdd.n31461 9.3
R40578 vdd.n31461 vdd.n31460 9.3
R40579 vdd.n32405 vdd.n32404 9.3
R40580 vdd.n32404 vdd.n32403 9.3
R40581 vdd.n32498 vdd.n32497 9.3
R40582 vdd.n32486 vdd.n32485 9.3
R40583 vdd.n32485 vdd.n32484 9.3
R40584 vdd.n32476 vdd.n32475 9.3
R40585 vdd.n32465 vdd.n32464 9.3
R40586 vdd.n32449 vdd.n32448 9.3
R40587 vdd.n32448 vdd.n32447 9.3
R40588 vdd.n31097 vdd.n31096 9.3
R40589 vdd.n31096 vdd.n31095 9.3
R40590 vdd.n31095 vdd.n31094 9.3
R40591 vdd.n31120 vdd.n31119 9.3
R40592 vdd.n31119 vdd.n31118 9.3
R40593 vdd.n31180 vdd.n31179 9.3
R40594 vdd.n31179 vdd.n31178 9.3
R40595 vdd.n12571 vdd.n10268 9.3
R40596 vdd.n10490 vdd.n10257 9.3
R40597 vdd.n10261 vdd.n10256 9.3
R40598 vdd.n12581 vdd.n10123 9.3
R40599 vdd.n12584 vdd.n12583 9.3
R40600 vdd.n10248 vdd.n10247 9.3
R40601 vdd.n10227 vdd.n10226 9.3
R40602 vdd.n10231 vdd.n10069 9.3
R40603 vdd.n10234 vdd.n10233 9.3
R40604 vdd.n10098 vdd.n10070 9.3
R40605 vdd.n10096 vdd.n10076 9.3
R40606 vdd.n12600 vdd.n12599 9.3
R40607 vdd.n12601 vdd.n12600 9.3
R40608 vdd.n10199 vdd.n10065 9.3
R40609 vdd.n12600 vdd.n10090 9.3
R40610 vdd.n10195 vdd.n10194 9.3
R40611 vdd.n12600 vdd.n10086 9.3
R40612 vdd.n11476 vdd.n11475 9.3
R40613 vdd.n11992 vdd.n11991 9.3
R40614 vdd.n11996 vdd.n11402 9.3
R40615 vdd.n12007 vdd.n12006 9.3
R40616 vdd.n11398 vdd.n11381 9.3
R40617 vdd.n11388 vdd.n11387 9.3
R40618 vdd.n12023 vdd.n12022 9.3
R40619 vdd.n11360 vdd.n11337 9.3
R40620 vdd.n11347 vdd.n11346 9.3
R40621 vdd.n11345 vdd.n11344 9.3
R40622 vdd.n12041 vdd.n11318 9.3
R40623 vdd.n12052 vdd.n12051 9.3
R40624 vdd.n11312 vdd.n11311 9.3
R40625 vdd.n11302 vdd.n11301 9.3
R40626 vdd.n11295 vdd.n11294 9.3
R40627 vdd.n12080 vdd.n12079 9.3
R40628 vdd.n11263 vdd.n11246 9.3
R40629 vdd.n11253 vdd.n11252 9.3
R40630 vdd.n12096 vdd.n12095 9.3
R40631 vdd.n12100 vdd.n11218 9.3
R40632 vdd.n12111 vdd.n12110 9.3
R40633 vdd.n11214 vdd.n11197 9.3
R40634 vdd.n11204 vdd.n11203 9.3
R40635 vdd.n12127 vdd.n11179 9.3
R40636 vdd.n12138 vdd.n12137 9.3
R40637 vdd.n11174 vdd.n11173 9.3
R40638 vdd.n11165 vdd.n11164 9.3
R40639 vdd.n11158 vdd.n11157 9.3
R40640 vdd.n12156 vdd.n11130 9.3
R40641 vdd.n12167 vdd.n12166 9.3
R40642 vdd.n11124 vdd.n11123 9.3
R40643 vdd.n12184 vdd.n12183 9.3
R40644 vdd.n12188 vdd.n11083 9.3
R40645 vdd.n12199 vdd.n12198 9.3
R40646 vdd.n11079 vdd.n11062 9.3
R40647 vdd.n11069 vdd.n11068 9.3
R40648 vdd.n12215 vdd.n12214 9.3
R40649 vdd.n12219 vdd.n11034 9.3
R40650 vdd.n12230 vdd.n12229 9.3
R40651 vdd.n11018 vdd.n11017 9.3
R40652 vdd.n11023 vdd.n11022 9.3
R40653 vdd.n12246 vdd.n10996 9.3
R40654 vdd.n12257 vdd.n12256 9.3
R40655 vdd.n10990 vdd.n10989 9.3
R40656 vdd.n10980 vdd.n10979 9.3
R40657 vdd.n10973 vdd.n10972 9.3
R40658 vdd.n10949 vdd.n10924 9.3
R40659 vdd.n10942 vdd.n10926 9.3
R40660 vdd.n10932 vdd.n10931 9.3
R40661 vdd.n12298 vdd.n12297 9.3
R40662 vdd.n12302 vdd.n10893 9.3
R40663 vdd.n12313 vdd.n12312 9.3
R40664 vdd.n10889 vdd.n10872 9.3
R40665 vdd.n10879 vdd.n10878 9.3
R40666 vdd.n12329 vdd.n12328 9.3
R40667 vdd.n10851 vdd.n10828 9.3
R40668 vdd.n10838 vdd.n10837 9.3
R40669 vdd.n10836 vdd.n10835 9.3
R40670 vdd.n12347 vdd.n10809 9.3
R40671 vdd.n12358 vdd.n12357 9.3
R40672 vdd.n10803 vdd.n10802 9.3
R40673 vdd.n10793 vdd.n10792 9.3
R40674 vdd.n10786 vdd.n10785 9.3
R40675 vdd.n12379 vdd.n10746 9.3
R40676 vdd.n12390 vdd.n12389 9.3
R40677 vdd.n10742 vdd.n10725 9.3
R40678 vdd.n10732 vdd.n10731 9.3
R40679 vdd.n12406 vdd.n12405 9.3
R40680 vdd.n12410 vdd.n10697 9.3
R40681 vdd.n12421 vdd.n12420 9.3
R40682 vdd.n10693 vdd.n10677 9.3
R40683 vdd.n10683 vdd.n10682 9.3
R40684 vdd.n12436 vdd.n10658 9.3
R40685 vdd.n12447 vdd.n12446 9.3
R40686 vdd.n10652 vdd.n10651 9.3
R40687 vdd.n10642 vdd.n10641 9.3
R40688 vdd.n10635 vdd.n10634 9.3
R40689 vdd.n12465 vdd.n10607 9.3
R40690 vdd.n12476 vdd.n12475 9.3
R40691 vdd.n10593 vdd.n10592 9.3
R40692 vdd.n12494 vdd.n12493 9.3
R40693 vdd.n12498 vdd.n10561 9.3
R40694 vdd.n12509 vdd.n12508 9.3
R40695 vdd.n10557 vdd.n10534 9.3
R40696 vdd.n10547 vdd.n10546 9.3
R40697 vdd.n10540 vdd.n10521 9.3
R40698 vdd.n11519 vdd.n11518 9.3
R40699 vdd.n11597 vdd.n11596 9.3
R40700 vdd.n11937 vdd.n11554 9.3
R40701 vdd.n11536 vdd.n11453 9.3
R40702 vdd.n11517 vdd.n11461 9.3
R40703 vdd.n11464 vdd.n11433 9.3
R40704 vdd.n11487 vdd.n11486 9.3
R40705 vdd.n11553 vdd.n11551 9.3
R40706 vdd.n11503 vdd.n11434 9.3
R40707 vdd.n11520 vdd.n11459 9.3
R40708 vdd.n11546 vdd.n11543 9.3
R40709 vdd.n11940 vdd.n11552 9.3
R40710 vdd.n9263 vdd.n9262 9.3
R40711 vdd.n11578 vdd.n9276 9.3
R40712 vdd.n8790 vdd.n8789 9.3
R40713 vdd.n13750 vdd.n8788 9.3
R40714 vdd.n13797 vdd.n8758 9.3
R40715 vdd.n8743 vdd.n8742 9.3
R40716 vdd.n13816 vdd.n13815 9.3
R40717 vdd.n8705 vdd.n8704 9.3
R40718 vdd.n8701 vdd.n8700 9.3
R40719 vdd.n13884 vdd.n8699 9.3
R40720 vdd.n13922 vdd.n8650 9.3
R40721 vdd.n8639 vdd.n8638 9.3
R40722 vdd.n13942 vdd.n8636 9.3
R40723 vdd.n13956 vdd.n8635 9.3
R40724 vdd.n8586 vdd.n8585 9.3
R40725 vdd.n14016 vdd.n8584 9.3
R40726 vdd.n14028 vdd.n8578 9.3
R40727 vdd.n14032 vdd.n14029 9.3
R40728 vdd.n14084 vdd.n8545 9.3
R40729 vdd.n8530 vdd.n8529 9.3
R40730 vdd.n14103 vdd.n14102 9.3
R40731 vdd.n8482 vdd.n8481 9.3
R40732 vdd.n8478 vdd.n8477 9.3
R40733 vdd.n14173 vdd.n8476 9.3
R40734 vdd.n14212 vdd.n8430 9.3
R40735 vdd.n8417 vdd.n8416 9.3
R40736 vdd.n14232 vdd.n8414 9.3
R40737 vdd.n14246 vdd.n8413 9.3
R40738 vdd.n8366 vdd.n8365 9.3
R40739 vdd.n8362 vdd.n8361 9.3
R40740 vdd.n14314 vdd.n8360 9.3
R40741 vdd.n14366 vdd.n8322 9.3
R40742 vdd.n8329 vdd.n8328 9.3
R40743 vdd.n14387 vdd.n8307 9.3
R40744 vdd.n8293 vdd.n8292 9.3
R40745 vdd.n8267 vdd.n8266 9.3
R40746 vdd.n14447 vdd.n8265 9.3
R40747 vdd.n14473 vdd.n14472 9.3
R40748 vdd.n14476 vdd.n8228 9.3
R40749 vdd.n14534 vdd.n8193 9.3
R40750 vdd.n14554 vdd.n8192 9.3
R40751 vdd.n14544 vdd.n14543 9.3
R40752 vdd.n14610 vdd.n14609 9.3
R40753 vdd.n14610 vdd.n8175 9.3
R40754 vdd.n8175 vdd.n8172 9.3
R40755 vdd.n14606 vdd.n14605 9.3
R40756 vdd.n14605 vdd.n14604 9.3
R40757 vdd.n14604 vdd.n14603 9.3
R40758 vdd.n14542 vdd.n8178 9.3
R40759 vdd.n14545 vdd.n14537 9.3
R40760 vdd.n14546 vdd.n14545 9.3
R40761 vdd.n14547 vdd.n14546 9.3
R40762 vdd.n14553 vdd.n14552 9.3
R40763 vdd.n14556 vdd.n14555 9.3
R40764 vdd.n14556 vdd.n8190 9.3
R40765 vdd.n8190 vdd.n8188 9.3
R40766 vdd.n14536 vdd.n14535 9.3
R40767 vdd.n14533 vdd.n8195 9.3
R40768 vdd.n14533 vdd.n14532 9.3
R40769 vdd.n14532 vdd.n14531 9.3
R40770 vdd.n14478 vdd.n14477 9.3
R40771 vdd.n14483 vdd.n14475 9.3
R40772 vdd.n14483 vdd.n14482 9.3
R40773 vdd.n14482 vdd.n8215 9.3
R40774 vdd.n14474 vdd.n8227 9.3
R40775 vdd.n14471 vdd.n8229 9.3
R40776 vdd.n14471 vdd.n8225 9.3
R40777 vdd.n8233 vdd.n8225 9.3
R40778 vdd.n14446 vdd.n14445 9.3
R40779 vdd.n14449 vdd.n14448 9.3
R40780 vdd.n14450 vdd.n14449 9.3
R40781 vdd.n14451 vdd.n14450 9.3
R40782 vdd.n14444 vdd.n14443 9.3
R40783 vdd.n14415 vdd.n14414 9.3
R40784 vdd.n14414 vdd.n8268 9.3
R40785 vdd.n8268 vdd.n8241 9.3
R40786 vdd.n14412 vdd.n14411 9.3
R40787 vdd.n14411 vdd.n14410 9.3
R40788 vdd.n14410 vdd.n14409 9.3
R40789 vdd.n14390 vdd.n14389 9.3
R40790 vdd.n14392 vdd.n14391 9.3
R40791 vdd.n14393 vdd.n14392 9.3
R40792 vdd.n14394 vdd.n14393 9.3
R40793 vdd.n14386 vdd.n14385 9.3
R40794 vdd.n8310 vdd.n8309 9.3
R40795 vdd.n8311 vdd.n8310 9.3
R40796 vdd.n8312 vdd.n8311 9.3
R40797 vdd.n8330 vdd.n8324 9.3
R40798 vdd.n14365 vdd.n14364 9.3
R40799 vdd.n14364 vdd.n14363 9.3
R40800 vdd.n14363 vdd.n14362 9.3
R40801 vdd.n14368 vdd.n14367 9.3
R40802 vdd.n8323 vdd.n8321 9.3
R40803 vdd.n8321 vdd.n8319 9.3
R40804 vdd.n8319 vdd.n8317 9.3
R40805 vdd.n14316 vdd.n14315 9.3
R40806 vdd.n14313 vdd.n14312 9.3
R40807 vdd.n14312 vdd.n14311 9.3
R40808 vdd.n14311 vdd.n14310 9.3
R40809 vdd.n14307 vdd.n14306 9.3
R40810 vdd.n14305 vdd.n14304 9.3
R40811 vdd.n14304 vdd.n14303 9.3
R40812 vdd.n14303 vdd.n14302 9.3
R40813 vdd.n14289 vdd.n14288 9.3
R40814 vdd.n14291 vdd.n14290 9.3
R40815 vdd.n14291 vdd.n8374 9.3
R40816 vdd.n8377 vdd.n8374 9.3
R40817 vdd.n14240 vdd.n14239 9.3
R40818 vdd.n14240 vdd.n8373 9.3
R40819 vdd.n14265 vdd.n8373 9.3
R40820 vdd.n14245 vdd.n14244 9.3
R40821 vdd.n14248 vdd.n14247 9.3
R40822 vdd.n14249 vdd.n14248 9.3
R40823 vdd.n14250 vdd.n14249 9.3
R40824 vdd.n14237 vdd.n14236 9.3
R40825 vdd.n14231 vdd.n14230 9.3
R40826 vdd.n14231 vdd.n8398 9.3
R40827 vdd.n14257 vdd.n8398 9.3
R40828 vdd.n14229 vdd.n14228 9.3
R40829 vdd.n8433 vdd.n8432 9.3
R40830 vdd.n8433 vdd.n8418 9.3
R40831 vdd.n8436 vdd.n8418 9.3
R40832 vdd.n14211 vdd.n14210 9.3
R40833 vdd.n14214 vdd.n14213 9.3
R40834 vdd.n14214 vdd.n8428 9.3
R40835 vdd.n8453 vdd.n8428 9.3
R40836 vdd.n8475 vdd.n8431 9.3
R40837 vdd.n14175 vdd.n14174 9.3
R40838 vdd.n14176 vdd.n14175 9.3
R40839 vdd.n14177 vdd.n14176 9.3
R40840 vdd.n14172 vdd.n14171 9.3
R40841 vdd.n14166 vdd.n14165 9.3
R40842 vdd.n14167 vdd.n14166 9.3
R40843 vdd.n14167 vdd.n8457 9.3
R40844 vdd.n14164 vdd.n14163 9.3
R40845 vdd.n14149 vdd.n14148 9.3
R40846 vdd.n14148 vdd.n8483 9.3
R40847 vdd.n8497 vdd.n8483 9.3
R40848 vdd.n14105 vdd.n8495 9.3
R40849 vdd.n14106 vdd.n14105 9.3
R40850 vdd.n14107 vdd.n14106 9.3
R40851 vdd.n14101 vdd.n8528 9.3
R40852 vdd.n14100 vdd.n14099 9.3
R40853 vdd.n14099 vdd.n14098 9.3
R40854 vdd.n14098 vdd.n14097 9.3
R40855 vdd.n8548 vdd.n8547 9.3
R40856 vdd.n14083 vdd.n14082 9.3
R40857 vdd.n14082 vdd.n14081 9.3
R40858 vdd.n14081 vdd.n14080 9.3
R40859 vdd.n14086 vdd.n14085 9.3
R40860 vdd.n8546 vdd.n8544 9.3
R40861 vdd.n8544 vdd.n8542 9.3
R40862 vdd.n8542 vdd.n8540 9.3
R40863 vdd.n14034 vdd.n14033 9.3
R40864 vdd.n14036 vdd.n14035 9.3
R40865 vdd.n14037 vdd.n14036 9.3
R40866 vdd.n14038 vdd.n14037 9.3
R40867 vdd.n14027 vdd.n14026 9.3
R40868 vdd.n8581 vdd.n8580 9.3
R40869 vdd.n14022 vdd.n8581 9.3
R40870 vdd.n14022 vdd.n14021 9.3
R40871 vdd.n14018 vdd.n14017 9.3
R40872 vdd.n14015 vdd.n14014 9.3
R40873 vdd.n14014 vdd.n14013 9.3
R40874 vdd.n14013 vdd.n14012 9.3
R40875 vdd.n13998 vdd.n13997 9.3
R40876 vdd.n14000 vdd.n13999 9.3
R40877 vdd.n14000 vdd.n8596 9.3
R40878 vdd.n8599 vdd.n8596 9.3
R40879 vdd.n13950 vdd.n13949 9.3
R40880 vdd.n13950 vdd.n8595 9.3
R40881 vdd.n13975 vdd.n8595 9.3
R40882 vdd.n13955 vdd.n13954 9.3
R40883 vdd.n13958 vdd.n13957 9.3
R40884 vdd.n13959 vdd.n13958 9.3
R40885 vdd.n13960 vdd.n13959 9.3
R40886 vdd.n13947 vdd.n13946 9.3
R40887 vdd.n13941 vdd.n13940 9.3
R40888 vdd.n13941 vdd.n8620 9.3
R40889 vdd.n13967 vdd.n8620 9.3
R40890 vdd.n13939 vdd.n13938 9.3
R40891 vdd.n8653 vdd.n8652 9.3
R40892 vdd.n8653 vdd.n8640 9.3
R40893 vdd.n8657 vdd.n8640 9.3
R40894 vdd.n13921 vdd.n13920 9.3
R40895 vdd.n13924 vdd.n13923 9.3
R40896 vdd.n13924 vdd.n8648 9.3
R40897 vdd.n8677 vdd.n8648 9.3
R40898 vdd.n8698 vdd.n8651 9.3
R40899 vdd.n13886 vdd.n13885 9.3
R40900 vdd.n13887 vdd.n13886 9.3
R40901 vdd.n13888 vdd.n13887 9.3
R40902 vdd.n13883 vdd.n13882 9.3
R40903 vdd.n13877 vdd.n13876 9.3
R40904 vdd.n13878 vdd.n13877 9.3
R40905 vdd.n13878 vdd.n8681 9.3
R40906 vdd.n13875 vdd.n13874 9.3
R40907 vdd.n13860 vdd.n13859 9.3
R40908 vdd.n13859 vdd.n8706 9.3
R40909 vdd.n8719 vdd.n8706 9.3
R40910 vdd.n13817 vdd.n8717 9.3
R40911 vdd.n13817 vdd.n8740 9.3
R40912 vdd.n8740 vdd.n8739 9.3
R40913 vdd.n13814 vdd.n8741 9.3
R40914 vdd.n13813 vdd.n13812 9.3
R40915 vdd.n13812 vdd.n13811 9.3
R40916 vdd.n13811 vdd.n13810 9.3
R40917 vdd.n8761 vdd.n8760 9.3
R40918 vdd.n13796 vdd.n13795 9.3
R40919 vdd.n13795 vdd.n13794 9.3
R40920 vdd.n13794 vdd.n13793 9.3
R40921 vdd.n13799 vdd.n13798 9.3
R40922 vdd.n8759 vdd.n8757 9.3
R40923 vdd.n8757 vdd.n8755 9.3
R40924 vdd.n8755 vdd.n8753 9.3
R40925 vdd.n13752 vdd.n13751 9.3
R40926 vdd.n13749 vdd.n13748 9.3
R40927 vdd.n13748 vdd.n13747 9.3
R40928 vdd.n13747 vdd.n13746 9.3
R40929 vdd.n9255 vdd.n9254 9.3
R40930 vdd.n13137 vdd.n13136 9.3
R40931 vdd.n11624 vdd.n11623 9.3
R40932 vdd.n11615 vdd.n11614 9.3
R40933 vdd.n11613 vdd.n9248 9.3
R40934 vdd.n9248 vdd.n9246 9.3
R40935 vdd.n9246 vdd.n9244 9.3
R40936 vdd.n9251 vdd.n9249 9.3
R40937 vdd.n9257 vdd.n9256 9.3
R40938 vdd.n9232 vdd.n9231 9.3
R40939 vdd.n13168 vdd.n9229 9.3
R40940 vdd.n13172 vdd.n9228 9.3
R40941 vdd.n13223 vdd.n9195 9.3
R40942 vdd.n9197 vdd.n9182 9.3
R40943 vdd.n13281 vdd.n9153 9.3
R40944 vdd.n13307 vdd.n9136 9.3
R40945 vdd.n13311 vdd.n9135 9.3
R40946 vdd.n9114 vdd.n9109 9.3
R40947 vdd.n9117 vdd.n9113 9.3
R40948 vdd.n9081 vdd.n9075 9.3
R40949 vdd.n9083 vdd.n9080 9.3
R40950 vdd.n13432 vdd.n9025 9.3
R40951 vdd.n9014 vdd.n9013 9.3
R40952 vdd.n13450 vdd.n9012 9.3
R40953 vdd.n13462 vdd.n9006 9.3
R40954 vdd.n13466 vdd.n13463 9.3
R40955 vdd.n13515 vdd.n8973 9.3
R40956 vdd.n8975 vdd.n8961 9.3
R40957 vdd.n13573 vdd.n8932 9.3
R40958 vdd.n13599 vdd.n8914 9.3
R40959 vdd.n13603 vdd.n8913 9.3
R40960 vdd.n8893 vdd.n8888 9.3
R40961 vdd.n8896 vdd.n8892 9.3
R40962 vdd.n8861 vdd.n8855 9.3
R40963 vdd.n8863 vdd.n8860 9.3
R40964 vdd.n13724 vdd.n8805 9.3
R40965 vdd.n8794 vdd.n8793 9.3
R40966 vdd.n9237 vdd.n9236 9.3
R40967 vdd.n13742 vdd.n13741 9.3
R40968 vdd.n13740 vdd.n13739 9.3
R40969 vdd.n13739 vdd.n13738 9.3
R40970 vdd.n13738 vdd.n13737 9.3
R40971 vdd.n8808 vdd.n8807 9.3
R40972 vdd.n13723 vdd.n13722 9.3
R40973 vdd.n13722 vdd.n13721 9.3
R40974 vdd.n13721 vdd.n13720 9.3
R40975 vdd.n13726 vdd.n13725 9.3
R40976 vdd.n8806 vdd.n8804 9.3
R40977 vdd.n8804 vdd.n8802 9.3
R40978 vdd.n8802 vdd.n8800 9.3
R40979 vdd.n13675 vdd.n13674 9.3
R40980 vdd.n13674 vdd.n8837 9.3
R40981 vdd.n8837 vdd.n8836 9.3
R40982 vdd.n8859 vdd.n8839 9.3
R40983 vdd.n8865 vdd.n8864 9.3
R40984 vdd.n8865 vdd.n8841 9.3
R40985 vdd.n13668 vdd.n8841 9.3
R40986 vdd.n8862 vdd.n8858 9.3
R40987 vdd.n13653 vdd.n8856 9.3
R40988 vdd.n13653 vdd.n13652 9.3
R40989 vdd.n13652 vdd.n13651 9.3
R40990 vdd.n8895 vdd.n8854 9.3
R40991 vdd.n8898 vdd.n8897 9.3
R40992 vdd.n8898 vdd.n8852 9.3
R40993 vdd.n8901 vdd.n8852 9.3
R40994 vdd.n8894 vdd.n8891 9.3
R40995 vdd.n13623 vdd.n8889 9.3
R40996 vdd.n13623 vdd.n13622 9.3
R40997 vdd.n13622 vdd.n8873 9.3
R40998 vdd.n13602 vdd.n8887 9.3
R40999 vdd.n13605 vdd.n13604 9.3
R41000 vdd.n13605 vdd.n8885 9.3
R41001 vdd.n8909 vdd.n8885 9.3
R41002 vdd.n13601 vdd.n13600 9.3
R41003 vdd.n13598 vdd.n8916 9.3
R41004 vdd.n13598 vdd.n13597 9.3
R41005 vdd.n13597 vdd.n13596 9.3
R41006 vdd.n13575 vdd.n13574 9.3
R41007 vdd.n13572 vdd.n13571 9.3
R41008 vdd.n13571 vdd.n8931 9.3
R41009 vdd.n8936 vdd.n8931 9.3
R41010 vdd.n13532 vdd.n8962 9.3
R41011 vdd.n13532 vdd.n13531 9.3
R41012 vdd.n13531 vdd.n13530 9.3
R41013 vdd.n8977 vdd.n8976 9.3
R41014 vdd.n13514 vdd.n13513 9.3
R41015 vdd.n13513 vdd.n13512 9.3
R41016 vdd.n13512 vdd.n13511 9.3
R41017 vdd.n13517 vdd.n13516 9.3
R41018 vdd.n8974 vdd.n8972 9.3
R41019 vdd.n8972 vdd.n8970 9.3
R41020 vdd.n8970 vdd.n8969 9.3
R41021 vdd.n13468 vdd.n13467 9.3
R41022 vdd.n13470 vdd.n13469 9.3
R41023 vdd.n13471 vdd.n13470 9.3
R41024 vdd.n13472 vdd.n13471 9.3
R41025 vdd.n13461 vdd.n13460 9.3
R41026 vdd.n9009 vdd.n9008 9.3
R41027 vdd.n13456 vdd.n9009 9.3
R41028 vdd.n13456 vdd.n13455 9.3
R41029 vdd.n13452 vdd.n13451 9.3
R41030 vdd.n13449 vdd.n13448 9.3
R41031 vdd.n13448 vdd.n13447 9.3
R41032 vdd.n13447 vdd.n13446 9.3
R41033 vdd.n9028 vdd.n9027 9.3
R41034 vdd.n13431 vdd.n13430 9.3
R41035 vdd.n13430 vdd.n13429 9.3
R41036 vdd.n13429 vdd.n13428 9.3
R41037 vdd.n13434 vdd.n13433 9.3
R41038 vdd.n9026 vdd.n9024 9.3
R41039 vdd.n9024 vdd.n9022 9.3
R41040 vdd.n9022 vdd.n9020 9.3
R41041 vdd.n13383 vdd.n13382 9.3
R41042 vdd.n13382 vdd.n9057 9.3
R41043 vdd.n9057 vdd.n9056 9.3
R41044 vdd.n9079 vdd.n9059 9.3
R41045 vdd.n9085 vdd.n9084 9.3
R41046 vdd.n9085 vdd.n9061 9.3
R41047 vdd.n13376 vdd.n9061 9.3
R41048 vdd.n9082 vdd.n9078 9.3
R41049 vdd.n13361 vdd.n9076 9.3
R41050 vdd.n13361 vdd.n13360 9.3
R41051 vdd.n13360 vdd.n13359 9.3
R41052 vdd.n9116 vdd.n9074 9.3
R41053 vdd.n9119 vdd.n9118 9.3
R41054 vdd.n9119 vdd.n9072 9.3
R41055 vdd.n9122 vdd.n9072 9.3
R41056 vdd.n9115 vdd.n9112 9.3
R41057 vdd.n13331 vdd.n9110 9.3
R41058 vdd.n13331 vdd.n13330 9.3
R41059 vdd.n13330 vdd.n9093 9.3
R41060 vdd.n13310 vdd.n9108 9.3
R41061 vdd.n13313 vdd.n13312 9.3
R41062 vdd.n13313 vdd.n9106 9.3
R41063 vdd.n9131 vdd.n9106 9.3
R41064 vdd.n13309 vdd.n13308 9.3
R41065 vdd.n13306 vdd.n9138 9.3
R41066 vdd.n13306 vdd.n13305 9.3
R41067 vdd.n13305 vdd.n13304 9.3
R41068 vdd.n13283 vdd.n13282 9.3
R41069 vdd.n13280 vdd.n13279 9.3
R41070 vdd.n13279 vdd.n9152 9.3
R41071 vdd.n9158 vdd.n9152 9.3
R41072 vdd.n13240 vdd.n9183 9.3
R41073 vdd.n13240 vdd.n13239 9.3
R41074 vdd.n13239 vdd.n13238 9.3
R41075 vdd.n9199 vdd.n9198 9.3
R41076 vdd.n13222 vdd.n13221 9.3
R41077 vdd.n13221 vdd.n13220 9.3
R41078 vdd.n13220 vdd.n13219 9.3
R41079 vdd.n13225 vdd.n13224 9.3
R41080 vdd.n9196 vdd.n9194 9.3
R41081 vdd.n9194 vdd.n9192 9.3
R41082 vdd.n9192 vdd.n9190 9.3
R41083 vdd.n13174 vdd.n13173 9.3
R41084 vdd.n13171 vdd.n13170 9.3
R41085 vdd.n13170 vdd.n13169 9.3
R41086 vdd.n13169 vdd.n9224 9.3
R41087 vdd.n13167 vdd.n13166 9.3
R41088 vdd.n13165 vdd.n13164 9.3
R41089 vdd.n13164 vdd.n13163 9.3
R41090 vdd.n13163 vdd.n13162 9.3
R41091 vdd.n13158 vdd.n13157 9.3
R41092 vdd.n13156 vdd.n13155 9.3
R41093 vdd.n13155 vdd.n13154 9.3
R41094 vdd.n13154 vdd.n13153 9.3
R41095 vdd.n9259 vdd.n9258 9.3
R41096 vdd.n10082 vdd.n10081 9.3
R41097 vdd.n10183 vdd.n10182 9.3
R41098 vdd.n12600 vdd.n10080 9.3
R41099 vdd.n12623 vdd.n12622 9.3
R41100 vdd.n10170 vdd.n10145 9.3
R41101 vdd.n10163 vdd.n10162 9.3
R41102 vdd.n12638 vdd.n10031 9.3
R41103 vdd.n10024 vdd.n10023 9.3
R41104 vdd.n10001 vdd.n10000 9.3
R41105 vdd.n9961 vdd.n9960 9.3
R41106 vdd.n9944 vdd.n9918 9.3
R41107 vdd.n12716 vdd.n12715 9.3
R41108 vdd.n9894 vdd.n9893 9.3
R41109 vdd.n12732 vdd.n12731 9.3
R41110 vdd.n9865 vdd.n9838 9.3
R41111 vdd.n9849 vdd.n9848 9.3
R41112 vdd.n12770 vdd.n12769 9.3
R41113 vdd.n9787 vdd.n9764 9.3
R41114 vdd.n12811 vdd.n12810 9.3
R41115 vdd.n9740 vdd.n9739 9.3
R41116 vdd.n12831 vdd.n12830 9.3
R41117 vdd.n9709 vdd.n9708 9.3
R41118 vdd.n12846 vdd.n9671 9.3
R41119 vdd.n9664 vdd.n9663 9.3
R41120 vdd.n9641 vdd.n9640 9.3
R41121 vdd.n9601 vdd.n9600 9.3
R41122 vdd.n9584 vdd.n9559 9.3
R41123 vdd.n12924 vdd.n12923 9.3
R41124 vdd.n9533 vdd.n9532 9.3
R41125 vdd.n12940 vdd.n12939 9.3
R41126 vdd.n9505 vdd.n9478 9.3
R41127 vdd.n9489 vdd.n9488 9.3
R41128 vdd.n12978 vdd.n12977 9.3
R41129 vdd.n9427 vdd.n9404 9.3
R41130 vdd.n13019 vdd.n13018 9.3
R41131 vdd.n9380 vdd.n9379 9.3
R41132 vdd.n13039 vdd.n13038 9.3
R41133 vdd.n9349 vdd.n9348 9.3
R41134 vdd.n13054 vdd.n9310 9.3
R41135 vdd.n9304 vdd.n9303 9.3
R41136 vdd.n10361 vdd.n10360 9.3
R41137 vdd.n10399 vdd.n10398 9.3
R41138 vdd.n10412 vdd.n10411 9.3
R41139 vdd.n10426 vdd.n10304 9.3
R41140 vdd.n10295 vdd.n10293 9.3
R41141 vdd.n10448 vdd.n10292 9.3
R41142 vdd.n10286 vdd.n10285 9.3
R41143 vdd.n12620 vdd.n12619 9.3
R41144 vdd.n10172 vdd.n10171 9.3
R41145 vdd.n12621 vdd.n10051 9.3
R41146 vdd.n10150 vdd.n10149 9.3
R41147 vdd.n12649 vdd.n12648 9.3
R41148 vdd.n10015 vdd.n9985 9.3
R41149 vdd.n9999 vdd.n9998 9.3
R41150 vdd.n12686 vdd.n12685 9.3
R41151 vdd.n9950 vdd.n9949 9.3
R41152 vdd.n12706 vdd.n12705 9.3
R41153 vdd.n9906 vdd.n9905 9.3
R41154 vdd.n9874 vdd.n9873 9.3
R41155 vdd.n9851 vdd.n9850 9.3
R41156 vdd.n12759 vdd.n9817 9.3
R41157 vdd.n9809 vdd.n9808 9.3
R41158 vdd.n9805 vdd.n9804 9.3
R41159 vdd.n12801 vdd.n12800 9.3
R41160 vdd.n9751 vdd.n9750 9.3
R41161 vdd.n9733 vdd.n9711 9.3
R41162 vdd.n9698 vdd.n9697 9.3
R41163 vdd.n12857 vdd.n12856 9.3
R41164 vdd.n9655 vdd.n9625 9.3
R41165 vdd.n9639 vdd.n9638 9.3
R41166 vdd.n12894 vdd.n12893 9.3
R41167 vdd.n9590 vdd.n9589 9.3
R41168 vdd.n12914 vdd.n12913 9.3
R41169 vdd.n9546 vdd.n9545 9.3
R41170 vdd.n9514 vdd.n9513 9.3
R41171 vdd.n9491 vdd.n9490 9.3
R41172 vdd.n12967 vdd.n9457 9.3
R41173 vdd.n9450 vdd.n9449 9.3
R41174 vdd.n9446 vdd.n9445 9.3
R41175 vdd.n13009 vdd.n13008 9.3
R41176 vdd.n9391 vdd.n9390 9.3
R41177 vdd.n9373 vdd.n9351 9.3
R41178 vdd.n9338 vdd.n9337 9.3
R41179 vdd.n13065 vdd.n13064 9.3
R41180 vdd.n10362 vdd.n9293 9.3
R41181 vdd.n10375 vdd.n10374 9.3
R41182 vdd.n10348 vdd.n10347 9.3
R41183 vdd.n10328 vdd.n10323 9.3
R41184 vdd.n10422 vdd.n10421 9.3
R41185 vdd.n10437 vdd.n10436 9.3
R41186 vdd.n10459 vdd.n10458 9.3
R41187 vdd.n10164 vdd.n10147 9.3
R41188 vdd.n10161 vdd.n10148 9.3
R41189 vdd.n10396 vdd.n10335 9.3
R41190 vdd.n10396 vdd.n10395 9.3
R41191 vdd.n10395 vdd.n10394 9.3
R41192 vdd.n10401 vdd.n10400 9.3
R41193 vdd.n10402 vdd.n10401 9.3
R41194 vdd.n10403 vdd.n10402 9.3
R41195 vdd.n10409 vdd.n10408 9.3
R41196 vdd.n10408 vdd.n10321 9.3
R41197 vdd.n10321 vdd.n10320 9.3
R41198 vdd.n10419 vdd.n10313 9.3
R41199 vdd.n10419 vdd.n10418 9.3
R41200 vdd.n10418 vdd.n10417 9.3
R41201 vdd.n10423 vdd.n10309 9.3
R41202 vdd.n10309 vdd.n10308 9.3
R41203 vdd.n10308 vdd.n10307 9.3
R41204 vdd.n10434 vdd.n10433 9.3
R41205 vdd.n10433 vdd.n10432 9.3
R41206 vdd.n10432 vdd.n10431 9.3
R41207 vdd.n10303 vdd.n10299 9.3
R41208 vdd.n10299 vdd.n10296 9.3
R41209 vdd.n10442 vdd.n10296 9.3
R41210 vdd.n10451 vdd.n10287 9.3
R41211 vdd.n10452 vdd.n10451 9.3
R41212 vdd.n10453 vdd.n10452 9.3
R41213 vdd.n10462 vdd.n10461 9.3
R41214 vdd.n10462 vdd.n10280 9.3
R41215 vdd.n10280 vdd.n10279 9.3
R41216 vdd.n10275 vdd.n10274 9.3
R41217 vdd.n10468 vdd.n10275 9.3
R41218 vdd.n10468 vdd.n10467 9.3
R41219 vdd.n10474 vdd.n10473 9.3
R41220 vdd.n10474 vdd.n10272 9.3
R41221 vdd.n12637 vdd.n12636 9.3
R41222 vdd.n12636 vdd.n12635 9.3
R41223 vdd.n12635 vdd.n12634 9.3
R41224 vdd.n12641 vdd.n10025 9.3
R41225 vdd.n12642 vdd.n12641 9.3
R41226 vdd.n12643 vdd.n12642 9.3
R41227 vdd.n12652 vdd.n12651 9.3
R41228 vdd.n12652 vdd.n10019 9.3
R41229 vdd.n10019 vdd.n10018 9.3
R41230 vdd.n12660 vdd.n10016 9.3
R41231 vdd.n12660 vdd.n12659 9.3
R41232 vdd.n12659 vdd.n12658 9.3
R41233 vdd.n10012 vdd.n9987 9.3
R41234 vdd.n10012 vdd.n9983 9.3
R41235 vdd.n9983 vdd.n9981 9.3
R41236 vdd.n10004 vdd.n10003 9.3
R41237 vdd.n10005 vdd.n10004 9.3
R41238 vdd.n10006 vdd.n10005 9.3
R41239 vdd.n9973 vdd.n9972 9.3
R41240 vdd.n12672 vdd.n9973 9.3
R41241 vdd.n12683 vdd.n12682 9.3
R41242 vdd.n12682 vdd.n12681 9.3
R41243 vdd.n12688 vdd.n12687 9.3
R41244 vdd.n12689 vdd.n12688 9.3
R41245 vdd.n12690 vdd.n12689 9.3
R41246 vdd.n9936 vdd.n9935 9.3
R41247 vdd.n9937 vdd.n9936 9.3
R41248 vdd.n9955 vdd.n9937 9.3
R41249 vdd.n9947 vdd.n9946 9.3
R41250 vdd.n9946 vdd.n9921 9.3
R41251 vdd.n9938 vdd.n9921 9.3
R41252 vdd.n12703 vdd.n12702 9.3
R41253 vdd.n12702 vdd.n9916 9.3
R41254 vdd.n9922 vdd.n9916 9.3
R41255 vdd.n12713 vdd.n9911 9.3
R41256 vdd.n12713 vdd.n12712 9.3
R41257 vdd.n12712 vdd.n12711 9.3
R41258 vdd.n12718 vdd.n12717 9.3
R41259 vdd.n12719 vdd.n12718 9.3
R41260 vdd.n12720 vdd.n12719 9.3
R41261 vdd.n9897 vdd.n9891 9.3
R41262 vdd.n9898 vdd.n9897 9.3
R41263 vdd.n9900 vdd.n9898 9.3
R41264 vdd.n12735 vdd.n12734 9.3
R41265 vdd.n12735 vdd.n9869 9.3
R41266 vdd.n9869 vdd.n9868 9.3
R41267 vdd.n12743 vdd.n9866 9.3
R41268 vdd.n12743 vdd.n12742 9.3
R41269 vdd.n12742 vdd.n12741 9.3
R41270 vdd.n9862 vdd.n9840 9.3
R41271 vdd.n9862 vdd.n9836 9.3
R41272 vdd.n9836 vdd.n9834 9.3
R41273 vdd.n9854 vdd.n9853 9.3
R41274 vdd.n9855 vdd.n9854 9.3
R41275 vdd.n9856 vdd.n9855 9.3
R41276 vdd.n12758 vdd.n12757 9.3
R41277 vdd.n12757 vdd.n12756 9.3
R41278 vdd.n12756 vdd.n12755 9.3
R41279 vdd.n12762 vdd.n9810 9.3
R41280 vdd.n12763 vdd.n12762 9.3
R41281 vdd.n12764 vdd.n12763 9.3
R41282 vdd.n12773 vdd.n12772 9.3
R41283 vdd.n12773 vdd.n9782 9.3
R41284 vdd.n9813 vdd.n9782 9.3
R41285 vdd.n12781 vdd.n12780 9.3
R41286 vdd.n12780 vdd.n12779 9.3
R41287 vdd.n9795 vdd.n9793 9.3
R41288 vdd.n9799 vdd.n9793 9.3
R41289 vdd.n9790 vdd.n9786 9.3
R41290 vdd.n9790 vdd.n9768 9.3
R41291 vdd.n9769 vdd.n9768 9.3
R41292 vdd.n12798 vdd.n12797 9.3
R41293 vdd.n12797 vdd.n9762 9.3
R41294 vdd.n9766 vdd.n9762 9.3
R41295 vdd.n12808 vdd.n9756 9.3
R41296 vdd.n12808 vdd.n12807 9.3
R41297 vdd.n12807 vdd.n12806 9.3
R41298 vdd.n12813 vdd.n12812 9.3
R41299 vdd.n12814 vdd.n12813 9.3
R41300 vdd.n12815 vdd.n12814 9.3
R41301 vdd.n9726 vdd.n9725 9.3
R41302 vdd.n9727 vdd.n9726 9.3
R41303 vdd.n9745 vdd.n9727 9.3
R41304 vdd.n9737 vdd.n9736 9.3
R41305 vdd.n9736 vdd.n9735 9.3
R41306 vdd.n9735 vdd.n9715 9.3
R41307 vdd.n12828 vdd.n12827 9.3
R41308 vdd.n12827 vdd.n9691 9.3
R41309 vdd.n9714 vdd.n9691 9.3
R41310 vdd.n9705 vdd.n9699 9.3
R41311 vdd.n9705 vdd.n9704 9.3
R41312 vdd.n9704 vdd.n9703 9.3
R41313 vdd.n12845 vdd.n12844 9.3
R41314 vdd.n12844 vdd.n12843 9.3
R41315 vdd.n12843 vdd.n12842 9.3
R41316 vdd.n12849 vdd.n9665 9.3
R41317 vdd.n12850 vdd.n12849 9.3
R41318 vdd.n12851 vdd.n12850 9.3
R41319 vdd.n12860 vdd.n12859 9.3
R41320 vdd.n12860 vdd.n9659 9.3
R41321 vdd.n9659 vdd.n9658 9.3
R41322 vdd.n12868 vdd.n9656 9.3
R41323 vdd.n12868 vdd.n12867 9.3
R41324 vdd.n12867 vdd.n12866 9.3
R41325 vdd.n9652 vdd.n9627 9.3
R41326 vdd.n9652 vdd.n9623 9.3
R41327 vdd.n9623 vdd.n9621 9.3
R41328 vdd.n9644 vdd.n9643 9.3
R41329 vdd.n9645 vdd.n9644 9.3
R41330 vdd.n9646 vdd.n9645 9.3
R41331 vdd.n9613 vdd.n9612 9.3
R41332 vdd.n12880 vdd.n9613 9.3
R41333 vdd.n12891 vdd.n12890 9.3
R41334 vdd.n12890 vdd.n12889 9.3
R41335 vdd.n12896 vdd.n12895 9.3
R41336 vdd.n12897 vdd.n12896 9.3
R41337 vdd.n12898 vdd.n12897 9.3
R41338 vdd.n9577 vdd.n9576 9.3
R41339 vdd.n9578 vdd.n9577 9.3
R41340 vdd.n9595 vdd.n9578 9.3
R41341 vdd.n9587 vdd.n9586 9.3
R41342 vdd.n9586 vdd.n9563 9.3
R41343 vdd.n9564 vdd.n9563 9.3
R41344 vdd.n12911 vdd.n12910 9.3
R41345 vdd.n12910 vdd.n9557 9.3
R41346 vdd.n9561 vdd.n9557 9.3
R41347 vdd.n12921 vdd.n9551 9.3
R41348 vdd.n12921 vdd.n12920 9.3
R41349 vdd.n12920 vdd.n12919 9.3
R41350 vdd.n12926 vdd.n12925 9.3
R41351 vdd.n12927 vdd.n12926 9.3
R41352 vdd.n12928 vdd.n12927 9.3
R41353 vdd.n9536 vdd.n9530 9.3
R41354 vdd.n9537 vdd.n9536 9.3
R41355 vdd.n9539 vdd.n9537 9.3
R41356 vdd.n12943 vdd.n12942 9.3
R41357 vdd.n12943 vdd.n9509 9.3
R41358 vdd.n9509 vdd.n9508 9.3
R41359 vdd.n12951 vdd.n9506 9.3
R41360 vdd.n12951 vdd.n12950 9.3
R41361 vdd.n12950 vdd.n12949 9.3
R41362 vdd.n9502 vdd.n9480 9.3
R41363 vdd.n9502 vdd.n9476 9.3
R41364 vdd.n9476 vdd.n9474 9.3
R41365 vdd.n9494 vdd.n9493 9.3
R41366 vdd.n9495 vdd.n9494 9.3
R41367 vdd.n9496 vdd.n9495 9.3
R41368 vdd.n12966 vdd.n12965 9.3
R41369 vdd.n12965 vdd.n12964 9.3
R41370 vdd.n12964 vdd.n12963 9.3
R41371 vdd.n12970 vdd.n9451 9.3
R41372 vdd.n12971 vdd.n12970 9.3
R41373 vdd.n12972 vdd.n12971 9.3
R41374 vdd.n12981 vdd.n12980 9.3
R41375 vdd.n12981 vdd.n9422 9.3
R41376 vdd.n9422 vdd.n9421 9.3
R41377 vdd.n12989 vdd.n12988 9.3
R41378 vdd.n12988 vdd.n12987 9.3
R41379 vdd.n9436 vdd.n9433 9.3
R41380 vdd.n9440 vdd.n9433 9.3
R41381 vdd.n9430 vdd.n9426 9.3
R41382 vdd.n9430 vdd.n9408 9.3
R41383 vdd.n9434 vdd.n9408 9.3
R41384 vdd.n13006 vdd.n13005 9.3
R41385 vdd.n13005 vdd.n9402 9.3
R41386 vdd.n9406 vdd.n9402 9.3
R41387 vdd.n13016 vdd.n9396 9.3
R41388 vdd.n13016 vdd.n13015 9.3
R41389 vdd.n13015 vdd.n13014 9.3
R41390 vdd.n13021 vdd.n13020 9.3
R41391 vdd.n13022 vdd.n13021 9.3
R41392 vdd.n13023 vdd.n13022 9.3
R41393 vdd.n9366 vdd.n9365 9.3
R41394 vdd.n9367 vdd.n9366 9.3
R41395 vdd.n9385 vdd.n9367 9.3
R41396 vdd.n9377 vdd.n9376 9.3
R41397 vdd.n9376 vdd.n9375 9.3
R41398 vdd.n9375 vdd.n9355 9.3
R41399 vdd.n13036 vdd.n13035 9.3
R41400 vdd.n13035 vdd.n9331 9.3
R41401 vdd.n9354 vdd.n9331 9.3
R41402 vdd.n9345 vdd.n9339 9.3
R41403 vdd.n9345 vdd.n9344 9.3
R41404 vdd.n9344 vdd.n9343 9.3
R41405 vdd.n13053 vdd.n13052 9.3
R41406 vdd.n13052 vdd.n13051 9.3
R41407 vdd.n13051 vdd.n13050 9.3
R41408 vdd.n13057 vdd.n9305 9.3
R41409 vdd.n13058 vdd.n13057 9.3
R41410 vdd.n13059 vdd.n13058 9.3
R41411 vdd.n13068 vdd.n13067 9.3
R41412 vdd.n13068 vdd.n9299 9.3
R41413 vdd.n9299 vdd.n9298 9.3
R41414 vdd.n13076 vdd.n9295 9.3
R41415 vdd.n13076 vdd.n13075 9.3
R41416 vdd.n13075 vdd.n13074 9.3
R41417 vdd.n10365 vdd.n10364 9.3
R41418 vdd.n10365 vdd.n9291 9.3
R41419 vdd.n9291 vdd.n9289 9.3
R41420 vdd.n10373 vdd.n10372 9.3
R41421 vdd.n10372 vdd.n10371 9.3
R41422 vdd.n10371 vdd.n10370 9.3
R41423 vdd.n10378 vdd.n10377 9.3
R41424 vdd.n10379 vdd.n10378 9.3
R41425 vdd.n10341 vdd.n10337 9.3
R41426 vdd.n10388 vdd.n10337 9.3
R41427 vdd.n10140 vdd.n10057 9.3
R41428 vdd.n10190 vdd.n10138 9.3
R41429 vdd.n12606 vdd.n12605 9.3
R41430 vdd.n10108 vdd.n10107 9.3
R41431 vdd.n10102 vdd.n10099 9.3
R41432 vdd.n10229 vdd.n10103 9.3
R41433 vdd.n10242 vdd.n10238 9.3
R41434 vdd.n10484 vdd.n10483 9.3
R41435 vdd.n10489 vdd.n10480 9.3
R41436 vdd.n12569 vdd.n12568 9.3
R41437 vdd.n12568 vdd.n12567 9.3
R41438 vdd.n10056 vdd.n10049 9.3
R41439 vdd.n10160 vdd.n10159 9.3
R41440 vdd.n10159 vdd.n10158 9.3
R41441 vdd.n10158 vdd.n10157 9.3
R41442 vdd.n11602 vdd.n11601 9.3
R41443 vdd.n11601 vdd.n11564 9.3
R41444 vdd.n11587 vdd.n11558 9.3
R41445 vdd.n11559 vdd.n11558 9.3
R41446 vdd.n11560 vdd.n11559 9.3
R41447 vdd.n11942 vdd.n11941 9.3
R41448 vdd.n11943 vdd.n11942 9.3
R41449 vdd.n11944 vdd.n11943 9.3
R41450 vdd.n11449 vdd.n11447 9.3
R41451 vdd.n11447 vdd.n11445 9.3
R41452 vdd.n11533 vdd.n11454 9.3
R41453 vdd.n11525 vdd.n11454 9.3
R41454 vdd.n11527 vdd.n11525 9.3
R41455 vdd.n11522 vdd.n11521 9.3
R41456 vdd.n11523 vdd.n11522 9.3
R41457 vdd.n11523 vdd.n11437 9.3
R41458 vdd.n11967 vdd.n11966 9.3
R41459 vdd.n11966 vdd.n11965 9.3
R41460 vdd.n11430 vdd.n11429 9.3
R41461 vdd.n11972 vdd.n11430 9.3
R41462 vdd.n11479 vdd.n11478 9.3
R41463 vdd.n11480 vdd.n11479 9.3
R41464 vdd.n11481 vdd.n11480 9.3
R41465 vdd.n11989 vdd.n11411 9.3
R41466 vdd.n11989 vdd.n11988 9.3
R41467 vdd.n11988 vdd.n11987 9.3
R41468 vdd.n11993 vdd.n11407 9.3
R41469 vdd.n11407 vdd.n11406 9.3
R41470 vdd.n11406 vdd.n11405 9.3
R41471 vdd.n12004 vdd.n12003 9.3
R41472 vdd.n12003 vdd.n12002 9.3
R41473 vdd.n12002 vdd.n12001 9.3
R41474 vdd.n11401 vdd.n11379 9.3
R41475 vdd.n11379 vdd.n11377 9.3
R41476 vdd.n11377 vdd.n11375 9.3
R41477 vdd.n11391 vdd.n11390 9.3
R41478 vdd.n11392 vdd.n11391 9.3
R41479 vdd.n11393 vdd.n11392 9.3
R41480 vdd.n12020 vdd.n11364 9.3
R41481 vdd.n12020 vdd.n12019 9.3
R41482 vdd.n12019 vdd.n12018 9.3
R41483 vdd.n12024 vdd.n11338 9.3
R41484 vdd.n11338 vdd.n11336 9.3
R41485 vdd.n11336 vdd.n11334 9.3
R41486 vdd.n11357 vdd.n11339 9.3
R41487 vdd.n11357 vdd.n11335 9.3
R41488 vdd.n11335 vdd.n11333 9.3
R41489 vdd.n11350 vdd.n11349 9.3
R41490 vdd.n11351 vdd.n11350 9.3
R41491 vdd.n11351 vdd.n11326 9.3
R41492 vdd.n12040 vdd.n12039 9.3
R41493 vdd.n12039 vdd.n12038 9.3
R41494 vdd.n12038 vdd.n12037 9.3
R41495 vdd.n12044 vdd.n11313 9.3
R41496 vdd.n12045 vdd.n12044 9.3
R41497 vdd.n12046 vdd.n12045 9.3
R41498 vdd.n12055 vdd.n12054 9.3
R41499 vdd.n12055 vdd.n11284 9.3
R41500 vdd.n11284 vdd.n11282 9.3
R41501 vdd.n11309 vdd.n11289 9.3
R41502 vdd.n11309 vdd.n11308 9.3
R41503 vdd.n11308 vdd.n11307 9.3
R41504 vdd.n11299 vdd.n11298 9.3
R41505 vdd.n11298 vdd.n11291 9.3
R41506 vdd.n11291 vdd.n11274 9.3
R41507 vdd.n12068 vdd.n11267 9.3
R41508 vdd.n12068 vdd.n12067 9.3
R41509 vdd.n12067 vdd.n12066 9.3
R41510 vdd.n12077 vdd.n12076 9.3
R41511 vdd.n11266 vdd.n11244 9.3
R41512 vdd.n11244 vdd.n11242 9.3
R41513 vdd.n11242 vdd.n11240 9.3
R41514 vdd.n11256 vdd.n11255 9.3
R41515 vdd.n11257 vdd.n11256 9.3
R41516 vdd.n11258 vdd.n11257 9.3
R41517 vdd.n12093 vdd.n11227 9.3
R41518 vdd.n12093 vdd.n12092 9.3
R41519 vdd.n12092 vdd.n12091 9.3
R41520 vdd.n12097 vdd.n11223 9.3
R41521 vdd.n11223 vdd.n11222 9.3
R41522 vdd.n11222 vdd.n11221 9.3
R41523 vdd.n12108 vdd.n12107 9.3
R41524 vdd.n12107 vdd.n12106 9.3
R41525 vdd.n12106 vdd.n12105 9.3
R41526 vdd.n11217 vdd.n11195 9.3
R41527 vdd.n11195 vdd.n11193 9.3
R41528 vdd.n11193 vdd.n11191 9.3
R41529 vdd.n11207 vdd.n11206 9.3
R41530 vdd.n11208 vdd.n11207 9.3
R41531 vdd.n11209 vdd.n11208 9.3
R41532 vdd.n12124 vdd.n11180 9.3
R41533 vdd.n12124 vdd.n12123 9.3
R41534 vdd.n12123 vdd.n12122 9.3
R41535 vdd.n12130 vdd.n11175 9.3
R41536 vdd.n12131 vdd.n12130 9.3
R41537 vdd.n12132 vdd.n12131 9.3
R41538 vdd.n12141 vdd.n12140 9.3
R41539 vdd.n12141 vdd.n11148 9.3
R41540 vdd.n11148 vdd.n11146 9.3
R41541 vdd.n11171 vdd.n11153 9.3
R41542 vdd.n11171 vdd.n11170 9.3
R41543 vdd.n11170 vdd.t298 9.3
R41544 vdd.n11162 vdd.n11161 9.3
R41545 vdd.n11161 vdd.n11155 9.3
R41546 vdd.n11155 vdd.n11138 9.3
R41547 vdd.n12155 vdd.n12154 9.3
R41548 vdd.n12154 vdd.n12153 9.3
R41549 vdd.n12153 vdd.n12152 9.3
R41550 vdd.n12159 vdd.n11125 9.3
R41551 vdd.n12160 vdd.n12159 9.3
R41552 vdd.n12161 vdd.n12160 9.3
R41553 vdd.n12170 vdd.n12169 9.3
R41554 vdd.n12170 vdd.n11108 9.3
R41555 vdd.n11108 vdd.n11106 9.3
R41556 vdd.n11121 vdd.n11113 9.3
R41557 vdd.n11121 vdd.n11120 9.3
R41558 vdd.n11120 vdd.n11119 9.3
R41559 vdd.n12181 vdd.n11091 9.3
R41560 vdd.n12185 vdd.n11088 9.3
R41561 vdd.n11088 vdd.n11087 9.3
R41562 vdd.n11087 vdd.n11086 9.3
R41563 vdd.n12196 vdd.n12195 9.3
R41564 vdd.n12195 vdd.n12194 9.3
R41565 vdd.n12194 vdd.n12193 9.3
R41566 vdd.n11082 vdd.n11060 9.3
R41567 vdd.n11060 vdd.n11058 9.3
R41568 vdd.n11058 vdd.n11056 9.3
R41569 vdd.n11072 vdd.n11071 9.3
R41570 vdd.n11073 vdd.n11072 9.3
R41571 vdd.n11074 vdd.n11073 9.3
R41572 vdd.n12212 vdd.n11042 9.3
R41573 vdd.n12212 vdd.n12211 9.3
R41574 vdd.n12211 vdd.n12210 9.3
R41575 vdd.n12216 vdd.n11038 9.3
R41576 vdd.n11038 vdd.n11037 9.3
R41577 vdd.n11047 vdd.n11037 9.3
R41578 vdd.n12227 vdd.n12226 9.3
R41579 vdd.n12226 vdd.n12225 9.3
R41580 vdd.n12225 vdd.n12224 9.3
R41581 vdd.n11033 vdd.n11015 9.3
R41582 vdd.n11015 vdd.n11013 9.3
R41583 vdd.n11013 vdd.n11011 9.3
R41584 vdd.n11026 vdd.n11025 9.3
R41585 vdd.n11027 vdd.n11026 9.3
R41586 vdd.n11027 vdd.n11004 9.3
R41587 vdd.n12245 vdd.n12244 9.3
R41588 vdd.n12244 vdd.n12243 9.3
R41589 vdd.n12243 vdd.n12242 9.3
R41590 vdd.n12249 vdd.n10991 9.3
R41591 vdd.n12250 vdd.n12249 9.3
R41592 vdd.n12251 vdd.n12250 9.3
R41593 vdd.n12260 vdd.n12259 9.3
R41594 vdd.n12260 vdd.n10962 9.3
R41595 vdd.n10962 vdd.n10960 9.3
R41596 vdd.n10987 vdd.n10967 9.3
R41597 vdd.n10987 vdd.n10986 9.3
R41598 vdd.n10986 vdd.n10985 9.3
R41599 vdd.n10977 vdd.n10976 9.3
R41600 vdd.n10976 vdd.n10969 9.3
R41601 vdd.n10969 vdd.n10952 9.3
R41602 vdd.n12273 vdd.n10950 9.3
R41603 vdd.n12273 vdd.n12272 9.3
R41604 vdd.n12272 vdd.n12271 9.3
R41605 vdd.n10946 vdd.n10920 9.3
R41606 vdd.n10921 vdd.n10920 9.3
R41607 vdd.n12278 vdd.n10921 9.3
R41608 vdd.n10945 vdd.n10919 9.3
R41609 vdd.n10935 vdd.n10934 9.3
R41610 vdd.n10936 vdd.n10935 9.3
R41611 vdd.n10937 vdd.n10936 9.3
R41612 vdd.n12295 vdd.n10902 9.3
R41613 vdd.n12295 vdd.n12294 9.3
R41614 vdd.n12294 vdd.n12293 9.3
R41615 vdd.n12299 vdd.n10898 9.3
R41616 vdd.n10898 vdd.n10897 9.3
R41617 vdd.n10897 vdd.n10896 9.3
R41618 vdd.n12310 vdd.n12309 9.3
R41619 vdd.n12309 vdd.n12308 9.3
R41620 vdd.n12308 vdd.n12307 9.3
R41621 vdd.n10892 vdd.n10870 9.3
R41622 vdd.n10870 vdd.n10868 9.3
R41623 vdd.n10868 vdd.n10866 9.3
R41624 vdd.n10882 vdd.n10881 9.3
R41625 vdd.n10883 vdd.n10882 9.3
R41626 vdd.n10884 vdd.n10883 9.3
R41627 vdd.n12326 vdd.n10855 9.3
R41628 vdd.n12326 vdd.n12325 9.3
R41629 vdd.n12325 vdd.n12324 9.3
R41630 vdd.n12330 vdd.n10829 9.3
R41631 vdd.n10829 vdd.n10827 9.3
R41632 vdd.n10827 vdd.n10825 9.3
R41633 vdd.n10848 vdd.n10830 9.3
R41634 vdd.n10848 vdd.n10826 9.3
R41635 vdd.n10826 vdd.n10824 9.3
R41636 vdd.n10841 vdd.n10840 9.3
R41637 vdd.n10842 vdd.n10841 9.3
R41638 vdd.n10842 vdd.n10817 9.3
R41639 vdd.n12346 vdd.n12345 9.3
R41640 vdd.n12345 vdd.n12344 9.3
R41641 vdd.n12344 vdd.n12343 9.3
R41642 vdd.n12350 vdd.n10804 9.3
R41643 vdd.n12351 vdd.n12350 9.3
R41644 vdd.n12352 vdd.n12351 9.3
R41645 vdd.n12361 vdd.n12360 9.3
R41646 vdd.n12361 vdd.n10776 9.3
R41647 vdd.n10776 vdd.n10774 9.3
R41648 vdd.n10800 vdd.n10781 9.3
R41649 vdd.n10800 vdd.n10799 9.3
R41650 vdd.n10799 vdd.n10798 9.3
R41651 vdd.n10790 vdd.n10789 9.3
R41652 vdd.n10789 vdd.n10783 9.3
R41653 vdd.n10783 vdd.n10764 9.3
R41654 vdd.n12375 vdd.n12374 9.3
R41655 vdd.n12374 vdd.n12373 9.3
R41656 vdd.n12373 vdd.n12372 9.3
R41657 vdd.n12376 vdd.n10751 9.3
R41658 vdd.n12387 vdd.n12386 9.3
R41659 vdd.n12386 vdd.n12385 9.3
R41660 vdd.n12385 vdd.n12384 9.3
R41661 vdd.n10745 vdd.n10723 9.3
R41662 vdd.n10723 vdd.n10721 9.3
R41663 vdd.n10721 vdd.n10719 9.3
R41664 vdd.n10735 vdd.n10734 9.3
R41665 vdd.n10736 vdd.n10735 9.3
R41666 vdd.n10737 vdd.n10736 9.3
R41667 vdd.n12403 vdd.n10705 9.3
R41668 vdd.n12403 vdd.n12402 9.3
R41669 vdd.n12402 vdd.n12401 9.3
R41670 vdd.n12407 vdd.n10701 9.3
R41671 vdd.n10701 vdd.n10700 9.3
R41672 vdd.n10710 vdd.n10700 9.3
R41673 vdd.n12418 vdd.n12417 9.3
R41674 vdd.n12417 vdd.n12416 9.3
R41675 vdd.n12416 vdd.n12415 9.3
R41676 vdd.n10696 vdd.n10675 9.3
R41677 vdd.n10675 vdd.n10673 9.3
R41678 vdd.n10673 vdd.n10671 9.3
R41679 vdd.n10686 vdd.n10685 9.3
R41680 vdd.n10687 vdd.n10686 9.3
R41681 vdd.n10688 vdd.n10687 9.3
R41682 vdd.n12435 vdd.n12434 9.3
R41683 vdd.n12434 vdd.n12433 9.3
R41684 vdd.n12433 vdd.n12432 9.3
R41685 vdd.n12439 vdd.n10653 9.3
R41686 vdd.n12440 vdd.n12439 9.3
R41687 vdd.n12441 vdd.n12440 9.3
R41688 vdd.n12450 vdd.n12449 9.3
R41689 vdd.n12450 vdd.n10625 9.3
R41690 vdd.n10625 vdd.n10623 9.3
R41691 vdd.n10649 vdd.n10630 9.3
R41692 vdd.n10649 vdd.n10648 9.3
R41693 vdd.n10648 vdd.n10647 9.3
R41694 vdd.n10639 vdd.n10638 9.3
R41695 vdd.n10638 vdd.n10632 9.3
R41696 vdd.n10632 vdd.n10615 9.3
R41697 vdd.n12464 vdd.n12463 9.3
R41698 vdd.n12463 vdd.n12462 9.3
R41699 vdd.n12462 vdd.n12461 9.3
R41700 vdd.n12468 vdd.n10602 9.3
R41701 vdd.n12469 vdd.n12468 9.3
R41702 vdd.n12470 vdd.n12469 9.3
R41703 vdd.n12479 vdd.n12478 9.3
R41704 vdd.n12479 vdd.n10586 9.3
R41705 vdd.n10586 vdd.n10584 9.3
R41706 vdd.n10601 vdd.n10600 9.3
R41707 vdd.n12491 vdd.n10570 9.3
R41708 vdd.n12491 vdd.n12490 9.3
R41709 vdd.n12490 vdd.n12489 9.3
R41710 vdd.n12495 vdd.n10566 9.3
R41711 vdd.n10566 vdd.n10565 9.3
R41712 vdd.n10565 vdd.n10564 9.3
R41713 vdd.n12506 vdd.n12505 9.3
R41714 vdd.n12505 vdd.n12504 9.3
R41715 vdd.n12504 vdd.n12503 9.3
R41716 vdd.n10560 vdd.n10532 9.3
R41717 vdd.n10532 vdd.n10530 9.3
R41718 vdd.n10530 vdd.n10528 9.3
R41719 vdd.n10550 vdd.n10549 9.3
R41720 vdd.n10551 vdd.n10550 9.3
R41721 vdd.n10552 vdd.n10551 9.3
R41722 vdd.n10543 vdd.n10539 9.3
R41723 vdd.n10543 vdd.n10522 9.3
R41724 vdd.n12520 vdd.n10522 9.3
R41725 vdd.n12526 vdd.n12525 9.3
R41726 vdd.n12527 vdd.n12526 9.3
R41727 vdd.n11781 vdd.n11779 9.3
R41728 vdd.n11672 vdd.n11670 9.3
R41729 vdd.n11736 vdd.n11735 9.3
R41730 vdd.n11734 vdd.n11731 9.3
R41731 vdd.n11737 vdd.n11725 9.3
R41732 vdd.n11738 vdd.n11737 9.3
R41733 vdd.n11743 vdd.n11742 9.3
R41734 vdd.n11704 vdd.n11703 9.3
R41735 vdd.n11709 vdd.n11700 9.3
R41736 vdd.n11698 vdd.n11697 9.3
R41737 vdd.n11690 vdd.n11684 9.3
R41738 vdd.n11696 vdd.n11687 9.3
R41739 vdd.n11699 vdd.n11694 9.3
R41740 vdd.n11711 vdd.n11710 9.3
R41741 vdd.n11708 vdd.n11707 9.3
R41742 vdd.n11706 vdd.n11705 9.3
R41743 vdd.n11702 vdd.n11691 9.3
R41744 vdd.n11718 vdd.n11717 9.3
R41745 vdd.n11828 vdd.n11815 9.3
R41746 vdd.n11822 vdd.n11815 9.3
R41747 vdd.n11831 vdd.n11814 9.3
R41748 vdd.n11830 vdd.n11829 9.3
R41749 vdd.n11827 vdd.n11817 9.3
R41750 vdd.n11827 vdd.n11826 9.3
R41751 vdd.n11820 vdd.n11816 9.3
R41752 vdd.n11847 vdd.n11842 9.3
R41753 vdd.n11852 vdd.n11851 9.3
R41754 vdd.n11860 vdd.n11810 9.3
R41755 vdd.n11863 vdd.n11862 9.3
R41756 vdd.n11866 vdd.n11865 9.3
R41757 vdd.n11853 vdd.n11839 9.3
R41758 vdd.n11850 vdd.n11841 9.3
R41759 vdd.n11849 vdd.n11848 9.3
R41760 vdd.n11846 vdd.n11845 9.3
R41761 vdd.n11857 vdd.n11838 9.3
R41762 vdd.n11859 vdd.n11858 9.3
R41763 vdd.n11913 vdd.n11912 9.3
R41764 vdd.n11920 vdd.n11919 9.3
R41765 vdd.n11920 vdd.n9287 9.3
R41766 vdd.n11659 vdd.n9287 9.3
R41767 vdd.n13085 vdd.n13084 9.3
R41768 vdd.n13123 vdd.n13122 9.3
R41769 vdd.n13125 vdd.n9269 9.3
R41770 vdd.n13193 vdd.n9217 9.3
R41771 vdd.n13183 vdd.n13182 9.3
R41772 vdd.n13208 vdd.n9205 9.3
R41773 vdd.n13249 vdd.n9176 9.3
R41774 vdd.n13272 vdd.n9161 9.3
R41775 vdd.n13292 vdd.n13291 9.3
R41776 vdd.n13293 vdd.n9145 9.3
R41777 vdd.n9145 vdd.n9143 9.3
R41778 vdd.n9143 vdd.n9140 9.3
R41779 vdd.n13290 vdd.n9147 9.3
R41780 vdd.n9163 vdd.n9162 9.3
R41781 vdd.n9164 vdd.n9163 9.3
R41782 vdd.n9179 vdd.n9164 9.3
R41783 vdd.n13251 vdd.n13250 9.3
R41784 vdd.n13181 vdd.n13180 9.3
R41785 vdd.n9268 vdd.n9218 9.3
R41786 vdd.n13121 vdd.n9270 9.3
R41787 vdd.n13121 vdd.n9265 9.3
R41788 vdd.n13117 vdd.n9265 9.3
R41789 vdd.n13124 vdd.n9267 9.3
R41790 vdd.n13128 vdd.n13126 9.3
R41791 vdd.n13128 vdd.n13127 9.3
R41792 vdd.n13127 vdd.n9239 9.3
R41793 vdd.n13195 vdd.n13194 9.3
R41794 vdd.n13195 vdd.n9215 9.3
R41795 vdd.n9215 vdd.n9213 9.3
R41796 vdd.n13192 vdd.n13191 9.3
R41797 vdd.n13184 vdd.n9219 9.3
R41798 vdd.n13185 vdd.n13184 9.3
R41799 vdd.n13186 vdd.n13185 9.3
R41800 vdd.n13207 vdd.n9207 9.3
R41801 vdd.n13207 vdd.n13206 9.3
R41802 vdd.n13206 vdd.n13205 9.3
R41803 vdd.n13210 vdd.n13209 9.3
R41804 vdd.n13213 vdd.n13212 9.3
R41805 vdd.n13213 vdd.n9171 9.3
R41806 vdd.n13217 vdd.n9171 9.3
R41807 vdd.n13253 vdd.n13252 9.3
R41808 vdd.n13253 vdd.n9172 9.3
R41809 vdd.n9185 vdd.n9172 9.3
R41810 vdd.n13271 vdd.n13270 9.3
R41811 vdd.n13274 vdd.n13273 9.3
R41812 vdd.n13275 vdd.n13274 9.3
R41813 vdd.n13276 vdd.n13275 9.3
R41814 vdd.n13297 vdd.n9146 9.3
R41815 vdd.n13341 vdd.n13340 9.3
R41816 vdd.n13415 vdd.n13414 9.3
R41817 vdd.n13418 vdd.n9038 9.3
R41818 vdd.n13487 vdd.n8997 9.3
R41819 vdd.n13477 vdd.n13476 9.3
R41820 vdd.n13564 vdd.n8939 9.3
R41821 vdd.n13584 vdd.n13583 9.3
R41822 vdd.n13589 vdd.n8925 9.3
R41823 vdd.n13633 vdd.n13632 9.3
R41824 vdd.n13709 vdd.n13708 9.3
R41825 vdd.n13711 vdd.n8817 9.3
R41826 vdd.n13767 vdd.n8780 9.3
R41827 vdd.n13757 vdd.n13756 9.3
R41828 vdd.n13846 vdd.n8723 9.3
R41829 vdd.n13850 vdd.n13847 9.3
R41830 vdd.n13893 vdd.n8686 9.3
R41831 vdd.n8674 vdd.n8673 9.3
R41832 vdd.n13985 vdd.n8606 9.3
R41833 vdd.n14057 vdd.n8569 9.3
R41834 vdd.n14047 vdd.n14046 9.3
R41835 vdd.n8557 vdd.n8556 9.3
R41836 vdd.n14135 vdd.n8502 9.3
R41837 vdd.n14139 vdd.n14136 9.3
R41838 vdd.n14182 vdd.n8462 9.3
R41839 vdd.n8450 vdd.n8449 9.3
R41840 vdd.n14275 vdd.n8384 9.3
R41841 vdd.n14332 vdd.n8351 9.3
R41842 vdd.n14331 vdd.n14330 9.3
R41843 vdd.n14274 vdd.n8382 9.3
R41844 vdd.n8402 vdd.n8400 9.3
R41845 vdd.n8400 vdd.n8397 9.3
R41846 vdd.n8446 vdd.n8445 9.3
R41847 vdd.n14199 vdd.n14198 9.3
R41848 vdd.n14198 vdd.n14197 9.3
R41849 vdd.n14197 vdd.n8426 9.3
R41850 vdd.n8466 vdd.n8465 9.3
R41851 vdd.n8463 vdd.n8461 9.3
R41852 vdd.n8461 vdd.n8459 9.3
R41853 vdd.n8485 vdd.n8459 9.3
R41854 vdd.n14141 vdd.n14140 9.3
R41855 vdd.n8505 vdd.n8504 9.3
R41856 vdd.n14129 vdd.n8505 9.3
R41857 vdd.n14129 vdd.n8489 9.3
R41858 vdd.n14074 vdd.n14073 9.3
R41859 vdd.n14056 vdd.n14055 9.3
R41860 vdd.n13984 vdd.n8604 9.3
R41861 vdd.n8624 vdd.n8622 9.3
R41862 vdd.n8622 vdd.n8619 9.3
R41863 vdd.n8669 vdd.n8668 9.3
R41864 vdd.n13909 vdd.n13908 9.3
R41865 vdd.n13908 vdd.n13907 9.3
R41866 vdd.n13907 vdd.n8646 9.3
R41867 vdd.n8689 vdd.n8688 9.3
R41868 vdd.n8687 vdd.n8685 9.3
R41869 vdd.n8685 vdd.n8683 9.3
R41870 vdd.n8708 vdd.n8683 9.3
R41871 vdd.n13852 vdd.n13851 9.3
R41872 vdd.n8726 vdd.n8725 9.3
R41873 vdd.n8727 vdd.n8726 9.3
R41874 vdd.n8727 vdd.n8712 9.3
R41875 vdd.n13755 vdd.n8770 9.3
R41876 vdd.n8816 vdd.n8781 9.3
R41877 vdd.n13688 vdd.n13687 9.3
R41878 vdd.n13648 vdd.n8849 9.3
R41879 vdd.n8869 vdd.n8849 9.3
R41880 vdd.n13662 vdd.n13661 9.3
R41881 vdd.n13634 vdd.n8877 9.3
R41882 vdd.n8877 vdd.n8875 9.3
R41883 vdd.n8883 vdd.n8875 9.3
R41884 vdd.n13631 vdd.n8879 9.3
R41885 vdd.n13585 vdd.n8924 9.3
R41886 vdd.n8924 vdd.n8922 9.3
R41887 vdd.n8922 vdd.n8918 9.3
R41888 vdd.n13582 vdd.n8926 9.3
R41889 vdd.n8942 vdd.n8941 9.3
R41890 vdd.n8943 vdd.n8942 9.3
R41891 vdd.n8958 vdd.n8943 9.3
R41892 vdd.n13475 vdd.n8985 9.3
R41893 vdd.n9037 vdd.n8998 9.3
R41894 vdd.n13396 vdd.n13395 9.3
R41895 vdd.n13356 vdd.n9069 9.3
R41896 vdd.n9089 vdd.n9069 9.3
R41897 vdd.n13370 vdd.n13369 9.3
R41898 vdd.n13342 vdd.n9097 9.3
R41899 vdd.n9097 vdd.n9095 9.3
R41900 vdd.n9104 vdd.n9095 9.3
R41901 vdd.n13339 vdd.n9100 9.3
R41902 vdd.n13299 vdd.n13298 9.3
R41903 vdd.n13296 vdd.n13295 9.3
R41904 vdd.n13295 vdd.n13294 9.3
R41905 vdd.n13294 vdd.n9132 9.3
R41906 vdd.n13344 vdd.n13343 9.3
R41907 vdd.n9124 vdd.n9123 9.3
R41908 vdd.n9125 vdd.n9124 9.3
R41909 vdd.n13401 vdd.n9048 9.3
R41910 vdd.n9048 vdd.n9046 9.3
R41911 vdd.n13399 vdd.n13398 9.3
R41912 vdd.n13393 vdd.n13392 9.3
R41913 vdd.n13392 vdd.n13391 9.3
R41914 vdd.n13413 vdd.n9039 9.3
R41915 vdd.n13413 vdd.n9034 9.3
R41916 vdd.n9034 vdd.n9032 9.3
R41917 vdd.n13416 vdd.n9036 9.3
R41918 vdd.n13422 vdd.n13419 9.3
R41919 vdd.n13422 vdd.n13421 9.3
R41920 vdd.n13421 vdd.n13420 9.3
R41921 vdd.n13489 vdd.n13488 9.3
R41922 vdd.n13489 vdd.n8995 9.3
R41923 vdd.n8995 vdd.n8993 9.3
R41924 vdd.n13486 vdd.n13485 9.3
R41925 vdd.n13478 vdd.n8999 9.3
R41926 vdd.n13479 vdd.n13478 9.3
R41927 vdd.n13480 vdd.n13479 9.3
R41928 vdd.n13502 vdd.n13501 9.3
R41929 vdd.n13501 vdd.n13500 9.3
R41930 vdd.n13500 vdd.n13499 9.3
R41931 vdd.n13506 vdd.n13505 9.3
R41932 vdd.n13506 vdd.n8951 9.3
R41933 vdd.n13510 vdd.n8951 9.3
R41934 vdd.n13544 vdd.n13543 9.3
R41935 vdd.n13544 vdd.n8952 9.3
R41936 vdd.n8964 vdd.n8952 9.3
R41937 vdd.n13563 vdd.n13562 9.3
R41938 vdd.n13566 vdd.n13565 9.3
R41939 vdd.n13567 vdd.n13566 9.3
R41940 vdd.n13568 vdd.n13567 9.3
R41941 vdd.n13591 vdd.n13590 9.3
R41942 vdd.n13588 vdd.n13587 9.3
R41943 vdd.n13587 vdd.n13586 9.3
R41944 vdd.n13586 vdd.n8910 9.3
R41945 vdd.n13636 vdd.n13635 9.3
R41946 vdd.n8903 vdd.n8902 9.3
R41947 vdd.n8904 vdd.n8903 9.3
R41948 vdd.n13694 vdd.n8827 9.3
R41949 vdd.n8827 vdd.n8825 9.3
R41950 vdd.n13692 vdd.n13691 9.3
R41951 vdd.n13685 vdd.n13684 9.3
R41952 vdd.n13684 vdd.n13683 9.3
R41953 vdd.n13707 vdd.n8818 9.3
R41954 vdd.n13707 vdd.n8813 9.3
R41955 vdd.n13703 vdd.n8813 9.3
R41956 vdd.n13710 vdd.n8815 9.3
R41957 vdd.n13714 vdd.n13712 9.3
R41958 vdd.n13714 vdd.n13713 9.3
R41959 vdd.n13713 vdd.n8796 9.3
R41960 vdd.n13769 vdd.n13768 9.3
R41961 vdd.n13769 vdd.n8778 9.3
R41962 vdd.n13745 vdd.n8778 9.3
R41963 vdd.n13766 vdd.n13765 9.3
R41964 vdd.n13758 vdd.n8782 9.3
R41965 vdd.n13759 vdd.n13758 9.3
R41966 vdd.n13760 vdd.n13759 9.3
R41967 vdd.n13782 vdd.n13781 9.3
R41968 vdd.n13781 vdd.n8767 9.3
R41969 vdd.n8767 vdd.n8765 9.3
R41970 vdd.n13787 vdd.n13786 9.3
R41971 vdd.n13787 vdd.n8732 9.3
R41972 vdd.n8749 vdd.n8732 9.3
R41973 vdd.n13829 vdd.n13828 9.3
R41974 vdd.n13829 vdd.n8733 9.3
R41975 vdd.n8738 vdd.n8733 9.3
R41976 vdd.n13845 vdd.n13844 9.3
R41977 vdd.n13854 vdd.n13853 9.3
R41978 vdd.n13855 vdd.n13854 9.3
R41979 vdd.n13856 vdd.n13855 9.3
R41980 vdd.n13895 vdd.n13894 9.3
R41981 vdd.n13892 vdd.n13891 9.3
R41982 vdd.n13891 vdd.n13890 9.3
R41983 vdd.n13890 vdd.n13889 9.3
R41984 vdd.n13911 vdd.n13910 9.3
R41985 vdd.n13914 vdd.n13913 9.3
R41986 vdd.n13915 vdd.n13914 9.3
R41987 vdd.n13977 vdd.n8613 9.3
R41988 vdd.n13977 vdd.n13976 9.3
R41989 vdd.n13982 vdd.n13981 9.3
R41990 vdd.n8610 vdd.n8602 9.3
R41991 vdd.n8602 vdd.n8601 9.3
R41992 vdd.n13988 vdd.n13986 9.3
R41993 vdd.n13988 vdd.n13987 9.3
R41994 vdd.n13987 vdd.n8588 9.3
R41995 vdd.n8605 vdd.n8570 9.3
R41996 vdd.n14059 vdd.n14058 9.3
R41997 vdd.n14059 vdd.n8567 9.3
R41998 vdd.n8567 vdd.n8565 9.3
R41999 vdd.n14048 vdd.n8571 9.3
R42000 vdd.n14049 vdd.n14048 9.3
R42001 vdd.n14050 vdd.n14049 9.3
R42002 vdd.n14045 vdd.n14042 9.3
R42003 vdd.n14044 vdd.n8559 9.3
R42004 vdd.n14070 vdd.n8559 9.3
R42005 vdd.n14070 vdd.n14069 9.3
R42006 vdd.n14076 vdd.n14075 9.3
R42007 vdd.n14077 vdd.n14076 9.3
R42008 vdd.n14078 vdd.n14077 9.3
R42009 vdd.n14115 vdd.n14114 9.3
R42010 vdd.n14115 vdd.n8514 9.3
R42011 vdd.n8535 vdd.n8514 9.3
R42012 vdd.n14111 vdd.n14110 9.3
R42013 vdd.n14110 vdd.n14109 9.3
R42014 vdd.n14109 vdd.n14108 9.3
R42015 vdd.n14134 vdd.n14133 9.3
R42016 vdd.n14143 vdd.n14142 9.3
R42017 vdd.n14144 vdd.n14143 9.3
R42018 vdd.n14145 vdd.n14144 9.3
R42019 vdd.n14184 vdd.n14183 9.3
R42020 vdd.n14181 vdd.n14180 9.3
R42021 vdd.n14180 vdd.n14179 9.3
R42022 vdd.n14179 vdd.n14178 9.3
R42023 vdd.n14201 vdd.n14200 9.3
R42024 vdd.n14204 vdd.n14203 9.3
R42025 vdd.n14205 vdd.n14204 9.3
R42026 vdd.n14267 vdd.n8391 9.3
R42027 vdd.n14267 vdd.n14266 9.3
R42028 vdd.n14272 vdd.n14271 9.3
R42029 vdd.n8388 vdd.n8380 9.3
R42030 vdd.n8380 vdd.n8379 9.3
R42031 vdd.n14279 vdd.n14276 9.3
R42032 vdd.n14279 vdd.n14278 9.3
R42033 vdd.n14278 vdd.n14277 9.3
R42034 vdd.n8383 vdd.n8353 9.3
R42035 vdd.n14334 vdd.n14333 9.3
R42036 vdd.n14334 vdd.n8349 9.3
R42037 vdd.n8349 vdd.n8347 9.3
R42038 vdd.n14322 vdd.n14321 9.3
R42039 vdd.n14350 vdd.n14349 9.3
R42040 vdd.n14352 vdd.n8338 9.3
R42041 vdd.n14424 vdd.n8278 9.3
R42042 vdd.n8246 vdd.n8244 9.3
R42043 vdd.n14455 vdd.n8247 9.3
R42044 vdd.n8256 vdd.n8255 9.3
R42045 vdd.n14493 vdd.n8218 9.3
R42046 vdd.n14936 vdd.n8003 9.3
R42047 vdd.n14917 vdd.n8013 9.3
R42048 vdd.n14902 vdd.n14901 9.3
R42049 vdd.n14866 vdd.n14865 9.3
R42050 vdd.n14866 vdd.n8037 9.3
R42051 vdd.n8037 vdd.n8035 9.3
R42052 vdd.n14838 vdd.n14837 9.3
R42053 vdd.n14837 vdd.n8045 9.3
R42054 vdd.n8045 vdd.n8044 9.3
R42055 vdd.n14825 vdd.n14824 9.3
R42056 vdd.n14825 vdd.n8057 9.3
R42057 vdd.n8057 vdd.n8055 9.3
R42058 vdd.n8077 vdd.n8065 9.3
R42059 vdd.n8065 vdd.n8064 9.3
R42060 vdd.n14769 vdd.n14768 9.3
R42061 vdd.n14753 vdd.n14752 9.3
R42062 vdd.n14737 vdd.n14736 9.3
R42063 vdd.n14681 vdd.n14680 9.3
R42064 vdd.n14681 vdd.n8118 9.3
R42065 vdd.n8119 vdd.n8118 9.3
R42066 vdd.n14676 vdd.n8132 9.3
R42067 vdd.n14676 vdd.n14675 9.3
R42068 vdd.n14675 vdd.n14674 9.3
R42069 vdd.n8158 vdd.n8152 9.3
R42070 vdd.n8159 vdd.n8158 9.3
R42071 vdd.n8160 vdd.n8159 9.3
R42072 vdd.n14653 vdd.n14652 9.3
R42073 vdd.n14653 vdd.n8148 9.3
R42074 vdd.n8148 vdd.n8146 9.3
R42075 vdd.n14650 vdd.n14649 9.3
R42076 vdd.n14651 vdd.n8150 9.3
R42077 vdd.n8157 vdd.n8156 9.3
R42078 vdd.n8155 vdd.n8137 9.3
R42079 vdd.n14666 vdd.n14665 9.3
R42080 vdd.n14665 vdd.n8135 9.3
R42081 vdd.n8141 vdd.n8135 9.3
R42082 vdd.n14669 vdd.n14668 9.3
R42083 vdd.n14667 vdd.n8136 9.3
R42084 vdd.n14677 vdd.n8130 9.3
R42085 vdd.n14679 vdd.n14678 9.3
R42086 vdd.n14692 vdd.n14691 9.3
R42087 vdd.n14692 vdd.n8127 9.3
R42088 vdd.n8127 vdd.n8125 9.3
R42089 vdd.n14689 vdd.n14688 9.3
R42090 vdd.n14690 vdd.n8129 9.3
R42091 vdd.n14710 vdd.n14709 9.3
R42092 vdd.n14711 vdd.n14710 9.3
R42093 vdd.n14712 vdd.n14711 9.3
R42094 vdd.n14717 vdd.n8110 9.3
R42095 vdd.n14720 vdd.n8108 9.3
R42096 vdd.n8108 vdd.n8106 9.3
R42097 vdd.n8106 vdd.n8104 9.3
R42098 vdd.n14719 vdd.n14718 9.3
R42099 vdd.n14735 vdd.n8109 9.3
R42100 vdd.n14734 vdd.n14733 9.3
R42101 vdd.n14733 vdd.n14732 9.3
R42102 vdd.n14732 vdd.n14731 9.3
R42103 vdd.n14726 vdd.n14721 9.3
R42104 vdd.n8098 vdd.n8097 9.3
R42105 vdd.n8099 vdd.n8098 9.3
R42106 vdd.n8100 vdd.n8099 9.3
R42107 vdd.n14725 vdd.n14724 9.3
R42108 vdd.n14754 vdd.n8096 9.3
R42109 vdd.n14756 vdd.n14755 9.3
R42110 vdd.n14757 vdd.n14756 9.3
R42111 vdd.n14758 vdd.n14757 9.3
R42112 vdd.n14763 vdd.n8091 9.3
R42113 vdd.n14766 vdd.n8086 9.3
R42114 vdd.n8086 vdd.n8084 9.3
R42115 vdd.n8084 vdd.n8082 9.3
R42116 vdd.n14765 vdd.n14764 9.3
R42117 vdd.n14767 vdd.n8090 9.3
R42118 vdd.n8089 vdd.n8068 9.3
R42119 vdd.n8089 vdd.n8088 9.3
R42120 vdd.n8088 vdd.n8087 9.3
R42121 vdd.n14793 vdd.n14792 9.3
R42122 vdd.n8076 vdd.n8071 9.3
R42123 vdd.n14788 vdd.n8071 9.3
R42124 vdd.n14797 vdd.n14796 9.3
R42125 vdd.n14804 vdd.n8062 9.3
R42126 vdd.n14804 vdd.n14803 9.3
R42127 vdd.n14803 vdd.n14802 9.3
R42128 vdd.n14807 vdd.n14806 9.3
R42129 vdd.n14805 vdd.n8060 9.3
R42130 vdd.n14823 vdd.n8059 9.3
R42131 vdd.n14822 vdd.n14821 9.3
R42132 vdd.n14814 vdd.n14808 9.3
R42133 vdd.n14815 vdd.n14814 9.3
R42134 vdd.n14816 vdd.n14815 9.3
R42135 vdd.n14811 vdd.n8047 9.3
R42136 vdd.n14813 vdd.n14812 9.3
R42137 vdd.n14839 vdd.n8046 9.3
R42138 vdd.n14841 vdd.n14840 9.3
R42139 vdd.n14848 vdd.n8042 9.3
R42140 vdd.n14848 vdd.n14847 9.3
R42141 vdd.n14847 vdd.n14846 9.3
R42142 vdd.n14851 vdd.n14850 9.3
R42143 vdd.n14849 vdd.n8040 9.3
R42144 vdd.n14864 vdd.n8039 9.3
R42145 vdd.n14863 vdd.n14862 9.3
R42146 vdd.n14855 vdd.n14852 9.3
R42147 vdd.n14856 vdd.n14855 9.3
R42148 vdd.n14856 vdd.n8030 9.3
R42149 vdd.n14882 vdd.n8024 9.3
R42150 vdd.n8024 vdd.n8022 9.3
R42151 vdd.n8022 vdd.n8020 9.3
R42152 vdd.n14900 vdd.n8025 9.3
R42153 vdd.n14899 vdd.n14898 9.3
R42154 vdd.n14898 vdd.n14897 9.3
R42155 vdd.n14897 vdd.n14896 9.3
R42156 vdd.n14891 vdd.n14883 9.3
R42157 vdd.n14888 vdd.n14887 9.3
R42158 vdd.n14887 vdd.n14886 9.3
R42159 vdd.n14886 vdd.n8016 9.3
R42160 vdd.n14890 vdd.n14889 9.3
R42161 vdd.n14919 vdd.n14918 9.3
R42162 vdd.n14920 vdd.n8012 9.3
R42163 vdd.n8012 vdd.n8011 9.3
R42164 vdd.n8011 vdd.n8009 9.3
R42165 vdd.n14922 vdd.n14921 9.3
R42166 vdd.n14935 vdd.n14934 9.3
R42167 vdd.n14934 vdd.n14933 9.3
R42168 vdd.n14933 vdd.n14932 9.3
R42169 vdd.n8005 vdd.n8004 9.3
R42170 vdd.n14938 vdd.n14937 9.3
R42171 vdd.n14939 vdd.n7982 9.3
R42172 vdd.n14939 vdd.n8002 9.3
R42173 vdd.n8002 vdd.n8001 9.3
R42174 vdd.n14496 vdd.n14495 9.3
R42175 vdd.n14496 vdd.n8217 9.3
R42176 vdd.n8223 vdd.n8217 9.3
R42177 vdd.n14492 vdd.n14491 9.3
R42178 vdd.n14454 vdd.n8250 9.3
R42179 vdd.n14454 vdd.n14453 9.3
R42180 vdd.n14453 vdd.n14452 9.3
R42181 vdd.n14457 vdd.n14456 9.3
R42182 vdd.n14423 vdd.n14422 9.3
R42183 vdd.n14422 vdd.n14421 9.3
R42184 vdd.n14421 vdd.n14420 9.3
R42185 vdd.n14426 vdd.n14425 9.3
R42186 vdd.n14351 vdd.n8336 9.3
R42187 vdd.n14323 vdd.n8354 9.3
R42188 vdd.n14324 vdd.n14323 9.3
R42189 vdd.n14325 vdd.n14324 9.3
R42190 vdd.n14320 vdd.n14319 9.3
R42191 vdd.n14348 vdd.n8339 9.3
R42192 vdd.n14348 vdd.n8334 9.3
R42193 vdd.n8334 vdd.n8327 9.3
R42194 vdd.n14356 vdd.n14353 9.3
R42195 vdd.n14356 vdd.n14355 9.3
R42196 vdd.n14355 vdd.n14354 9.3
R42197 vdd.n8337 vdd.n8300 9.3
R42198 vdd.n14400 vdd.n14399 9.3
R42199 vdd.n14399 vdd.n8298 9.3
R42200 vdd.n14395 vdd.n8298 9.3
R42201 vdd.n8279 vdd.n8277 9.3
R42202 vdd.n8277 vdd.n8275 9.3
R42203 vdd.n14408 vdd.n8275 9.3
R42204 vdd.n8281 vdd.n8280 9.3
R42205 vdd.n14459 vdd.n14458 9.3
R42206 vdd.n14460 vdd.n14459 9.3
R42207 vdd.n14461 vdd.n14460 9.3
R42208 vdd.n8258 vdd.n8257 9.3
R42209 vdd.n8254 vdd.n8219 9.3
R42210 vdd.n8254 vdd.n8253 9.3
R42211 vdd.n8253 vdd.n8234 9.3
R42212 vdd.n22136 vdd.n22135 9.3
R42213 vdd.n22110 vdd.n22109 9.3
R42214 vdd.n22073 vdd.n22072 9.3
R42215 vdd.n22057 vdd.n22056 9.3
R42216 vdd.n22334 vdd.n22333 9.3
R42217 vdd.n22234 vdd.n22233 9.3
R42218 vdd.n22209 vdd.n22208 9.3
R42219 vdd.n22199 vdd.n22198 9.3
R42220 vdd.n22362 vdd.n22361 9.3
R42221 vdd.n22361 vdd.n22360 9.3
R42222 vdd.n22360 vdd.n22359 9.3
R42223 vdd.n22239 vdd.n22238 9.3
R42224 vdd.n22227 vdd.n22226 9.3
R42225 vdd.n22226 vdd.n22225 9.3
R42226 vdd.n22339 vdd.n22338 9.3
R42227 vdd.n22253 vdd.n22252 9.3
R42228 vdd.n22252 vdd.n22251 9.3
R42229 vdd.n22141 vdd.n22140 9.3
R42230 vdd.n22129 vdd.n22128 9.3
R42231 vdd.n22128 vdd.n22127 9.3
R42232 vdd.n22115 vdd.n22114 9.3
R42233 vdd.n22103 vdd.n22102 9.3
R42234 vdd.n22102 vdd.n22101 9.3
R42235 vdd.n22091 vdd.n22090 9.3
R42236 vdd.n22090 vdd.n22089 9.3
R42237 vdd.n22089 vdd.n22088 9.3
R42238 vdd.n22278 vdd.n22277 9.3
R42239 vdd.n22277 vdd.n22276 9.3
R42240 vdd.n22304 vdd.n22303 9.3
R42241 vdd.n22303 vdd.n22302 9.3
R42242 vdd.n24363 vdd.n24362 9.3
R42243 vdd.n24362 vdd.n24361 9.3
R42244 vdd.n24337 vdd.n24336 9.3
R42245 vdd.n24336 vdd.n24335 9.3
R42246 vdd.n24335 vdd.n24334 9.3
R42247 vdd.n22052 vdd.n22051 9.3
R42248 vdd.n22051 vdd.n22050 9.3
R42249 vdd.n24348 vdd.n24347 9.3
R42250 vdd.n24347 vdd.n24346 9.3
R42251 vdd.n22289 vdd.n22288 9.3
R42252 vdd.n22288 vdd.n22287 9.3
R42253 vdd.n22311 vdd.n22310 9.3
R42254 vdd.n22320 vdd.n22319 9.3
R42255 vdd.n22319 vdd.n22318 9.3
R42256 vdd.n22267 vdd.n22266 9.3
R42257 vdd.n22266 vdd.n22265 9.3
R42258 vdd.n22163 vdd.n22162 9.3
R42259 vdd.n22162 vdd.n22161 9.3
R42260 vdd.n24276 vdd.n24275 9.3
R42261 vdd.n24275 vdd.n24274 9.3
R42262 vdd.n24246 vdd.n24245 9.3
R42263 vdd.n24245 vdd.n24244 9.3
R42264 vdd.n24220 vdd.n24219 9.3
R42265 vdd.n24219 vdd.n24218 9.3
R42266 vdd.n24218 vdd.n24217 9.3
R42267 vdd.n22173 vdd.n22172 9.3
R42268 vdd.n22172 vdd.n22171 9.3
R42269 vdd.n24231 vdd.n24230 9.3
R42270 vdd.n24230 vdd.n24229 9.3
R42271 vdd.n24261 vdd.n24260 9.3
R42272 vdd.n24260 vdd.n24259 9.3
R42273 vdd.n24283 vdd.n24282 9.3
R42274 vdd.n24292 vdd.n24291 9.3
R42275 vdd.n24291 vdd.n24290 9.3
R42276 vdd.n22152 vdd.n22151 9.3
R42277 vdd.n22151 vdd.n22150 9.3
R42278 vdd.n24202 vdd.n24201 9.3
R42279 vdd.n24201 vdd.n24200 9.3
R42280 vdd.n24200 vdd.n24199 9.3
R42281 vdd.n24176 vdd.n24175 9.3
R42282 vdd.n24190 vdd.n24189 9.3
R42283 vdd.n24192 vdd.n24191 9.3
R42284 vdd.n24164 vdd.n24163 9.3
R42285 vdd.n24150 vdd.n24149 9.3
R42286 vdd.n24136 vdd.n24135 9.3
R42287 vdd.n24122 vdd.n24121 9.3
R42288 vdd.n24108 vdd.n24107 9.3
R42289 vdd.n24094 vdd.n24093 9.3
R42290 vdd.n24080 vdd.n24079 9.3
R42291 vdd.n24066 vdd.n24065 9.3
R42292 vdd.n24052 vdd.n24051 9.3
R42293 vdd.n24038 vdd.n24037 9.3
R42294 vdd.n24024 vdd.n24023 9.3
R42295 vdd.n24010 vdd.n24009 9.3
R42296 vdd.n23996 vdd.n23995 9.3
R42297 vdd.n23982 vdd.n23981 9.3
R42298 vdd.n23960 vdd.n23959 9.3
R42299 vdd.n23946 vdd.n23945 9.3
R42300 vdd.n23932 vdd.n23931 9.3
R42301 vdd.n23918 vdd.n23917 9.3
R42302 vdd.n23904 vdd.n23903 9.3
R42303 vdd.n23890 vdd.n23889 9.3
R42304 vdd.n23876 vdd.n23875 9.3
R42305 vdd.n23862 vdd.n23861 9.3
R42306 vdd.n23848 vdd.n23847 9.3
R42307 vdd.n23834 vdd.n23833 9.3
R42308 vdd.n23820 vdd.n23819 9.3
R42309 vdd.n23806 vdd.n23805 9.3
R42310 vdd.n23792 vdd.n23791 9.3
R42311 vdd.n23778 vdd.n23777 9.3
R42312 vdd.n23764 vdd.n23763 9.3
R42313 vdd.n23750 vdd.n23749 9.3
R42314 vdd.n23728 vdd.n23727 9.3
R42315 vdd.n23714 vdd.n23713 9.3
R42316 vdd.n23700 vdd.n23699 9.3
R42317 vdd.n23686 vdd.n23685 9.3
R42318 vdd.n23672 vdd.n23671 9.3
R42319 vdd.n23658 vdd.n23657 9.3
R42320 vdd.n23644 vdd.n23643 9.3
R42321 vdd.n23640 vdd.n23639 9.3
R42322 vdd.n23639 vdd.n23638 9.3
R42323 vdd.n23638 vdd.n23637 9.3
R42324 vdd.n23748 vdd.n23747 9.3
R42325 vdd.n23747 vdd.n23746 9.3
R42326 vdd.n23746 vdd.n23745 9.3
R42327 vdd.n23776 vdd.n23775 9.3
R42328 vdd.n23775 vdd.n23774 9.3
R42329 vdd.n23774 vdd.n23773 9.3
R42330 vdd.n23804 vdd.n23803 9.3
R42331 vdd.n23803 vdd.n23802 9.3
R42332 vdd.n23802 vdd.n23801 9.3
R42333 vdd.n23832 vdd.n23831 9.3
R42334 vdd.n23831 vdd.n23830 9.3
R42335 vdd.n23830 vdd.n23829 9.3
R42336 vdd.n23980 vdd.n23979 9.3
R42337 vdd.n23979 vdd.n23978 9.3
R42338 vdd.n23978 vdd.n23977 9.3
R42339 vdd.n24008 vdd.n24007 9.3
R42340 vdd.n24007 vdd.n24006 9.3
R42341 vdd.n24006 vdd.n24005 9.3
R42342 vdd.n24036 vdd.n24035 9.3
R42343 vdd.n24035 vdd.n24034 9.3
R42344 vdd.n24034 vdd.n24033 9.3
R42345 vdd.n24064 vdd.n24063 9.3
R42346 vdd.n24063 vdd.n24062 9.3
R42347 vdd.n24062 vdd.n24061 9.3
R42348 vdd.n24162 vdd.n24161 9.3
R42349 vdd.n24174 vdd.n24173 9.3
R42350 vdd.n24173 vdd.n24172 9.3
R42351 vdd.n24172 vdd.n24171 9.3
R42352 vdd.n24160 vdd.n24159 9.3
R42353 vdd.n24159 vdd.n24158 9.3
R42354 vdd.n24158 vdd.n24157 9.3
R42355 vdd.n24148 vdd.n24147 9.3
R42356 vdd.n24134 vdd.n24133 9.3
R42357 vdd.n24146 vdd.n24145 9.3
R42358 vdd.n24145 vdd.n24144 9.3
R42359 vdd.n24144 vdd.n24143 9.3
R42360 vdd.n24132 vdd.n24131 9.3
R42361 vdd.n24131 vdd.n24130 9.3
R42362 vdd.n24130 vdd.n24129 9.3
R42363 vdd.n24120 vdd.n24119 9.3
R42364 vdd.n24106 vdd.n24105 9.3
R42365 vdd.n24118 vdd.n24117 9.3
R42366 vdd.n24117 vdd.n24116 9.3
R42367 vdd.n24116 vdd.n24115 9.3
R42368 vdd.n24104 vdd.n24103 9.3
R42369 vdd.n24103 vdd.n24102 9.3
R42370 vdd.n24102 vdd.n24101 9.3
R42371 vdd.n24092 vdd.n24091 9.3
R42372 vdd.n24082 vdd.n24081 9.3
R42373 vdd.n24078 vdd.n24077 9.3
R42374 vdd.n24077 vdd.n24076 9.3
R42375 vdd.n24076 vdd.n24075 9.3
R42376 vdd.n24068 vdd.n24067 9.3
R42377 vdd.n24054 vdd.n24053 9.3
R42378 vdd.n24050 vdd.n24049 9.3
R42379 vdd.n24049 vdd.n24048 9.3
R42380 vdd.n24048 vdd.n24047 9.3
R42381 vdd.n24040 vdd.n24039 9.3
R42382 vdd.n24026 vdd.n24025 9.3
R42383 vdd.n24022 vdd.n24021 9.3
R42384 vdd.n24021 vdd.n24020 9.3
R42385 vdd.n24020 vdd.n24019 9.3
R42386 vdd.n24012 vdd.n24011 9.3
R42387 vdd.n23998 vdd.n23997 9.3
R42388 vdd.n23994 vdd.n23993 9.3
R42389 vdd.n23993 vdd.n23992 9.3
R42390 vdd.n23992 vdd.n23991 9.3
R42391 vdd.n23984 vdd.n23983 9.3
R42392 vdd.n23958 vdd.n23957 9.3
R42393 vdd.n23970 vdd.n23969 9.3
R42394 vdd.n23969 vdd.n23968 9.3
R42395 vdd.n23968 vdd.n23967 9.3
R42396 vdd.n23956 vdd.n23955 9.3
R42397 vdd.n23955 vdd.n23954 9.3
R42398 vdd.n23954 vdd.n23953 9.3
R42399 vdd.n23944 vdd.n23943 9.3
R42400 vdd.n23930 vdd.n23929 9.3
R42401 vdd.n23942 vdd.n23941 9.3
R42402 vdd.n23941 vdd.n23940 9.3
R42403 vdd.n23940 vdd.n23939 9.3
R42404 vdd.n23928 vdd.n23927 9.3
R42405 vdd.n23927 vdd.n23926 9.3
R42406 vdd.n23926 vdd.n23925 9.3
R42407 vdd.n23916 vdd.n23915 9.3
R42408 vdd.n23902 vdd.n23901 9.3
R42409 vdd.n23914 vdd.n23913 9.3
R42410 vdd.n23913 vdd.n23912 9.3
R42411 vdd.n23912 vdd.n23911 9.3
R42412 vdd.n23900 vdd.n23899 9.3
R42413 vdd.n23899 vdd.n23898 9.3
R42414 vdd.n23898 vdd.n23897 9.3
R42415 vdd.n23888 vdd.n23887 9.3
R42416 vdd.n23874 vdd.n23873 9.3
R42417 vdd.n23886 vdd.n23885 9.3
R42418 vdd.n23885 vdd.n23884 9.3
R42419 vdd.n23884 vdd.n23883 9.3
R42420 vdd.n23872 vdd.n23871 9.3
R42421 vdd.n23871 vdd.n23870 9.3
R42422 vdd.n23870 vdd.n23869 9.3
R42423 vdd.n23860 vdd.n23859 9.3
R42424 vdd.n23850 vdd.n23849 9.3
R42425 vdd.n23846 vdd.n23845 9.3
R42426 vdd.n23845 vdd.n23844 9.3
R42427 vdd.n23844 vdd.n23843 9.3
R42428 vdd.n23836 vdd.n23835 9.3
R42429 vdd.n23822 vdd.n23821 9.3
R42430 vdd.n23818 vdd.n23817 9.3
R42431 vdd.n23817 vdd.n23816 9.3
R42432 vdd.n23816 vdd.n23815 9.3
R42433 vdd.n23808 vdd.n23807 9.3
R42434 vdd.n23794 vdd.n23793 9.3
R42435 vdd.n23790 vdd.n23789 9.3
R42436 vdd.n23789 vdd.n23788 9.3
R42437 vdd.n23788 vdd.n23787 9.3
R42438 vdd.n23780 vdd.n23779 9.3
R42439 vdd.n23766 vdd.n23765 9.3
R42440 vdd.n23762 vdd.n23761 9.3
R42441 vdd.n23761 vdd.n23760 9.3
R42442 vdd.n23760 vdd.n23759 9.3
R42443 vdd.n23752 vdd.n23751 9.3
R42444 vdd.n23726 vdd.n23725 9.3
R42445 vdd.n23738 vdd.n23737 9.3
R42446 vdd.n23737 vdd.n23736 9.3
R42447 vdd.n23736 vdd.n23735 9.3
R42448 vdd.n23724 vdd.n23723 9.3
R42449 vdd.n23723 vdd.n23722 9.3
R42450 vdd.n23722 vdd.n23721 9.3
R42451 vdd.n23712 vdd.n23711 9.3
R42452 vdd.n23698 vdd.n23697 9.3
R42453 vdd.n23710 vdd.n23709 9.3
R42454 vdd.n23709 vdd.n23708 9.3
R42455 vdd.n23708 vdd.n23707 9.3
R42456 vdd.n23696 vdd.n23695 9.3
R42457 vdd.n23695 vdd.n23694 9.3
R42458 vdd.n23694 vdd.n23693 9.3
R42459 vdd.n23684 vdd.n23683 9.3
R42460 vdd.n23670 vdd.n23669 9.3
R42461 vdd.n23682 vdd.n23681 9.3
R42462 vdd.n23681 vdd.n23680 9.3
R42463 vdd.n23680 vdd.n23679 9.3
R42464 vdd.n23668 vdd.n23667 9.3
R42465 vdd.n23667 vdd.n23666 9.3
R42466 vdd.n23666 vdd.n23665 9.3
R42467 vdd.n23656 vdd.n23655 9.3
R42468 vdd.n23642 vdd.n23641 9.3
R42469 vdd.n23654 vdd.n23653 9.3
R42470 vdd.n23653 vdd.n23652 9.3
R42471 vdd.n23652 vdd.n23651 9.3
R42472 vdd.n23628 vdd.n23627 9.3
R42473 vdd.n23630 vdd.n23629 9.3
R42474 vdd.n24178 vdd.n24177 9.3
R42475 vdd.n24188 vdd.n24187 9.3
R42476 vdd.n24187 vdd.n24186 9.3
R42477 vdd.n24186 vdd.n24185 9.3
R42478 vdd.n23624 vdd.n23623 9.3
R42479 vdd.n23610 vdd.n23609 9.3
R42480 vdd.n23596 vdd.n23595 9.3
R42481 vdd.n23582 vdd.n23581 9.3
R42482 vdd.n23568 vdd.n23567 9.3
R42483 vdd.n23554 vdd.n23553 9.3
R42484 vdd.n23540 vdd.n23539 9.3
R42485 vdd.n23526 vdd.n23525 9.3
R42486 vdd.n23504 vdd.n23503 9.3
R42487 vdd.n23490 vdd.n23489 9.3
R42488 vdd.n23476 vdd.n23475 9.3
R42489 vdd.n23462 vdd.n23461 9.3
R42490 vdd.n23448 vdd.n23447 9.3
R42491 vdd.n23434 vdd.n23433 9.3
R42492 vdd.n23420 vdd.n23419 9.3
R42493 vdd.n23406 vdd.n23405 9.3
R42494 vdd.n23392 vdd.n23391 9.3
R42495 vdd.n23378 vdd.n23377 9.3
R42496 vdd.n23364 vdd.n23363 9.3
R42497 vdd.n23350 vdd.n23349 9.3
R42498 vdd.n23336 vdd.n23335 9.3
R42499 vdd.n23322 vdd.n23321 9.3
R42500 vdd.n23308 vdd.n23307 9.3
R42501 vdd.n23294 vdd.n23293 9.3
R42502 vdd.n23272 vdd.n23271 9.3
R42503 vdd.n23258 vdd.n23257 9.3
R42504 vdd.n23244 vdd.n23243 9.3
R42505 vdd.n23230 vdd.n23229 9.3
R42506 vdd.n23216 vdd.n23215 9.3
R42507 vdd.n23202 vdd.n23201 9.3
R42508 vdd.n23188 vdd.n23187 9.3
R42509 vdd.n23174 vdd.n23173 9.3
R42510 vdd.n23160 vdd.n23159 9.3
R42511 vdd.n23146 vdd.n23145 9.3
R42512 vdd.n23132 vdd.n23131 9.3
R42513 vdd.n23118 vdd.n23117 9.3
R42514 vdd.n23104 vdd.n23103 9.3
R42515 vdd.n23090 vdd.n23089 9.3
R42516 vdd.n23076 vdd.n23075 9.3
R42517 vdd.n23612 vdd.n23611 9.3
R42518 vdd.n23584 vdd.n23583 9.3
R42519 vdd.n23556 vdd.n23555 9.3
R42520 vdd.n23528 vdd.n23527 9.3
R42521 vdd.n23514 vdd.n23513 9.3
R42522 vdd.n23513 vdd.n23512 9.3
R42523 vdd.n23512 vdd.n23511 9.3
R42524 vdd.n23502 vdd.n23501 9.3
R42525 vdd.n23486 vdd.n23485 9.3
R42526 vdd.n23485 vdd.n23484 9.3
R42527 vdd.n23484 vdd.n23483 9.3
R42528 vdd.n23474 vdd.n23473 9.3
R42529 vdd.n23458 vdd.n23457 9.3
R42530 vdd.n23457 vdd.n23456 9.3
R42531 vdd.n23456 vdd.n23455 9.3
R42532 vdd.n23446 vdd.n23445 9.3
R42533 vdd.n23430 vdd.n23429 9.3
R42534 vdd.n23429 vdd.n23428 9.3
R42535 vdd.n23428 vdd.n23427 9.3
R42536 vdd.n23418 vdd.n23417 9.3
R42537 vdd.n23380 vdd.n23379 9.3
R42538 vdd.n23352 vdd.n23351 9.3
R42539 vdd.n23324 vdd.n23323 9.3
R42540 vdd.n23296 vdd.n23295 9.3
R42541 vdd.n23282 vdd.n23281 9.3
R42542 vdd.n23281 vdd.n23280 9.3
R42543 vdd.n23280 vdd.n23279 9.3
R42544 vdd.n23270 vdd.n23269 9.3
R42545 vdd.n23254 vdd.n23253 9.3
R42546 vdd.n23253 vdd.n23252 9.3
R42547 vdd.n23252 vdd.n23251 9.3
R42548 vdd.n23242 vdd.n23241 9.3
R42549 vdd.n23226 vdd.n23225 9.3
R42550 vdd.n23225 vdd.n23224 9.3
R42551 vdd.n23224 vdd.n23223 9.3
R42552 vdd.n23214 vdd.n23213 9.3
R42553 vdd.n23198 vdd.n23197 9.3
R42554 vdd.n23197 vdd.n23196 9.3
R42555 vdd.n23196 vdd.n23195 9.3
R42556 vdd.n23186 vdd.n23185 9.3
R42557 vdd.n23148 vdd.n23147 9.3
R42558 vdd.n23120 vdd.n23119 9.3
R42559 vdd.n23092 vdd.n23091 9.3
R42560 vdd.n23074 vdd.n23073 9.3
R42561 vdd.n23073 vdd.n23072 9.3
R42562 vdd.n23072 vdd.n23071 9.3
R42563 vdd.n23078 vdd.n23077 9.3
R42564 vdd.n23088 vdd.n23087 9.3
R42565 vdd.n23087 vdd.n23086 9.3
R42566 vdd.n23086 vdd.n23085 9.3
R42567 vdd.n23102 vdd.n23101 9.3
R42568 vdd.n23101 vdd.n23100 9.3
R42569 vdd.n23100 vdd.n23099 9.3
R42570 vdd.n23106 vdd.n23105 9.3
R42571 vdd.n23116 vdd.n23115 9.3
R42572 vdd.n23115 vdd.n23114 9.3
R42573 vdd.n23114 vdd.n23113 9.3
R42574 vdd.n23130 vdd.n23129 9.3
R42575 vdd.n23129 vdd.n23128 9.3
R42576 vdd.n23128 vdd.n23127 9.3
R42577 vdd.n23134 vdd.n23133 9.3
R42578 vdd.n23144 vdd.n23143 9.3
R42579 vdd.n23143 vdd.n23142 9.3
R42580 vdd.n23142 vdd.n23141 9.3
R42581 vdd.n23158 vdd.n23157 9.3
R42582 vdd.n23157 vdd.n23156 9.3
R42583 vdd.n23156 vdd.n23155 9.3
R42584 vdd.n23162 vdd.n23161 9.3
R42585 vdd.n23172 vdd.n23171 9.3
R42586 vdd.n23184 vdd.n23183 9.3
R42587 vdd.n23183 vdd.n23182 9.3
R42588 vdd.n23182 vdd.n23181 9.3
R42589 vdd.n23200 vdd.n23199 9.3
R42590 vdd.n23212 vdd.n23211 9.3
R42591 vdd.n23211 vdd.n23210 9.3
R42592 vdd.n23210 vdd.n23209 9.3
R42593 vdd.n23228 vdd.n23227 9.3
R42594 vdd.n23240 vdd.n23239 9.3
R42595 vdd.n23239 vdd.n23238 9.3
R42596 vdd.n23238 vdd.n23237 9.3
R42597 vdd.n23256 vdd.n23255 9.3
R42598 vdd.n23268 vdd.n23267 9.3
R42599 vdd.n23267 vdd.n23266 9.3
R42600 vdd.n23266 vdd.n23265 9.3
R42601 vdd.n23292 vdd.n23291 9.3
R42602 vdd.n23291 vdd.n23290 9.3
R42603 vdd.n23290 vdd.n23289 9.3
R42604 vdd.n23306 vdd.n23305 9.3
R42605 vdd.n23305 vdd.n23304 9.3
R42606 vdd.n23304 vdd.n23303 9.3
R42607 vdd.n23310 vdd.n23309 9.3
R42608 vdd.n23320 vdd.n23319 9.3
R42609 vdd.n23319 vdd.n23318 9.3
R42610 vdd.n23318 vdd.n23317 9.3
R42611 vdd.n23334 vdd.n23333 9.3
R42612 vdd.n23333 vdd.n23332 9.3
R42613 vdd.n23332 vdd.n23331 9.3
R42614 vdd.n23338 vdd.n23337 9.3
R42615 vdd.n23348 vdd.n23347 9.3
R42616 vdd.n23347 vdd.n23346 9.3
R42617 vdd.n23346 vdd.n23345 9.3
R42618 vdd.n23362 vdd.n23361 9.3
R42619 vdd.n23361 vdd.n23360 9.3
R42620 vdd.n23360 vdd.n23359 9.3
R42621 vdd.n23366 vdd.n23365 9.3
R42622 vdd.n23376 vdd.n23375 9.3
R42623 vdd.n23375 vdd.n23374 9.3
R42624 vdd.n23374 vdd.n23373 9.3
R42625 vdd.n23390 vdd.n23389 9.3
R42626 vdd.n23389 vdd.n23388 9.3
R42627 vdd.n23388 vdd.n23387 9.3
R42628 vdd.n23394 vdd.n23393 9.3
R42629 vdd.n23404 vdd.n23403 9.3
R42630 vdd.n23416 vdd.n23415 9.3
R42631 vdd.n23415 vdd.n23414 9.3
R42632 vdd.n23414 vdd.n23413 9.3
R42633 vdd.n23432 vdd.n23431 9.3
R42634 vdd.n23444 vdd.n23443 9.3
R42635 vdd.n23443 vdd.n23442 9.3
R42636 vdd.n23442 vdd.n23441 9.3
R42637 vdd.n23460 vdd.n23459 9.3
R42638 vdd.n23472 vdd.n23471 9.3
R42639 vdd.n23471 vdd.n23470 9.3
R42640 vdd.n23470 vdd.n23469 9.3
R42641 vdd.n23488 vdd.n23487 9.3
R42642 vdd.n23500 vdd.n23499 9.3
R42643 vdd.n23499 vdd.n23498 9.3
R42644 vdd.n23498 vdd.n23497 9.3
R42645 vdd.n23524 vdd.n23523 9.3
R42646 vdd.n23523 vdd.n23522 9.3
R42647 vdd.n23522 vdd.n23521 9.3
R42648 vdd.n23538 vdd.n23537 9.3
R42649 vdd.n23537 vdd.n23536 9.3
R42650 vdd.n23536 vdd.n23535 9.3
R42651 vdd.n23542 vdd.n23541 9.3
R42652 vdd.n23552 vdd.n23551 9.3
R42653 vdd.n23551 vdd.n23550 9.3
R42654 vdd.n23550 vdd.n23549 9.3
R42655 vdd.n23566 vdd.n23565 9.3
R42656 vdd.n23565 vdd.n23564 9.3
R42657 vdd.n23564 vdd.n23563 9.3
R42658 vdd.n23570 vdd.n23569 9.3
R42659 vdd.n23580 vdd.n23579 9.3
R42660 vdd.n23579 vdd.n23578 9.3
R42661 vdd.n23578 vdd.n23577 9.3
R42662 vdd.n23594 vdd.n23593 9.3
R42663 vdd.n23593 vdd.n23592 9.3
R42664 vdd.n23592 vdd.n23591 9.3
R42665 vdd.n23598 vdd.n23597 9.3
R42666 vdd.n23608 vdd.n23607 9.3
R42667 vdd.n23607 vdd.n23606 9.3
R42668 vdd.n23606 vdd.n23605 9.3
R42669 vdd.n23622 vdd.n23621 9.3
R42670 vdd.n23621 vdd.n23620 9.3
R42671 vdd.n23620 vdd.n23619 9.3
R42672 vdd.n23626 vdd.n23625 9.3
R42673 vdd.n23060 vdd.n23059 9.3
R42674 vdd.n23059 vdd.n23058 9.3
R42675 vdd.n23058 vdd.n23057 9.3
R42676 vdd.n23064 vdd.n23063 9.3
R42677 vdd.n23062 vdd.n23061 9.3
R42678 vdd.n22483 vdd.n22482 9.3
R42679 vdd.n22497 vdd.n22496 9.3
R42680 vdd.n22511 vdd.n22510 9.3
R42681 vdd.n22525 vdd.n22524 9.3
R42682 vdd.n22539 vdd.n22538 9.3
R42683 vdd.n22553 vdd.n22552 9.3
R42684 vdd.n22567 vdd.n22566 9.3
R42685 vdd.n22581 vdd.n22580 9.3
R42686 vdd.n22595 vdd.n22594 9.3
R42687 vdd.n22609 vdd.n22608 9.3
R42688 vdd.n22623 vdd.n22622 9.3
R42689 vdd.n22637 vdd.n22636 9.3
R42690 vdd.n22651 vdd.n22650 9.3
R42691 vdd.n22665 vdd.n22664 9.3
R42692 vdd.n22679 vdd.n22678 9.3
R42693 vdd.n22693 vdd.n22692 9.3
R42694 vdd.n22715 vdd.n22714 9.3
R42695 vdd.n22729 vdd.n22728 9.3
R42696 vdd.n22743 vdd.n22742 9.3
R42697 vdd.n22757 vdd.n22756 9.3
R42698 vdd.n22771 vdd.n22770 9.3
R42699 vdd.n22785 vdd.n22784 9.3
R42700 vdd.n22799 vdd.n22798 9.3
R42701 vdd.n22813 vdd.n22812 9.3
R42702 vdd.n22827 vdd.n22826 9.3
R42703 vdd.n22841 vdd.n22840 9.3
R42704 vdd.n22855 vdd.n22854 9.3
R42705 vdd.n22869 vdd.n22868 9.3
R42706 vdd.n22883 vdd.n22882 9.3
R42707 vdd.n22897 vdd.n22896 9.3
R42708 vdd.n22911 vdd.n22910 9.3
R42709 vdd.n22925 vdd.n22924 9.3
R42710 vdd.n22947 vdd.n22946 9.3
R42711 vdd.n22961 vdd.n22960 9.3
R42712 vdd.n22975 vdd.n22974 9.3
R42713 vdd.n22989 vdd.n22988 9.3
R42714 vdd.n23003 vdd.n23002 9.3
R42715 vdd.n23017 vdd.n23016 9.3
R42716 vdd.n23031 vdd.n23030 9.3
R42717 vdd.n23045 vdd.n23044 9.3
R42718 vdd.n22935 vdd.n22934 9.3
R42719 vdd.n22934 vdd.n22933 9.3
R42720 vdd.n22933 vdd.n22932 9.3
R42721 vdd.n22907 vdd.n22906 9.3
R42722 vdd.n22906 vdd.n22905 9.3
R42723 vdd.n22905 vdd.n22904 9.3
R42724 vdd.n22879 vdd.n22878 9.3
R42725 vdd.n22878 vdd.n22877 9.3
R42726 vdd.n22877 vdd.n22876 9.3
R42727 vdd.n22851 vdd.n22850 9.3
R42728 vdd.n22850 vdd.n22849 9.3
R42729 vdd.n22849 vdd.n22848 9.3
R42730 vdd.n22703 vdd.n22702 9.3
R42731 vdd.n22702 vdd.n22701 9.3
R42732 vdd.n22701 vdd.n22700 9.3
R42733 vdd.n22675 vdd.n22674 9.3
R42734 vdd.n22674 vdd.n22673 9.3
R42735 vdd.n22673 vdd.n22672 9.3
R42736 vdd.n22647 vdd.n22646 9.3
R42737 vdd.n22646 vdd.n22645 9.3
R42738 vdd.n22645 vdd.n22644 9.3
R42739 vdd.n22619 vdd.n22618 9.3
R42740 vdd.n22618 vdd.n22617 9.3
R42741 vdd.n22617 vdd.n22616 9.3
R42742 vdd.n22485 vdd.n22484 9.3
R42743 vdd.n22481 vdd.n22480 9.3
R42744 vdd.n22480 vdd.n22479 9.3
R42745 vdd.n22479 vdd.n22478 9.3
R42746 vdd.n22495 vdd.n22494 9.3
R42747 vdd.n22494 vdd.n22493 9.3
R42748 vdd.n22493 vdd.n22492 9.3
R42749 vdd.n22499 vdd.n22498 9.3
R42750 vdd.n22513 vdd.n22512 9.3
R42751 vdd.n22509 vdd.n22508 9.3
R42752 vdd.n22508 vdd.n22507 9.3
R42753 vdd.n22507 vdd.n22506 9.3
R42754 vdd.n22523 vdd.n22522 9.3
R42755 vdd.n22522 vdd.n22521 9.3
R42756 vdd.n22521 vdd.n22520 9.3
R42757 vdd.n22527 vdd.n22526 9.3
R42758 vdd.n22541 vdd.n22540 9.3
R42759 vdd.n22537 vdd.n22536 9.3
R42760 vdd.n22536 vdd.n22535 9.3
R42761 vdd.n22535 vdd.n22534 9.3
R42762 vdd.n22551 vdd.n22550 9.3
R42763 vdd.n22550 vdd.n22549 9.3
R42764 vdd.n22549 vdd.n22548 9.3
R42765 vdd.n22555 vdd.n22554 9.3
R42766 vdd.n22569 vdd.n22568 9.3
R42767 vdd.n22565 vdd.n22564 9.3
R42768 vdd.n22564 vdd.n22563 9.3
R42769 vdd.n22563 vdd.n22562 9.3
R42770 vdd.n22579 vdd.n22578 9.3
R42771 vdd.n22578 vdd.n22577 9.3
R42772 vdd.n22577 vdd.n22576 9.3
R42773 vdd.n22583 vdd.n22582 9.3
R42774 vdd.n22593 vdd.n22592 9.3
R42775 vdd.n22605 vdd.n22604 9.3
R42776 vdd.n22604 vdd.n22603 9.3
R42777 vdd.n22603 vdd.n22602 9.3
R42778 vdd.n22607 vdd.n22606 9.3
R42779 vdd.n22621 vdd.n22620 9.3
R42780 vdd.n22633 vdd.n22632 9.3
R42781 vdd.n22632 vdd.n22631 9.3
R42782 vdd.n22631 vdd.n22630 9.3
R42783 vdd.n22635 vdd.n22634 9.3
R42784 vdd.n22649 vdd.n22648 9.3
R42785 vdd.n22661 vdd.n22660 9.3
R42786 vdd.n22660 vdd.n22659 9.3
R42787 vdd.n22659 vdd.n22658 9.3
R42788 vdd.n22663 vdd.n22662 9.3
R42789 vdd.n22677 vdd.n22676 9.3
R42790 vdd.n22689 vdd.n22688 9.3
R42791 vdd.n22688 vdd.n22687 9.3
R42792 vdd.n22687 vdd.n22686 9.3
R42793 vdd.n22691 vdd.n22690 9.3
R42794 vdd.n22717 vdd.n22716 9.3
R42795 vdd.n22713 vdd.n22712 9.3
R42796 vdd.n22712 vdd.n22711 9.3
R42797 vdd.n22711 vdd.n22710 9.3
R42798 vdd.n22727 vdd.n22726 9.3
R42799 vdd.n22726 vdd.n22725 9.3
R42800 vdd.n22725 vdd.n22724 9.3
R42801 vdd.n22731 vdd.n22730 9.3
R42802 vdd.n22745 vdd.n22744 9.3
R42803 vdd.n22741 vdd.n22740 9.3
R42804 vdd.n22740 vdd.n22739 9.3
R42805 vdd.n22739 vdd.n22738 9.3
R42806 vdd.n22755 vdd.n22754 9.3
R42807 vdd.n22754 vdd.n22753 9.3
R42808 vdd.n22753 vdd.n22752 9.3
R42809 vdd.n22759 vdd.n22758 9.3
R42810 vdd.n22773 vdd.n22772 9.3
R42811 vdd.n22769 vdd.n22768 9.3
R42812 vdd.n22768 vdd.n22767 9.3
R42813 vdd.n22767 vdd.n22766 9.3
R42814 vdd.n22783 vdd.n22782 9.3
R42815 vdd.n22782 vdd.n22781 9.3
R42816 vdd.n22781 vdd.n22780 9.3
R42817 vdd.n22787 vdd.n22786 9.3
R42818 vdd.n22801 vdd.n22800 9.3
R42819 vdd.n22797 vdd.n22796 9.3
R42820 vdd.n22796 vdd.n22795 9.3
R42821 vdd.n22795 vdd.n22794 9.3
R42822 vdd.n22811 vdd.n22810 9.3
R42823 vdd.n22810 vdd.n22809 9.3
R42824 vdd.n22809 vdd.n22808 9.3
R42825 vdd.n22815 vdd.n22814 9.3
R42826 vdd.n22825 vdd.n22824 9.3
R42827 vdd.n22837 vdd.n22836 9.3
R42828 vdd.n22836 vdd.n22835 9.3
R42829 vdd.n22835 vdd.n22834 9.3
R42830 vdd.n22839 vdd.n22838 9.3
R42831 vdd.n22853 vdd.n22852 9.3
R42832 vdd.n22865 vdd.n22864 9.3
R42833 vdd.n22864 vdd.n22863 9.3
R42834 vdd.n22863 vdd.n22862 9.3
R42835 vdd.n22867 vdd.n22866 9.3
R42836 vdd.n22881 vdd.n22880 9.3
R42837 vdd.n22893 vdd.n22892 9.3
R42838 vdd.n22892 vdd.n22891 9.3
R42839 vdd.n22891 vdd.n22890 9.3
R42840 vdd.n22895 vdd.n22894 9.3
R42841 vdd.n22909 vdd.n22908 9.3
R42842 vdd.n22921 vdd.n22920 9.3
R42843 vdd.n22920 vdd.n22919 9.3
R42844 vdd.n22919 vdd.n22918 9.3
R42845 vdd.n22923 vdd.n22922 9.3
R42846 vdd.n22949 vdd.n22948 9.3
R42847 vdd.n22945 vdd.n22944 9.3
R42848 vdd.n22944 vdd.n22943 9.3
R42849 vdd.n22943 vdd.n22942 9.3
R42850 vdd.n22959 vdd.n22958 9.3
R42851 vdd.n22958 vdd.n22957 9.3
R42852 vdd.n22957 vdd.n22956 9.3
R42853 vdd.n22963 vdd.n22962 9.3
R42854 vdd.n22977 vdd.n22976 9.3
R42855 vdd.n22973 vdd.n22972 9.3
R42856 vdd.n22972 vdd.n22971 9.3
R42857 vdd.n22971 vdd.n22970 9.3
R42858 vdd.n22987 vdd.n22986 9.3
R42859 vdd.n22986 vdd.n22985 9.3
R42860 vdd.n22985 vdd.n22984 9.3
R42861 vdd.n22991 vdd.n22990 9.3
R42862 vdd.n23005 vdd.n23004 9.3
R42863 vdd.n23001 vdd.n23000 9.3
R42864 vdd.n23000 vdd.n22999 9.3
R42865 vdd.n22999 vdd.n22998 9.3
R42866 vdd.n23015 vdd.n23014 9.3
R42867 vdd.n23014 vdd.n23013 9.3
R42868 vdd.n23013 vdd.n23012 9.3
R42869 vdd.n23019 vdd.n23018 9.3
R42870 vdd.n23033 vdd.n23032 9.3
R42871 vdd.n23029 vdd.n23028 9.3
R42872 vdd.n23028 vdd.n23027 9.3
R42873 vdd.n23027 vdd.n23026 9.3
R42874 vdd.n23043 vdd.n23042 9.3
R42875 vdd.n23042 vdd.n23041 9.3
R42876 vdd.n23041 vdd.n23040 9.3
R42877 vdd.n23050 vdd.n23049 9.3
R42878 vdd.n22184 vdd.n22183 9.3
R42879 vdd.n22183 vdd.n22182 9.3
R42880 vdd.n22448 vdd.n22447 9.3
R42881 vdd.n22447 vdd.n22446 9.3
R42882 vdd.n22418 vdd.n22417 9.3
R42883 vdd.n22417 vdd.n22416 9.3
R42884 vdd.n22392 vdd.n22391 9.3
R42885 vdd.n22391 vdd.n22390 9.3
R42886 vdd.n22390 vdd.n22389 9.3
R42887 vdd.n22194 vdd.n22193 9.3
R42888 vdd.n22193 vdd.n22192 9.3
R42889 vdd.n22403 vdd.n22402 9.3
R42890 vdd.n22402 vdd.n22401 9.3
R42891 vdd.n22433 vdd.n22432 9.3
R42892 vdd.n22432 vdd.n22431 9.3
R42893 vdd.n22455 vdd.n22454 9.3
R42894 vdd.n22464 vdd.n22463 9.3
R42895 vdd.n22463 vdd.n22462 9.3
R42896 vdd.n15120 vdd.n15067 9.3
R42897 vdd.n15066 vdd.n15065 9.3
R42898 vdd.n15054 vdd.n15053 9.3
R42899 vdd.n15048 vdd.n15047 9.3
R42900 vdd.n16676 vdd.n16675 9.3
R42901 vdd.n16587 vdd.n16586 9.3
R42902 vdd.n16595 vdd.n16594 9.3
R42903 vdd.n16689 vdd.n16688 9.3
R42904 vdd.n16743 vdd.n16742 9.3
R42905 vdd.n16743 vdd.n16690 9.3
R42906 vdd.n21079 vdd.n21078 9.3
R42907 vdd.n21063 vdd.n21062 9.3
R42908 vdd.n21047 vdd.n21046 9.3
R42909 vdd.n21031 vdd.n21030 9.3
R42910 vdd.n21017 vdd.n21016 9.3
R42911 vdd.n19134 vdd.n19133 9.3
R42912 vdd.n19119 vdd.n19118 9.3
R42913 vdd.n19103 vdd.n19102 9.3
R42914 vdd.n19087 vdd.n19086 9.3
R42915 vdd.n19071 vdd.n19070 9.3
R42916 vdd.n19055 vdd.n19054 9.3
R42917 vdd.n19039 vdd.n19038 9.3
R42918 vdd.n19004 vdd.n19003 9.3
R42919 vdd.n18988 vdd.n18987 9.3
R42920 vdd.n18972 vdd.n18971 9.3
R42921 vdd.n18956 vdd.n18955 9.3
R42922 vdd.n18940 vdd.n18939 9.3
R42923 vdd.n18924 vdd.n18923 9.3
R42924 vdd.n18908 vdd.n18907 9.3
R42925 vdd.n18876 vdd.n18875 9.3
R42926 vdd.n18860 vdd.n18859 9.3
R42927 vdd.n18844 vdd.n18843 9.3
R42928 vdd.n18828 vdd.n18827 9.3
R42929 vdd.n18812 vdd.n18811 9.3
R42930 vdd.n18796 vdd.n18795 9.3
R42931 vdd.n18780 vdd.n18779 9.3
R42932 vdd.n18745 vdd.n18744 9.3
R42933 vdd.n18729 vdd.n18728 9.3
R42934 vdd.n18713 vdd.n18712 9.3
R42935 vdd.n18697 vdd.n18696 9.3
R42936 vdd.n18681 vdd.n18680 9.3
R42937 vdd.n18665 vdd.n18664 9.3
R42938 vdd.n18649 vdd.n18648 9.3
R42939 vdd.n18617 vdd.n18616 9.3
R42940 vdd.n18601 vdd.n18600 9.3
R42941 vdd.n18585 vdd.n18584 9.3
R42942 vdd.n18569 vdd.n18568 9.3
R42943 vdd.n18553 vdd.n18552 9.3
R42944 vdd.n18537 vdd.n18536 9.3
R42945 vdd.n18521 vdd.n18520 9.3
R42946 vdd.n18519 vdd.n18518 9.3
R42947 vdd.n18535 vdd.n18534 9.3
R42948 vdd.n18551 vdd.n18550 9.3
R42949 vdd.n18567 vdd.n18566 9.3
R42950 vdd.n18583 vdd.n18582 9.3
R42951 vdd.n18599 vdd.n18598 9.3
R42952 vdd.n18615 vdd.n18614 9.3
R42953 vdd.n18651 vdd.n18650 9.3
R42954 vdd.n18667 vdd.n18666 9.3
R42955 vdd.n18683 vdd.n18682 9.3
R42956 vdd.n18699 vdd.n18698 9.3
R42957 vdd.n18715 vdd.n18714 9.3
R42958 vdd.n18731 vdd.n18730 9.3
R42959 vdd.n18747 vdd.n18746 9.3
R42960 vdd.n18778 vdd.n18777 9.3
R42961 vdd.n18794 vdd.n18793 9.3
R42962 vdd.n18810 vdd.n18809 9.3
R42963 vdd.n18826 vdd.n18825 9.3
R42964 vdd.n18842 vdd.n18841 9.3
R42965 vdd.n18858 vdd.n18857 9.3
R42966 vdd.n18874 vdd.n18873 9.3
R42967 vdd.n18910 vdd.n18909 9.3
R42968 vdd.n18926 vdd.n18925 9.3
R42969 vdd.n18942 vdd.n18941 9.3
R42970 vdd.n18958 vdd.n18957 9.3
R42971 vdd.n18974 vdd.n18973 9.3
R42972 vdd.n18990 vdd.n18989 9.3
R42973 vdd.n19006 vdd.n19005 9.3
R42974 vdd.n19037 vdd.n19036 9.3
R42975 vdd.n19053 vdd.n19052 9.3
R42976 vdd.n19069 vdd.n19068 9.3
R42977 vdd.n19085 vdd.n19084 9.3
R42978 vdd.n19101 vdd.n19100 9.3
R42979 vdd.n19117 vdd.n19116 9.3
R42980 vdd.n19132 vdd.n19131 9.3
R42981 vdd.n21019 vdd.n21018 9.3
R42982 vdd.n21033 vdd.n21032 9.3
R42983 vdd.n21049 vdd.n21048 9.3
R42984 vdd.n21065 vdd.n21064 9.3
R42985 vdd.n21687 vdd.n21686 9.3
R42986 vdd.n21623 vdd.n21622 9.3
R42987 vdd.n21597 vdd.n21596 9.3
R42988 vdd.n21581 vdd.n21580 9.3
R42989 vdd.n21565 vdd.n21564 9.3
R42990 vdd.n21549 vdd.n21548 9.3
R42991 vdd.n21533 vdd.n21532 9.3
R42992 vdd.n21501 vdd.n21500 9.3
R42993 vdd.n21485 vdd.n21484 9.3
R42994 vdd.n21469 vdd.n21468 9.3
R42995 vdd.n21453 vdd.n21452 9.3
R42996 vdd.n21437 vdd.n21436 9.3
R42997 vdd.n21421 vdd.n21420 9.3
R42998 vdd.n21405 vdd.n21404 9.3
R42999 vdd.n21370 vdd.n21369 9.3
R43000 vdd.n21354 vdd.n21353 9.3
R43001 vdd.n21338 vdd.n21337 9.3
R43002 vdd.n21322 vdd.n21321 9.3
R43003 vdd.n21306 vdd.n21305 9.3
R43004 vdd.n21290 vdd.n21289 9.3
R43005 vdd.n21274 vdd.n21273 9.3
R43006 vdd.n21242 vdd.n21241 9.3
R43007 vdd.n21226 vdd.n21225 9.3
R43008 vdd.n21210 vdd.n21209 9.3
R43009 vdd.n21194 vdd.n21193 9.3
R43010 vdd.n21178 vdd.n21177 9.3
R43011 vdd.n21162 vdd.n21161 9.3
R43012 vdd.n21146 vdd.n21145 9.3
R43013 vdd.n21111 vdd.n21110 9.3
R43014 vdd.n21095 vdd.n21094 9.3
R43015 vdd.n21621 vdd.n21620 9.3
R43016 vdd.n21092 vdd.n21091 9.3
R43017 vdd.n21097 vdd.n21096 9.3
R43018 vdd.n21113 vdd.n21112 9.3
R43019 vdd.n21144 vdd.n21143 9.3
R43020 vdd.n21160 vdd.n21159 9.3
R43021 vdd.n21176 vdd.n21175 9.3
R43022 vdd.n21192 vdd.n21191 9.3
R43023 vdd.n21208 vdd.n21207 9.3
R43024 vdd.n21224 vdd.n21223 9.3
R43025 vdd.n21240 vdd.n21239 9.3
R43026 vdd.n21276 vdd.n21275 9.3
R43027 vdd.n21292 vdd.n21291 9.3
R43028 vdd.n21308 vdd.n21307 9.3
R43029 vdd.n21324 vdd.n21323 9.3
R43030 vdd.n21340 vdd.n21339 9.3
R43031 vdd.n21356 vdd.n21355 9.3
R43032 vdd.n21372 vdd.n21371 9.3
R43033 vdd.n21403 vdd.n21402 9.3
R43034 vdd.n21419 vdd.n21418 9.3
R43035 vdd.n21435 vdd.n21434 9.3
R43036 vdd.n21451 vdd.n21450 9.3
R43037 vdd.n21467 vdd.n21466 9.3
R43038 vdd.n21483 vdd.n21482 9.3
R43039 vdd.n21499 vdd.n21498 9.3
R43040 vdd.n21535 vdd.n21534 9.3
R43041 vdd.n21551 vdd.n21550 9.3
R43042 vdd.n21567 vdd.n21566 9.3
R43043 vdd.n21583 vdd.n21582 9.3
R43044 vdd.n21599 vdd.n21598 9.3
R43045 vdd.n15340 vdd.n15339 9.3
R43046 vdd.n15339 vdd.n15338 9.3
R43047 vdd.n15326 vdd.n15325 9.3
R43048 vdd.n15325 vdd.n15324 9.3
R43049 vdd.n15305 vdd.n15304 9.3
R43050 vdd.n15304 vdd.n15303 9.3
R43051 vdd.n15289 vdd.n15288 9.3
R43052 vdd.n15288 vdd.n15287 9.3
R43053 vdd.n15275 vdd.n15274 9.3
R43054 vdd.n15274 vdd.n15273 9.3
R43055 vdd.n15264 vdd.n15263 9.3
R43056 vdd.n15263 vdd.n15262 9.3
R43057 vdd.n15412 vdd.n15411 9.3
R43058 vdd.n15411 vdd.n15410 9.3
R43059 vdd.n15397 vdd.n15396 9.3
R43060 vdd.n15396 vdd.n15395 9.3
R43061 vdd.n15383 vdd.n15382 9.3
R43062 vdd.n15382 vdd.n15381 9.3
R43063 vdd.n15369 vdd.n15368 9.3
R43064 vdd.n15368 vdd.n15367 9.3
R43065 vdd.n15355 vdd.n15354 9.3
R43066 vdd.n15354 vdd.n15353 9.3
R43067 vdd.n16538 vdd.n16537 9.3
R43068 vdd.n16537 vdd.n16536 9.3
R43069 vdd.n16521 vdd.n16520 9.3
R43070 vdd.n16520 vdd.n16519 9.3
R43071 vdd.n16504 vdd.n16503 9.3
R43072 vdd.n16503 vdd.n16502 9.3
R43073 vdd.n16487 vdd.n16486 9.3
R43074 vdd.n16486 vdd.n16485 9.3
R43075 vdd.n16467 vdd.n16466 9.3
R43076 vdd.n16466 vdd.n16465 9.3
R43077 vdd.n16450 vdd.n16449 9.3
R43078 vdd.n16449 vdd.n16448 9.3
R43079 vdd.n15134 vdd.n15133 9.3
R43080 vdd.n15133 vdd.n15132 9.3
R43081 vdd.n15148 vdd.n15147 9.3
R43082 vdd.n15147 vdd.n15146 9.3
R43083 vdd.n16430 vdd.n16429 9.3
R43084 vdd.n16429 vdd.n16428 9.3
R43085 vdd.n16413 vdd.n16412 9.3
R43086 vdd.n16412 vdd.n16411 9.3
R43087 vdd.n16396 vdd.n16395 9.3
R43088 vdd.n16395 vdd.n16394 9.3
R43089 vdd.n16379 vdd.n16378 9.3
R43090 vdd.n16378 vdd.n16377 9.3
R43091 vdd.n16362 vdd.n16361 9.3
R43092 vdd.n16361 vdd.n16360 9.3
R43093 vdd.n16345 vdd.n16344 9.3
R43094 vdd.n16344 vdd.n16343 9.3
R43095 vdd.n16328 vdd.n16327 9.3
R43096 vdd.n16327 vdd.n16326 9.3
R43097 vdd.n16301 vdd.n16300 9.3
R43098 vdd.n16300 vdd.n16299 9.3
R43099 vdd.n16282 vdd.n16281 9.3
R43100 vdd.n16281 vdd.n16280 9.3
R43101 vdd.n16265 vdd.n16264 9.3
R43102 vdd.n16264 vdd.n16263 9.3
R43103 vdd.n16248 vdd.n16247 9.3
R43104 vdd.n16247 vdd.n16246 9.3
R43105 vdd.n16231 vdd.n16230 9.3
R43106 vdd.n16230 vdd.n16229 9.3
R43107 vdd.n16211 vdd.n16210 9.3
R43108 vdd.n16210 vdd.n16209 9.3
R43109 vdd.n16194 vdd.n16193 9.3
R43110 vdd.n16193 vdd.n16192 9.3
R43111 vdd.n15162 vdd.n15161 9.3
R43112 vdd.n15161 vdd.n15160 9.3
R43113 vdd.n15176 vdd.n15175 9.3
R43114 vdd.n15175 vdd.n15174 9.3
R43115 vdd.n16174 vdd.n16173 9.3
R43116 vdd.n16173 vdd.n16172 9.3
R43117 vdd.n16157 vdd.n16156 9.3
R43118 vdd.n16156 vdd.n16155 9.3
R43119 vdd.n16140 vdd.n16139 9.3
R43120 vdd.n16139 vdd.n16138 9.3
R43121 vdd.n16123 vdd.n16122 9.3
R43122 vdd.n16122 vdd.n16121 9.3
R43123 vdd.n16106 vdd.n16105 9.3
R43124 vdd.n16105 vdd.n16104 9.3
R43125 vdd.n16089 vdd.n16088 9.3
R43126 vdd.n16088 vdd.n16087 9.3
R43127 vdd.n16072 vdd.n16071 9.3
R43128 vdd.n16071 vdd.n16070 9.3
R43129 vdd.n16045 vdd.n16044 9.3
R43130 vdd.n16044 vdd.n16043 9.3
R43131 vdd.n16026 vdd.n16025 9.3
R43132 vdd.n16025 vdd.n16024 9.3
R43133 vdd.n16009 vdd.n16008 9.3
R43134 vdd.n16008 vdd.n16007 9.3
R43135 vdd.n15992 vdd.n15991 9.3
R43136 vdd.n15991 vdd.n15990 9.3
R43137 vdd.n15975 vdd.n15974 9.3
R43138 vdd.n15974 vdd.n15973 9.3
R43139 vdd.n15955 vdd.n15954 9.3
R43140 vdd.n15954 vdd.n15953 9.3
R43141 vdd.n15938 vdd.n15937 9.3
R43142 vdd.n15937 vdd.n15936 9.3
R43143 vdd.n15193 vdd.n15192 9.3
R43144 vdd.n15194 vdd.n15193 9.3
R43145 vdd.n15204 vdd.n15203 9.3
R43146 vdd.n15203 vdd.n15202 9.3
R43147 vdd.n15918 vdd.n15917 9.3
R43148 vdd.n15917 vdd.n15916 9.3
R43149 vdd.n15901 vdd.n15900 9.3
R43150 vdd.n15900 vdd.n15899 9.3
R43151 vdd.n15884 vdd.n15883 9.3
R43152 vdd.n15883 vdd.n15882 9.3
R43153 vdd.n15867 vdd.n15866 9.3
R43154 vdd.n15866 vdd.n15865 9.3
R43155 vdd.n15850 vdd.n15849 9.3
R43156 vdd.n15849 vdd.n15848 9.3
R43157 vdd.n15833 vdd.n15832 9.3
R43158 vdd.n15832 vdd.n15831 9.3
R43159 vdd.n15816 vdd.n15815 9.3
R43160 vdd.n15815 vdd.n15814 9.3
R43161 vdd.n15789 vdd.n15788 9.3
R43162 vdd.n15788 vdd.n15787 9.3
R43163 vdd.n15770 vdd.n15769 9.3
R43164 vdd.n15769 vdd.n15768 9.3
R43165 vdd.n15753 vdd.n15752 9.3
R43166 vdd.n15752 vdd.n15751 9.3
R43167 vdd.n15736 vdd.n15735 9.3
R43168 vdd.n15735 vdd.n15734 9.3
R43169 vdd.n15719 vdd.n15718 9.3
R43170 vdd.n15718 vdd.n15717 9.3
R43171 vdd.n15699 vdd.n15698 9.3
R43172 vdd.n15698 vdd.n15697 9.3
R43173 vdd.n15682 vdd.n15681 9.3
R43174 vdd.n15681 vdd.n15680 9.3
R43175 vdd.n15218 vdd.n15217 9.3
R43176 vdd.n15217 vdd.n15216 9.3
R43177 vdd.n15232 vdd.n15231 9.3
R43178 vdd.n15231 vdd.n15230 9.3
R43179 vdd.n15662 vdd.n15661 9.3
R43180 vdd.n15661 vdd.n15660 9.3
R43181 vdd.n15645 vdd.n15644 9.3
R43182 vdd.n15644 vdd.n15643 9.3
R43183 vdd.n15628 vdd.n15627 9.3
R43184 vdd.n15627 vdd.n15626 9.3
R43185 vdd.n15611 vdd.n15610 9.3
R43186 vdd.n15610 vdd.n15609 9.3
R43187 vdd.n15594 vdd.n15593 9.3
R43188 vdd.n15593 vdd.n15592 9.3
R43189 vdd.n15577 vdd.n15576 9.3
R43190 vdd.n15576 vdd.n15575 9.3
R43191 vdd.n15560 vdd.n15559 9.3
R43192 vdd.n15559 vdd.n15558 9.3
R43193 vdd.n15533 vdd.n15532 9.3
R43194 vdd.n15532 vdd.n15531 9.3
R43195 vdd.n15514 vdd.n15513 9.3
R43196 vdd.n15513 vdd.n15512 9.3
R43197 vdd.n15497 vdd.n15496 9.3
R43198 vdd.n15496 vdd.n15495 9.3
R43199 vdd.n15480 vdd.n15479 9.3
R43200 vdd.n15479 vdd.n15478 9.3
R43201 vdd.n15463 vdd.n15462 9.3
R43202 vdd.n15462 vdd.n15461 9.3
R43203 vdd.n15443 vdd.n15442 9.3
R43204 vdd.n15442 vdd.n15441 9.3
R43205 vdd.n15429 vdd.n15428 9.3
R43206 vdd.n15428 vdd.n15427 9.3
R43207 vdd.n15243 vdd.n15242 9.3
R43208 vdd.n15242 vdd.n15241 9.3
R43209 vdd.n15254 vdd.n15253 9.3
R43210 vdd.n15253 vdd.n15252 9.3
R43211 vdd.n16552 vdd.n16551 9.3
R43212 vdd.n16616 vdd.n16615 9.3
R43213 vdd.n16624 vdd.n16623 9.3
R43214 vdd.n16632 vdd.n16631 9.3
R43215 vdd.n16644 vdd.n16643 9.3
R43216 vdd.n16665 vdd.n16664 9.3
R43217 vdd.n16656 vdd.n16655 9.3
R43218 vdd.n15079 vdd.n15078 9.3
R43219 vdd.n15118 vdd.n15117 9.3
R43220 vdd.n15117 vdd.n15116 9.3
R43221 vdd.n16558 vdd.n16557 9.3
R43222 vdd.n16574 vdd.n16573 9.3
R43223 vdd.n16573 vdd.n16572 9.3
R43224 vdd.n16572 vdd.n16571 9.3
R43225 vdd.n21703 vdd.n21702 9.3
R43226 vdd.n21704 vdd.n21703 9.3
R43227 vdd.n15015 vdd.n15014 9.3
R43228 vdd.n18399 vdd.n18398 9.3
R43229 vdd.n15025 vdd.n15024 9.3
R43230 vdd.n15024 vdd.n15023 9.3
R43231 vdd.n18367 vdd.n18366 9.3
R43232 vdd.n18366 vdd.n18365 9.3
R43233 vdd.n18346 vdd.n18345 9.3
R43234 vdd.n18345 vdd.n18344 9.3
R43235 vdd.n18329 vdd.n18328 9.3
R43236 vdd.n18328 vdd.n18327 9.3
R43237 vdd.n15036 vdd.n15035 9.3
R43238 vdd.n15035 vdd.n15034 9.3
R43239 vdd.n18304 vdd.n18303 9.3
R43240 vdd.n18303 vdd.n18302 9.3
R43241 vdd.n18289 vdd.n18288 9.3
R43242 vdd.n18288 vdd.n18287 9.3
R43243 vdd.n18274 vdd.n18273 9.3
R43244 vdd.n18273 vdd.n18272 9.3
R43245 vdd.n18259 vdd.n18258 9.3
R43246 vdd.n18258 vdd.n18257 9.3
R43247 vdd.n18244 vdd.n18243 9.3
R43248 vdd.n18243 vdd.n18242 9.3
R43249 vdd.n18229 vdd.n18228 9.3
R43250 vdd.n18228 vdd.n18227 9.3
R43251 vdd.n18214 vdd.n18213 9.3
R43252 vdd.n18213 vdd.n18212 9.3
R43253 vdd.n18198 vdd.n18197 9.3
R43254 vdd.n18197 vdd.n18196 9.3
R43255 vdd.n18178 vdd.n18177 9.3
R43256 vdd.n18177 vdd.n18176 9.3
R43257 vdd.n18162 vdd.n18161 9.3
R43258 vdd.n18161 vdd.n18160 9.3
R43259 vdd.n18146 vdd.n18145 9.3
R43260 vdd.n18145 vdd.n18144 9.3
R43261 vdd.n18130 vdd.n18129 9.3
R43262 vdd.n18129 vdd.n18128 9.3
R43263 vdd.n18114 vdd.n18113 9.3
R43264 vdd.n18113 vdd.n18112 9.3
R43265 vdd.n18098 vdd.n18097 9.3
R43266 vdd.n18097 vdd.n18096 9.3
R43267 vdd.n18082 vdd.n18081 9.3
R43268 vdd.n18081 vdd.n18080 9.3
R43269 vdd.n18066 vdd.n18065 9.3
R43270 vdd.n18065 vdd.n18064 9.3
R43271 vdd.n18038 vdd.n18037 9.3
R43272 vdd.n18037 vdd.n18036 9.3
R43273 vdd.n18022 vdd.n18021 9.3
R43274 vdd.n18021 vdd.n18020 9.3
R43275 vdd.n18006 vdd.n18005 9.3
R43276 vdd.n18005 vdd.n18004 9.3
R43277 vdd.n17990 vdd.n17989 9.3
R43278 vdd.n17989 vdd.n17988 9.3
R43279 vdd.n17974 vdd.n17973 9.3
R43280 vdd.n17973 vdd.n17972 9.3
R43281 vdd.n17958 vdd.n17957 9.3
R43282 vdd.n17957 vdd.n17956 9.3
R43283 vdd.n17942 vdd.n17941 9.3
R43284 vdd.n17941 vdd.n17940 9.3
R43285 vdd.n17926 vdd.n17925 9.3
R43286 vdd.n17925 vdd.n17924 9.3
R43287 vdd.n17906 vdd.n17905 9.3
R43288 vdd.n17905 vdd.n17904 9.3
R43289 vdd.n17890 vdd.n17889 9.3
R43290 vdd.n17889 vdd.n17888 9.3
R43291 vdd.n17874 vdd.n17873 9.3
R43292 vdd.n17873 vdd.t258 9.3
R43293 vdd.n17859 vdd.n17858 9.3
R43294 vdd.n17858 vdd.n17857 9.3
R43295 vdd.n17843 vdd.n17842 9.3
R43296 vdd.n17842 vdd.n17841 9.3
R43297 vdd.n17827 vdd.n17826 9.3
R43298 vdd.n17826 vdd.n17825 9.3
R43299 vdd.n17811 vdd.n17810 9.3
R43300 vdd.n17810 vdd.n17809 9.3
R43301 vdd.n17795 vdd.n17794 9.3
R43302 vdd.n17794 vdd.n17793 9.3
R43303 vdd.n17767 vdd.n17766 9.3
R43304 vdd.n17766 vdd.n17765 9.3
R43305 vdd.n17751 vdd.n17750 9.3
R43306 vdd.n17750 vdd.n17749 9.3
R43307 vdd.n17735 vdd.n17734 9.3
R43308 vdd.n17734 vdd.n17733 9.3
R43309 vdd.n17719 vdd.n17718 9.3
R43310 vdd.n17718 vdd.n17717 9.3
R43311 vdd.n17703 vdd.n17702 9.3
R43312 vdd.n17702 vdd.n17701 9.3
R43313 vdd.n17687 vdd.n17686 9.3
R43314 vdd.n17686 vdd.n17685 9.3
R43315 vdd.n17671 vdd.n17670 9.3
R43316 vdd.n17670 vdd.n17669 9.3
R43317 vdd.n17655 vdd.n17654 9.3
R43318 vdd.n17654 vdd.n17653 9.3
R43319 vdd.n17635 vdd.n17634 9.3
R43320 vdd.n17634 vdd.n17633 9.3
R43321 vdd.n17619 vdd.n17618 9.3
R43322 vdd.n17618 vdd.n17617 9.3
R43323 vdd.n17603 vdd.n17602 9.3
R43324 vdd.n17602 vdd.n17601 9.3
R43325 vdd.n17595 vdd.n17594 9.3
R43326 vdd.n17596 vdd.n17595 9.3
R43327 vdd.n17585 vdd.n17584 9.3
R43328 vdd.n17584 vdd.n17583 9.3
R43329 vdd.n17569 vdd.n17568 9.3
R43330 vdd.n17568 vdd.n17567 9.3
R43331 vdd.n17553 vdd.n17552 9.3
R43332 vdd.n17552 vdd.n17551 9.3
R43333 vdd.n17537 vdd.n17536 9.3
R43334 vdd.n17536 vdd.n17535 9.3
R43335 vdd.n17509 vdd.n17508 9.3
R43336 vdd.n17508 vdd.n17507 9.3
R43337 vdd.n17493 vdd.n17492 9.3
R43338 vdd.n17492 vdd.n17491 9.3
R43339 vdd.n17477 vdd.n17476 9.3
R43340 vdd.n17476 vdd.n17475 9.3
R43341 vdd.n17461 vdd.n17460 9.3
R43342 vdd.n17460 vdd.n17459 9.3
R43343 vdd.n17445 vdd.n17444 9.3
R43344 vdd.n17444 vdd.n17443 9.3
R43345 vdd.n17429 vdd.n17428 9.3
R43346 vdd.n17428 vdd.n17427 9.3
R43347 vdd.n17413 vdd.n17412 9.3
R43348 vdd.n17412 vdd.n17411 9.3
R43349 vdd.n17397 vdd.n17396 9.3
R43350 vdd.n17396 vdd.n17395 9.3
R43351 vdd.n17377 vdd.n17376 9.3
R43352 vdd.n17376 vdd.n17375 9.3
R43353 vdd.n17361 vdd.n17360 9.3
R43354 vdd.n17360 vdd.n17359 9.3
R43355 vdd.n17345 vdd.n17344 9.3
R43356 vdd.n17344 vdd.n17343 9.3
R43357 vdd.n17329 vdd.n17328 9.3
R43358 vdd.n17328 vdd.n17327 9.3
R43359 vdd.n17313 vdd.n17312 9.3
R43360 vdd.n17312 vdd.n17311 9.3
R43361 vdd.n17297 vdd.n17296 9.3
R43362 vdd.n17296 vdd.n17295 9.3
R43363 vdd.n17281 vdd.n17280 9.3
R43364 vdd.n17280 vdd.n17279 9.3
R43365 vdd.n17265 vdd.n17264 9.3
R43366 vdd.n17264 vdd.n17263 9.3
R43367 vdd.n17237 vdd.n17236 9.3
R43368 vdd.n17236 vdd.n17235 9.3
R43369 vdd.n17221 vdd.n17220 9.3
R43370 vdd.n17220 vdd.n17219 9.3
R43371 vdd.n17205 vdd.n17204 9.3
R43372 vdd.n17204 vdd.n17203 9.3
R43373 vdd.n17189 vdd.n17188 9.3
R43374 vdd.n17188 vdd.n17187 9.3
R43375 vdd.n17173 vdd.n17172 9.3
R43376 vdd.n17172 vdd.n17171 9.3
R43377 vdd.n17157 vdd.n17156 9.3
R43378 vdd.n17156 vdd.n17155 9.3
R43379 vdd.n17141 vdd.n17140 9.3
R43380 vdd.n17140 vdd.n17139 9.3
R43381 vdd.n17125 vdd.n17124 9.3
R43382 vdd.n17124 vdd.n17123 9.3
R43383 vdd.n17105 vdd.n17104 9.3
R43384 vdd.n17104 vdd.n17103 9.3
R43385 vdd.n17089 vdd.n17088 9.3
R43386 vdd.n17088 vdd.n17087 9.3
R43387 vdd.n17073 vdd.n17072 9.3
R43388 vdd.n17072 vdd.n17071 9.3
R43389 vdd.n17057 vdd.n17056 9.3
R43390 vdd.n17056 vdd.n17055 9.3
R43391 vdd.n17041 vdd.n17040 9.3
R43392 vdd.n17040 vdd.n17039 9.3
R43393 vdd.n17025 vdd.n17024 9.3
R43394 vdd.n17024 vdd.n17023 9.3
R43395 vdd.n17009 vdd.n17008 9.3
R43396 vdd.n17008 vdd.n17007 9.3
R43397 vdd.n16993 vdd.n16992 9.3
R43398 vdd.n16992 vdd.n16991 9.3
R43399 vdd.n16965 vdd.n16964 9.3
R43400 vdd.n16964 vdd.n16963 9.3
R43401 vdd.n16949 vdd.n16948 9.3
R43402 vdd.n16948 vdd.n16947 9.3
R43403 vdd.n16933 vdd.n16932 9.3
R43404 vdd.n16932 vdd.n16931 9.3
R43405 vdd.n16917 vdd.n16916 9.3
R43406 vdd.n16916 vdd.n16915 9.3
R43407 vdd.n16901 vdd.n16900 9.3
R43408 vdd.n16900 vdd.n16899 9.3
R43409 vdd.n16885 vdd.n16884 9.3
R43410 vdd.n16884 vdd.n16883 9.3
R43411 vdd.n16871 vdd.n16870 9.3
R43412 vdd.n16870 vdd.n16869 9.3
R43413 vdd.n18500 vdd.n18499 9.3
R43414 vdd.n18499 vdd.n18498 9.3
R43415 vdd.n18498 vdd.n18497 9.3
R43416 vdd.n18517 vdd.n18516 9.3
R43417 vdd.n18516 vdd.n18515 9.3
R43418 vdd.n18515 vdd.n18514 9.3
R43419 vdd.n18533 vdd.n18532 9.3
R43420 vdd.n18532 vdd.n18531 9.3
R43421 vdd.n18531 vdd.n18530 9.3
R43422 vdd.n18549 vdd.n18548 9.3
R43423 vdd.n18548 vdd.n18547 9.3
R43424 vdd.n18547 vdd.n18546 9.3
R43425 vdd.n18565 vdd.n18564 9.3
R43426 vdd.n18564 vdd.n18563 9.3
R43427 vdd.n18563 vdd.n18562 9.3
R43428 vdd.n18581 vdd.n18580 9.3
R43429 vdd.n18580 vdd.n18579 9.3
R43430 vdd.n18579 vdd.n18578 9.3
R43431 vdd.n18597 vdd.n18596 9.3
R43432 vdd.n18596 vdd.n18595 9.3
R43433 vdd.n18595 vdd.n18594 9.3
R43434 vdd.n18613 vdd.n18612 9.3
R43435 vdd.n18612 vdd.n18611 9.3
R43436 vdd.n18611 vdd.n18610 9.3
R43437 vdd.n18629 vdd.n18628 9.3
R43438 vdd.n18628 vdd.n18627 9.3
R43439 vdd.n18627 vdd.n18626 9.3
R43440 vdd.n18647 vdd.n18646 9.3
R43441 vdd.n18646 vdd.n18645 9.3
R43442 vdd.n18645 vdd.n18644 9.3
R43443 vdd.n18663 vdd.n18662 9.3
R43444 vdd.n18662 vdd.n18661 9.3
R43445 vdd.n18661 vdd.n18660 9.3
R43446 vdd.n18679 vdd.n18678 9.3
R43447 vdd.n18678 vdd.n18677 9.3
R43448 vdd.n18677 vdd.n18676 9.3
R43449 vdd.n18695 vdd.n18694 9.3
R43450 vdd.n18694 vdd.n18693 9.3
R43451 vdd.n18693 vdd.n18692 9.3
R43452 vdd.n18711 vdd.n18710 9.3
R43453 vdd.n18710 vdd.n18709 9.3
R43454 vdd.n18709 vdd.n18708 9.3
R43455 vdd.n18727 vdd.n18726 9.3
R43456 vdd.n18726 vdd.n18725 9.3
R43457 vdd.n18725 vdd.n18724 9.3
R43458 vdd.n18743 vdd.n18742 9.3
R43459 vdd.n18742 vdd.n18741 9.3
R43460 vdd.n18741 vdd.n18740 9.3
R43461 vdd.n18759 vdd.n18758 9.3
R43462 vdd.n18758 vdd.n18757 9.3
R43463 vdd.n18757 vdd.n18756 9.3
R43464 vdd.n18776 vdd.n18775 9.3
R43465 vdd.n18775 vdd.n18774 9.3
R43466 vdd.n18774 vdd.n18773 9.3
R43467 vdd.n18792 vdd.n18791 9.3
R43468 vdd.n18791 vdd.n18790 9.3
R43469 vdd.n18790 vdd.n18789 9.3
R43470 vdd.n18808 vdd.n18807 9.3
R43471 vdd.n18807 vdd.n18806 9.3
R43472 vdd.n18806 vdd.n18805 9.3
R43473 vdd.n18824 vdd.n18823 9.3
R43474 vdd.n18823 vdd.n18822 9.3
R43475 vdd.n18822 vdd.n18821 9.3
R43476 vdd.n18840 vdd.n18839 9.3
R43477 vdd.n18839 vdd.n18838 9.3
R43478 vdd.n18838 vdd.n18837 9.3
R43479 vdd.n18856 vdd.n18855 9.3
R43480 vdd.n18855 vdd.n18854 9.3
R43481 vdd.n18854 vdd.n18853 9.3
R43482 vdd.n18872 vdd.n18871 9.3
R43483 vdd.n18871 vdd.n18870 9.3
R43484 vdd.n18870 vdd.n18869 9.3
R43485 vdd.n18888 vdd.n18887 9.3
R43486 vdd.n18887 vdd.n18886 9.3
R43487 vdd.n18886 vdd.n18885 9.3
R43488 vdd.n18906 vdd.n18905 9.3
R43489 vdd.n18905 vdd.n18904 9.3
R43490 vdd.n18904 vdd.n18903 9.3
R43491 vdd.n18922 vdd.n18921 9.3
R43492 vdd.n18921 vdd.n18920 9.3
R43493 vdd.n18920 vdd.n18919 9.3
R43494 vdd.n18938 vdd.n18937 9.3
R43495 vdd.n18937 vdd.n18936 9.3
R43496 vdd.n18936 vdd.n18935 9.3
R43497 vdd.n18954 vdd.n18953 9.3
R43498 vdd.n18953 vdd.n18952 9.3
R43499 vdd.n18952 vdd.n18951 9.3
R43500 vdd.n18970 vdd.n18969 9.3
R43501 vdd.n18969 vdd.n18968 9.3
R43502 vdd.n18968 vdd.n18967 9.3
R43503 vdd.n18986 vdd.n18985 9.3
R43504 vdd.n18985 vdd.n18984 9.3
R43505 vdd.n18984 vdd.n18983 9.3
R43506 vdd.n19002 vdd.n19001 9.3
R43507 vdd.n19001 vdd.n19000 9.3
R43508 vdd.n19000 vdd.n18999 9.3
R43509 vdd.n19018 vdd.n19017 9.3
R43510 vdd.n19017 vdd.n19016 9.3
R43511 vdd.n19016 vdd.n19015 9.3
R43512 vdd.n19035 vdd.n19034 9.3
R43513 vdd.n19034 vdd.n19033 9.3
R43514 vdd.n19033 vdd.n19032 9.3
R43515 vdd.n19051 vdd.n19050 9.3
R43516 vdd.n19050 vdd.n19049 9.3
R43517 vdd.n19049 vdd.n19048 9.3
R43518 vdd.n19067 vdd.n19066 9.3
R43519 vdd.n19066 vdd.n19065 9.3
R43520 vdd.n19065 vdd.n19064 9.3
R43521 vdd.n19083 vdd.n19082 9.3
R43522 vdd.n19082 vdd.n19081 9.3
R43523 vdd.n19081 vdd.n19080 9.3
R43524 vdd.n19099 vdd.n19098 9.3
R43525 vdd.n19098 vdd.n19097 9.3
R43526 vdd.n19097 vdd.n19096 9.3
R43527 vdd.n19115 vdd.n19114 9.3
R43528 vdd.n19114 vdd.n19113 9.3
R43529 vdd.n19113 vdd.n19112 9.3
R43530 vdd.n19130 vdd.n19129 9.3
R43531 vdd.n19129 vdd.n19128 9.3
R43532 vdd.n19128 vdd.n19127 9.3
R43533 vdd.n19140 vdd.n19139 9.3
R43534 vdd.n19139 vdd.n19138 9.3
R43535 vdd.n21015 vdd.n21014 9.3
R43536 vdd.n19147 vdd.n19146 9.3
R43537 vdd.n21029 vdd.n21028 9.3
R43538 vdd.n21028 vdd.n21027 9.3
R43539 vdd.n21027 vdd.n21026 9.3
R43540 vdd.n21045 vdd.n21044 9.3
R43541 vdd.n21044 vdd.n21043 9.3
R43542 vdd.n21043 vdd.n21042 9.3
R43543 vdd.n21061 vdd.n21060 9.3
R43544 vdd.n21060 vdd.n21059 9.3
R43545 vdd.n21059 vdd.n21058 9.3
R43546 vdd.n21077 vdd.n21076 9.3
R43547 vdd.n21076 vdd.n21075 9.3
R43548 vdd.n21075 vdd.n21074 9.3
R43549 vdd.n21088 vdd.n21087 9.3
R43550 vdd.n21087 vdd.n21086 9.3
R43551 vdd.n21109 vdd.n21108 9.3
R43552 vdd.n21108 vdd.n21107 9.3
R43553 vdd.n21107 vdd.n21106 9.3
R43554 vdd.n21125 vdd.n21124 9.3
R43555 vdd.n21124 vdd.n21123 9.3
R43556 vdd.n21123 vdd.n21122 9.3
R43557 vdd.n21142 vdd.n21141 9.3
R43558 vdd.n21141 vdd.n21140 9.3
R43559 vdd.n21140 vdd.n21139 9.3
R43560 vdd.n21158 vdd.n21157 9.3
R43561 vdd.n21157 vdd.n21156 9.3
R43562 vdd.n21156 vdd.n21155 9.3
R43563 vdd.n21174 vdd.n21173 9.3
R43564 vdd.n21173 vdd.n21172 9.3
R43565 vdd.n21172 vdd.n21171 9.3
R43566 vdd.n21190 vdd.n21189 9.3
R43567 vdd.n21189 vdd.n21188 9.3
R43568 vdd.n21188 vdd.n21187 9.3
R43569 vdd.n21206 vdd.n21205 9.3
R43570 vdd.n21205 vdd.n21204 9.3
R43571 vdd.n21204 vdd.n21203 9.3
R43572 vdd.n21222 vdd.n21221 9.3
R43573 vdd.n21221 vdd.n21220 9.3
R43574 vdd.n21220 vdd.n21219 9.3
R43575 vdd.n21238 vdd.n21237 9.3
R43576 vdd.n21237 vdd.n21236 9.3
R43577 vdd.n21236 vdd.n21235 9.3
R43578 vdd.n21254 vdd.n21253 9.3
R43579 vdd.n21253 vdd.n21252 9.3
R43580 vdd.n21252 vdd.n21251 9.3
R43581 vdd.n21272 vdd.n21271 9.3
R43582 vdd.n21271 vdd.n21270 9.3
R43583 vdd.n21270 vdd.n21269 9.3
R43584 vdd.n21288 vdd.n21287 9.3
R43585 vdd.n21287 vdd.n21286 9.3
R43586 vdd.n21286 vdd.n21285 9.3
R43587 vdd.n21304 vdd.n21303 9.3
R43588 vdd.n21303 vdd.n21302 9.3
R43589 vdd.n21302 vdd.n21301 9.3
R43590 vdd.n21320 vdd.n21319 9.3
R43591 vdd.n21319 vdd.n21318 9.3
R43592 vdd.n21318 vdd.n21317 9.3
R43593 vdd.n21336 vdd.n21335 9.3
R43594 vdd.n21335 vdd.n21334 9.3
R43595 vdd.n21334 vdd.n21333 9.3
R43596 vdd.n21352 vdd.n21351 9.3
R43597 vdd.n21351 vdd.n21350 9.3
R43598 vdd.n21350 vdd.n21349 9.3
R43599 vdd.n21368 vdd.n21367 9.3
R43600 vdd.n21367 vdd.n21366 9.3
R43601 vdd.n21366 vdd.n21365 9.3
R43602 vdd.n21384 vdd.n21383 9.3
R43603 vdd.n21383 vdd.n21382 9.3
R43604 vdd.n21382 vdd.n21381 9.3
R43605 vdd.n21401 vdd.n21400 9.3
R43606 vdd.n21400 vdd.n21399 9.3
R43607 vdd.n21399 vdd.n21398 9.3
R43608 vdd.n21417 vdd.n21416 9.3
R43609 vdd.n21416 vdd.n21415 9.3
R43610 vdd.n21415 vdd.n21414 9.3
R43611 vdd.n21433 vdd.n21432 9.3
R43612 vdd.n21432 vdd.n21431 9.3
R43613 vdd.n21431 vdd.n21430 9.3
R43614 vdd.n21449 vdd.n21448 9.3
R43615 vdd.n21448 vdd.n21447 9.3
R43616 vdd.n21447 vdd.n21446 9.3
R43617 vdd.n21465 vdd.n21464 9.3
R43618 vdd.n21464 vdd.n21463 9.3
R43619 vdd.n21463 vdd.n21462 9.3
R43620 vdd.n21481 vdd.n21480 9.3
R43621 vdd.n21480 vdd.n21479 9.3
R43622 vdd.n21479 vdd.n21478 9.3
R43623 vdd.n21497 vdd.n21496 9.3
R43624 vdd.n21496 vdd.n21495 9.3
R43625 vdd.n21495 vdd.n21494 9.3
R43626 vdd.n21513 vdd.n21512 9.3
R43627 vdd.n21512 vdd.n21511 9.3
R43628 vdd.n21511 vdd.n21510 9.3
R43629 vdd.n21531 vdd.n21530 9.3
R43630 vdd.n21530 vdd.n21529 9.3
R43631 vdd.n21529 vdd.n21528 9.3
R43632 vdd.n21547 vdd.n21546 9.3
R43633 vdd.n21546 vdd.n21545 9.3
R43634 vdd.n21545 vdd.n21544 9.3
R43635 vdd.n21563 vdd.n21562 9.3
R43636 vdd.n21562 vdd.n21561 9.3
R43637 vdd.n21561 vdd.n21560 9.3
R43638 vdd.n21579 vdd.n21578 9.3
R43639 vdd.n21578 vdd.n21577 9.3
R43640 vdd.n21577 vdd.n21576 9.3
R43641 vdd.n21595 vdd.n21594 9.3
R43642 vdd.n21594 vdd.n21593 9.3
R43643 vdd.n21593 vdd.n21592 9.3
R43644 vdd.n21619 vdd.n21618 9.3
R43645 vdd.n21618 vdd.n21617 9.3
R43646 vdd.n21617 vdd.n21616 9.3
R43647 vdd.n21607 vdd.n21606 9.3
R43648 vdd.n21664 vdd.n21663 9.3
R43649 vdd.n21676 vdd.n21675 9.3
R43650 vdd.n21675 vdd.n21674 9.3
R43651 vdd.n21674 vdd.n21673 9.3
R43652 vdd.n20067 vdd.n20066 9.3
R43653 vdd.n20083 vdd.n20082 9.3
R43654 vdd.n20099 vdd.n20098 9.3
R43655 vdd.n20115 vdd.n20114 9.3
R43656 vdd.n20131 vdd.n20130 9.3
R43657 vdd.n20175 vdd.n20174 9.3
R43658 vdd.n20191 vdd.n20190 9.3
R43659 vdd.n20207 vdd.n20206 9.3
R43660 vdd.n20223 vdd.n20222 9.3
R43661 vdd.n20239 vdd.n20238 9.3
R43662 vdd.n20255 vdd.n20254 9.3
R43663 vdd.n20287 vdd.n20286 9.3
R43664 vdd.n20303 vdd.n20302 9.3
R43665 vdd.n20319 vdd.n20318 9.3
R43666 vdd.n20335 vdd.n20334 9.3
R43667 vdd.n20351 vdd.n20350 9.3
R43668 vdd.n20367 vdd.n20366 9.3
R43669 vdd.n20411 vdd.n20410 9.3
R43670 vdd.n20427 vdd.n20426 9.3
R43671 vdd.n20443 vdd.n20442 9.3
R43672 vdd.n20458 vdd.n20457 9.3
R43673 vdd.n20468 vdd.n20467 9.3
R43674 vdd.n20469 vdd.n20468 9.3
R43675 vdd.n20470 vdd.n20469 9.3
R43676 vdd.n20464 vdd.n20463 9.3
R43677 vdd.n20463 vdd.n20462 9.3
R43678 vdd.n20456 vdd.n20455 9.3
R43679 vdd.n20454 vdd.n20453 9.3
R43680 vdd.n20453 vdd.n20452 9.3
R43681 vdd.n20452 vdd.n20451 9.3
R43682 vdd.n20441 vdd.n20440 9.3
R43683 vdd.n20439 vdd.n20438 9.3
R43684 vdd.n20438 vdd.n20437 9.3
R43685 vdd.n20437 vdd.n20436 9.3
R43686 vdd.n20425 vdd.n20424 9.3
R43687 vdd.n20423 vdd.n20422 9.3
R43688 vdd.n20422 vdd.n20421 9.3
R43689 vdd.n20421 vdd.n20420 9.3
R43690 vdd.n20409 vdd.n20408 9.3
R43691 vdd.n20407 vdd.n20406 9.3
R43692 vdd.n20406 vdd.n20405 9.3
R43693 vdd.n20405 vdd.n20404 9.3
R43694 vdd.n20384 vdd.n20383 9.3
R43695 vdd.n20383 vdd.n20382 9.3
R43696 vdd.n20382 vdd.n20381 9.3
R43697 vdd.n20369 vdd.n20368 9.3
R43698 vdd.n20365 vdd.n20364 9.3
R43699 vdd.n20364 vdd.n20363 9.3
R43700 vdd.n20363 vdd.n20362 9.3
R43701 vdd.n20353 vdd.n20352 9.3
R43702 vdd.n20349 vdd.n20348 9.3
R43703 vdd.n20348 vdd.n20347 9.3
R43704 vdd.n20347 vdd.n20346 9.3
R43705 vdd.n20337 vdd.n20336 9.3
R43706 vdd.n20333 vdd.n20332 9.3
R43707 vdd.n20332 vdd.n20331 9.3
R43708 vdd.n20331 vdd.n20330 9.3
R43709 vdd.n20321 vdd.n20320 9.3
R43710 vdd.n20317 vdd.n20316 9.3
R43711 vdd.n20316 vdd.n20315 9.3
R43712 vdd.n20315 vdd.n20314 9.3
R43713 vdd.n20305 vdd.n20304 9.3
R43714 vdd.n20301 vdd.n20300 9.3
R43715 vdd.n20300 vdd.n20299 9.3
R43716 vdd.n20299 vdd.n20298 9.3
R43717 vdd.n20289 vdd.n20288 9.3
R43718 vdd.n20285 vdd.n20284 9.3
R43719 vdd.n20284 vdd.n20283 9.3
R43720 vdd.n20283 vdd.n20282 9.3
R43721 vdd.n20273 vdd.n20272 9.3
R43722 vdd.n20000 vdd.n19999 9.3
R43723 vdd.n19999 vdd.n19998 9.3
R43724 vdd.n20012 vdd.n20011 9.3
R43725 vdd.n20011 vdd.n20010 9.3
R43726 vdd.n20269 vdd.n20268 9.3
R43727 vdd.n20267 vdd.n20266 9.3
R43728 vdd.n20266 vdd.n20265 9.3
R43729 vdd.n20265 vdd.n20264 9.3
R43730 vdd.n20253 vdd.n20252 9.3
R43731 vdd.n20251 vdd.n20250 9.3
R43732 vdd.n20250 vdd.n20249 9.3
R43733 vdd.n20249 vdd.n20248 9.3
R43734 vdd.n20237 vdd.n20236 9.3
R43735 vdd.n20235 vdd.n20234 9.3
R43736 vdd.n20234 vdd.n20233 9.3
R43737 vdd.n20233 vdd.n20232 9.3
R43738 vdd.n20221 vdd.n20220 9.3
R43739 vdd.n20219 vdd.n20218 9.3
R43740 vdd.n20218 vdd.n20217 9.3
R43741 vdd.n20217 vdd.n20216 9.3
R43742 vdd.n20205 vdd.n20204 9.3
R43743 vdd.n20203 vdd.n20202 9.3
R43744 vdd.n20202 vdd.n20201 9.3
R43745 vdd.n20201 vdd.n20200 9.3
R43746 vdd.n20189 vdd.n20188 9.3
R43747 vdd.n20187 vdd.n20186 9.3
R43748 vdd.n20186 vdd.n20185 9.3
R43749 vdd.n20185 vdd.n20184 9.3
R43750 vdd.n20173 vdd.n20172 9.3
R43751 vdd.n20171 vdd.n20170 9.3
R43752 vdd.n20170 vdd.n20169 9.3
R43753 vdd.n20169 vdd.n20168 9.3
R43754 vdd.n20148 vdd.n20147 9.3
R43755 vdd.n20147 vdd.n20146 9.3
R43756 vdd.n20146 vdd.n20145 9.3
R43757 vdd.n20133 vdd.n20132 9.3
R43758 vdd.n20129 vdd.n20128 9.3
R43759 vdd.n20128 vdd.n20127 9.3
R43760 vdd.n20127 vdd.n20126 9.3
R43761 vdd.n20117 vdd.n20116 9.3
R43762 vdd.n20113 vdd.n20112 9.3
R43763 vdd.n20112 vdd.n20111 9.3
R43764 vdd.n20111 vdd.n20110 9.3
R43765 vdd.n20101 vdd.n20100 9.3
R43766 vdd.n20097 vdd.n20096 9.3
R43767 vdd.n20096 vdd.n20095 9.3
R43768 vdd.n20095 vdd.n20094 9.3
R43769 vdd.n20085 vdd.n20084 9.3
R43770 vdd.n20081 vdd.n20080 9.3
R43771 vdd.n20080 vdd.n20079 9.3
R43772 vdd.n20079 vdd.n20078 9.3
R43773 vdd.n20069 vdd.n20068 9.3
R43774 vdd.n20065 vdd.n20064 9.3
R43775 vdd.n20064 vdd.n20063 9.3
R43776 vdd.n20063 vdd.n20062 9.3
R43777 vdd.n20549 vdd.n20548 9.3
R43778 vdd.n20565 vdd.n20564 9.3
R43779 vdd.n20581 vdd.n20580 9.3
R43780 vdd.n20597 vdd.n20596 9.3
R43781 vdd.n20613 vdd.n20612 9.3
R43782 vdd.n20648 vdd.n20647 9.3
R43783 vdd.n20664 vdd.n20663 9.3
R43784 vdd.n20680 vdd.n20679 9.3
R43785 vdd.n20692 vdd.n20691 9.3
R43786 vdd.n20691 vdd.n20690 9.3
R43787 vdd.n20690 vdd.n20689 9.3
R43788 vdd.n20678 vdd.n20677 9.3
R43789 vdd.n20676 vdd.n20675 9.3
R43790 vdd.n20675 vdd.n20674 9.3
R43791 vdd.n20674 vdd.n20673 9.3
R43792 vdd.n20662 vdd.n20661 9.3
R43793 vdd.n20660 vdd.n20659 9.3
R43794 vdd.n20659 vdd.n20658 9.3
R43795 vdd.n20658 vdd.n20657 9.3
R43796 vdd.n20646 vdd.n20645 9.3
R43797 vdd.n20644 vdd.n20643 9.3
R43798 vdd.n20643 vdd.n20642 9.3
R43799 vdd.n20642 vdd.n20641 9.3
R43800 vdd.n20627 vdd.n20626 9.3
R43801 vdd.n20626 vdd.n20625 9.3
R43802 vdd.n20625 vdd.n20624 9.3
R43803 vdd.n20615 vdd.n20614 9.3
R43804 vdd.n20611 vdd.n20610 9.3
R43805 vdd.n20610 vdd.n20609 9.3
R43806 vdd.n20609 vdd.n20608 9.3
R43807 vdd.n20599 vdd.n20598 9.3
R43808 vdd.n20595 vdd.n20594 9.3
R43809 vdd.n20594 vdd.n20593 9.3
R43810 vdd.n20593 vdd.n20592 9.3
R43811 vdd.n20583 vdd.n20582 9.3
R43812 vdd.n20579 vdd.n20578 9.3
R43813 vdd.n20578 vdd.n20577 9.3
R43814 vdd.n20577 vdd.n20576 9.3
R43815 vdd.n20567 vdd.n20566 9.3
R43816 vdd.n20563 vdd.n20562 9.3
R43817 vdd.n20562 vdd.n20561 9.3
R43818 vdd.n20561 vdd.n20560 9.3
R43819 vdd.n20551 vdd.n20550 9.3
R43820 vdd.n20547 vdd.n20546 9.3
R43821 vdd.n20546 vdd.n20545 9.3
R43822 vdd.n20545 vdd.n20544 9.3
R43823 vdd.n20696 vdd.n20695 9.3
R43824 vdd.n20711 vdd.n20710 9.3
R43825 vdd.n20755 vdd.n20754 9.3
R43826 vdd.n20770 vdd.n19900 9.3
R43827 vdd.n20786 vdd.n20785 9.3
R43828 vdd.n20802 vdd.n20801 9.3
R43829 vdd.n20863 vdd.n20862 9.3
R43830 vdd.n20868 vdd.n20867 9.3
R43831 vdd.n20884 vdd.n20883 9.3
R43832 vdd.n20900 vdd.n20899 9.3
R43833 vdd.n20945 vdd.n20944 9.3
R43834 vdd.n20961 vdd.n20960 9.3
R43835 vdd.n20977 vdd.n20976 9.3
R43836 vdd.n20993 vdd.n20992 9.3
R43837 vdd.n19796 vdd.n19795 9.3
R43838 vdd.n19780 vdd.n19779 9.3
R43839 vdd.n19764 vdd.n19763 9.3
R43840 vdd.n19748 vdd.n19747 9.3
R43841 vdd.n19703 vdd.n19702 9.3
R43842 vdd.n19687 vdd.n19686 9.3
R43843 vdd.n19671 vdd.n19670 9.3
R43844 vdd.n19655 vdd.n19654 9.3
R43845 vdd.n19594 vdd.n19593 9.3
R43846 vdd.n19578 vdd.n19577 9.3
R43847 vdd.n19562 vdd.n19561 9.3
R43848 vdd.n19546 vdd.n19545 9.3
R43849 vdd.n19502 vdd.n19501 9.3
R43850 vdd.n19487 vdd.n19486 9.3
R43851 vdd.n19485 vdd.n19484 9.3
R43852 vdd.n19499 vdd.n19498 9.3
R43853 vdd.n19498 vdd.n19497 9.3
R43854 vdd.n19497 vdd.n19496 9.3
R43855 vdd.n19500 vdd.n19284 9.3
R43856 vdd.n19514 vdd.n19513 9.3
R43857 vdd.n19513 vdd.n19512 9.3
R43858 vdd.n19512 vdd.n19511 9.3
R43859 vdd.n19516 vdd.n19515 9.3
R43860 vdd.n19281 vdd.n19280 9.3
R43861 vdd.n19280 vdd.n19279 9.3
R43862 vdd.n19519 vdd.n19518 9.3
R43863 vdd.n19269 vdd.n19268 9.3
R43864 vdd.n19268 vdd.n19267 9.3
R43865 vdd.n19257 vdd.n19256 9.3
R43866 vdd.n19256 vdd.n19255 9.3
R43867 vdd.n19529 vdd.n19528 9.3
R43868 vdd.n19245 vdd.n19244 9.3
R43869 vdd.n19244 vdd.n19243 9.3
R43870 vdd.n19532 vdd.n19531 9.3
R43871 vdd.n19544 vdd.n19543 9.3
R43872 vdd.n19543 vdd.n19542 9.3
R43873 vdd.n19542 vdd.n19541 9.3
R43874 vdd.n19548 vdd.n19547 9.3
R43875 vdd.n19560 vdd.n19559 9.3
R43876 vdd.n19559 vdd.n19558 9.3
R43877 vdd.n19558 vdd.n19557 9.3
R43878 vdd.n19564 vdd.n19563 9.3
R43879 vdd.n19576 vdd.n19575 9.3
R43880 vdd.n19575 vdd.n19574 9.3
R43881 vdd.n19574 vdd.n19573 9.3
R43882 vdd.n19580 vdd.n19579 9.3
R43883 vdd.n19592 vdd.n19591 9.3
R43884 vdd.n19591 vdd.n19590 9.3
R43885 vdd.n19590 vdd.n19589 9.3
R43886 vdd.n19596 vdd.n19595 9.3
R43887 vdd.n19608 vdd.n19607 9.3
R43888 vdd.n19607 vdd.n19606 9.3
R43889 vdd.n19606 vdd.n19605 9.3
R43890 vdd.n19624 vdd.n19623 9.3
R43891 vdd.n19623 vdd.n19622 9.3
R43892 vdd.n19622 vdd.n19621 9.3
R43893 vdd.n19638 vdd.n19637 9.3
R43894 vdd.n19637 vdd.n19636 9.3
R43895 vdd.n19636 vdd.n19635 9.3
R43896 vdd.n19651 vdd.n19650 9.3
R43897 vdd.n19650 vdd.n19649 9.3
R43898 vdd.n19649 vdd.n19648 9.3
R43899 vdd.n19653 vdd.n19652 9.3
R43900 vdd.n19667 vdd.n19666 9.3
R43901 vdd.n19666 vdd.n19665 9.3
R43902 vdd.n19665 vdd.n19664 9.3
R43903 vdd.n19669 vdd.n19668 9.3
R43904 vdd.n19683 vdd.n19682 9.3
R43905 vdd.n19682 vdd.n19681 9.3
R43906 vdd.n19681 vdd.n19680 9.3
R43907 vdd.n19685 vdd.n19684 9.3
R43908 vdd.n19699 vdd.n19698 9.3
R43909 vdd.n19698 vdd.n19697 9.3
R43910 vdd.n19697 vdd.n19696 9.3
R43911 vdd.n19701 vdd.n19700 9.3
R43912 vdd.n19715 vdd.n19714 9.3
R43913 vdd.n19714 vdd.n19713 9.3
R43914 vdd.n19713 vdd.n19712 9.3
R43915 vdd.n19717 vdd.n19716 9.3
R43916 vdd.n19225 vdd.n19224 9.3
R43917 vdd.n19224 vdd.n19223 9.3
R43918 vdd.n19720 vdd.n19719 9.3
R43919 vdd.n19213 vdd.n19212 9.3
R43920 vdd.n19212 vdd.n19211 9.3
R43921 vdd.n19201 vdd.n19200 9.3
R43922 vdd.n19200 vdd.n19199 9.3
R43923 vdd.n19730 vdd.n19729 9.3
R43924 vdd.n19188 vdd.n19187 9.3
R43925 vdd.n19187 vdd.n19186 9.3
R43926 vdd.n19734 vdd.n19733 9.3
R43927 vdd.n19746 vdd.n19745 9.3
R43928 vdd.n19745 vdd.n19744 9.3
R43929 vdd.n19744 vdd.n19743 9.3
R43930 vdd.n19750 vdd.n19749 9.3
R43931 vdd.n19762 vdd.n19761 9.3
R43932 vdd.n19761 vdd.n19760 9.3
R43933 vdd.n19760 vdd.n19759 9.3
R43934 vdd.n19766 vdd.n19765 9.3
R43935 vdd.n19778 vdd.n19777 9.3
R43936 vdd.n19777 vdd.n19776 9.3
R43937 vdd.n19776 vdd.n19775 9.3
R43938 vdd.n19782 vdd.n19781 9.3
R43939 vdd.n19794 vdd.n19793 9.3
R43940 vdd.n19793 vdd.n19792 9.3
R43941 vdd.n19792 vdd.n19791 9.3
R43942 vdd.n19798 vdd.n19797 9.3
R43943 vdd.n19810 vdd.n19809 9.3
R43944 vdd.n19809 vdd.n19808 9.3
R43945 vdd.n19808 vdd.n19807 9.3
R43946 vdd.n19826 vdd.n19825 9.3
R43947 vdd.n19825 vdd.n19824 9.3
R43948 vdd.n19824 vdd.n19823 9.3
R43949 vdd.n19172 vdd.n19171 9.3
R43950 vdd.n19171 vdd.n19170 9.3
R43951 vdd.n20997 vdd.n20996 9.3
R43952 vdd.n20998 vdd.n20997 9.3
R43953 vdd.n20999 vdd.n20998 9.3
R43954 vdd.n20995 vdd.n20994 9.3
R43955 vdd.n20991 vdd.n20990 9.3
R43956 vdd.n20990 vdd.n20989 9.3
R43957 vdd.n20989 vdd.n20988 9.3
R43958 vdd.n20979 vdd.n20978 9.3
R43959 vdd.n20975 vdd.n20974 9.3
R43960 vdd.n20974 vdd.n20973 9.3
R43961 vdd.n20973 vdd.n20972 9.3
R43962 vdd.n20963 vdd.n20962 9.3
R43963 vdd.n20959 vdd.n20958 9.3
R43964 vdd.n20958 vdd.n20957 9.3
R43965 vdd.n20957 vdd.n20956 9.3
R43966 vdd.n20947 vdd.n20946 9.3
R43967 vdd.n20943 vdd.n20942 9.3
R43968 vdd.n20942 vdd.n20941 9.3
R43969 vdd.n20941 vdd.n20940 9.3
R43970 vdd.n20931 vdd.n20930 9.3
R43971 vdd.n19842 vdd.n19841 9.3
R43972 vdd.n19841 vdd.n19840 9.3
R43973 vdd.n20927 vdd.n20926 9.3
R43974 vdd.n19855 vdd.n19854 9.3
R43975 vdd.n19854 vdd.n19853 9.3
R43976 vdd.n19867 vdd.n19866 9.3
R43977 vdd.n19866 vdd.n19865 9.3
R43978 vdd.n20917 vdd.n20916 9.3
R43979 vdd.n19879 vdd.n19878 9.3
R43980 vdd.n19878 vdd.n19877 9.3
R43981 vdd.n20914 vdd.n20913 9.3
R43982 vdd.n20912 vdd.n20911 9.3
R43983 vdd.n20911 vdd.n20910 9.3
R43984 vdd.n20910 vdd.n20909 9.3
R43985 vdd.n20898 vdd.n20897 9.3
R43986 vdd.n20896 vdd.n20895 9.3
R43987 vdd.n20895 vdd.n20894 9.3
R43988 vdd.n20894 vdd.n20893 9.3
R43989 vdd.n20882 vdd.n20881 9.3
R43990 vdd.n20880 vdd.n20879 9.3
R43991 vdd.n20879 vdd.n20878 9.3
R43992 vdd.n20878 vdd.n20877 9.3
R43993 vdd.n20866 vdd.n20865 9.3
R43994 vdd.n20864 vdd.n19892 9.3
R43995 vdd.n19892 vdd.n19891 9.3
R43996 vdd.n19891 vdd.n19890 9.3
R43997 vdd.n20861 vdd.n20860 9.3
R43998 vdd.n20859 vdd.n20858 9.3
R43999 vdd.n20858 vdd.n20857 9.3
R44000 vdd.n20857 vdd.n20856 9.3
R44001 vdd.n20846 vdd.n20845 9.3
R44002 vdd.n20845 vdd.n20844 9.3
R44003 vdd.n20844 vdd.n20843 9.3
R44004 vdd.n20829 vdd.n20828 9.3
R44005 vdd.n20828 vdd.n20827 9.3
R44006 vdd.n20827 vdd.n20826 9.3
R44007 vdd.n20816 vdd.n20815 9.3
R44008 vdd.n20815 vdd.n20814 9.3
R44009 vdd.n20814 vdd.n20813 9.3
R44010 vdd.n20804 vdd.n20803 9.3
R44011 vdd.n20800 vdd.n20799 9.3
R44012 vdd.n20799 vdd.n20798 9.3
R44013 vdd.n20798 vdd.n20797 9.3
R44014 vdd.n20788 vdd.n20787 9.3
R44015 vdd.n20784 vdd.n20783 9.3
R44016 vdd.n20783 vdd.n20782 9.3
R44017 vdd.n20782 vdd.n20781 9.3
R44018 vdd.n20772 vdd.n20771 9.3
R44019 vdd.n20769 vdd.n20768 9.3
R44020 vdd.n20768 vdd.n20767 9.3
R44021 vdd.n20767 vdd.n20766 9.3
R44022 vdd.n20757 vdd.n20756 9.3
R44023 vdd.n20753 vdd.n20752 9.3
R44024 vdd.n20752 vdd.n20751 9.3
R44025 vdd.n20751 vdd.n20750 9.3
R44026 vdd.n20741 vdd.n20740 9.3
R44027 vdd.n19911 vdd.n19910 9.3
R44028 vdd.n19910 vdd.n19909 9.3
R44029 vdd.n20738 vdd.n20737 9.3
R44030 vdd.n19923 vdd.n19922 9.3
R44031 vdd.n19922 vdd.n19921 9.3
R44032 vdd.n19935 vdd.n19934 9.3
R44033 vdd.n19934 vdd.n19933 9.3
R44034 vdd.n20728 vdd.n20727 9.3
R44035 vdd.n19947 vdd.n19946 9.3
R44036 vdd.n19946 vdd.n19945 9.3
R44037 vdd.n20725 vdd.n20724 9.3
R44038 vdd.n20723 vdd.n20722 9.3
R44039 vdd.n20722 vdd.n20721 9.3
R44040 vdd.n20721 vdd.n20720 9.3
R44041 vdd.n20709 vdd.n19950 9.3
R44042 vdd.n20708 vdd.n20707 9.3
R44043 vdd.n20707 vdd.n20706 9.3
R44044 vdd.n20706 vdd.n20705 9.3
R44045 vdd.n20694 vdd.n20693 9.3
R44046 vdd.n19471 vdd.n19470 9.3
R44047 vdd.n19455 vdd.n19454 9.3
R44048 vdd.n19439 vdd.n19438 9.3
R44049 vdd.n19404 vdd.n19403 9.3
R44050 vdd.n19388 vdd.n19387 9.3
R44051 vdd.n19372 vdd.n19371 9.3
R44052 vdd.n19356 vdd.n19355 9.3
R44053 vdd.n19340 vdd.n19339 9.3
R44054 vdd.n19338 vdd.n19337 9.3
R44055 vdd.n19337 vdd.n19336 9.3
R44056 vdd.n19336 vdd.n19335 9.3
R44057 vdd.n19342 vdd.n19341 9.3
R44058 vdd.n19354 vdd.n19353 9.3
R44059 vdd.n19353 vdd.n19352 9.3
R44060 vdd.n19352 vdd.n19351 9.3
R44061 vdd.n19358 vdd.n19357 9.3
R44062 vdd.n19370 vdd.n19369 9.3
R44063 vdd.n19369 vdd.n19368 9.3
R44064 vdd.n19368 vdd.n19367 9.3
R44065 vdd.n19374 vdd.n19373 9.3
R44066 vdd.n19386 vdd.n19385 9.3
R44067 vdd.n19385 vdd.n19384 9.3
R44068 vdd.n19384 vdd.n19383 9.3
R44069 vdd.n19390 vdd.n19389 9.3
R44070 vdd.n19402 vdd.n19401 9.3
R44071 vdd.n19401 vdd.n19400 9.3
R44072 vdd.n19400 vdd.n19399 9.3
R44073 vdd.n19406 vdd.n19405 9.3
R44074 vdd.n19421 vdd.n19420 9.3
R44075 vdd.n19420 vdd.n19419 9.3
R44076 vdd.n19419 vdd.n19418 9.3
R44077 vdd.n19435 vdd.n19434 9.3
R44078 vdd.n19434 vdd.n19433 9.3
R44079 vdd.n19433 vdd.n19432 9.3
R44080 vdd.n19437 vdd.n19436 9.3
R44081 vdd.n19451 vdd.n19450 9.3
R44082 vdd.n19450 vdd.n19449 9.3
R44083 vdd.n19449 vdd.n19448 9.3
R44084 vdd.n19453 vdd.n19452 9.3
R44085 vdd.n19467 vdd.n19466 9.3
R44086 vdd.n19466 vdd.n19465 9.3
R44087 vdd.n19465 vdd.n19464 9.3
R44088 vdd.n19469 vdd.n19468 9.3
R44089 vdd.n19483 vdd.n19482 9.3
R44090 vdd.n19482 vdd.n19481 9.3
R44091 vdd.n19481 vdd.n19480 9.3
R44092 vdd.n21812 vdd.n21811 9.3
R44093 vdd.n21810 vdd.n21809 9.3
R44094 vdd.n21820 vdd.n21819 9.3
R44095 vdd.n21819 vdd.n21818 9.3
R44096 vdd.n21776 vdd.n21775 9.3
R44097 vdd.n21783 vdd.n21782 9.3
R44098 vdd.n21793 vdd.n21792 9.3
R44099 vdd.n21766 vdd.n21765 9.3
R44100 vdd.n21796 vdd.n21795 9.3
R44101 vdd.n21791 vdd.n21790 9.3
R44102 vdd.n21785 vdd.n21784 9.3
R44103 vdd.n21781 vdd.n21780 9.3
R44104 vdd.n21778 vdd.n21777 9.3
R44105 vdd.n21774 vdd.n21773 9.3
R44106 vdd.n21919 vdd.n21906 9.3
R44107 vdd.n21913 vdd.n21906 9.3
R44108 vdd.n21922 vdd.n21905 9.3
R44109 vdd.n21921 vdd.n21920 9.3
R44110 vdd.n21918 vdd.n21908 9.3
R44111 vdd.n21918 vdd.n21917 9.3
R44112 vdd.n21911 vdd.n21907 9.3
R44113 vdd.n21938 vdd.n21933 9.3
R44114 vdd.n21943 vdd.n21942 9.3
R44115 vdd.n21951 vdd.n21901 9.3
R44116 vdd.n21954 vdd.n21953 9.3
R44117 vdd.n21957 vdd.n21956 9.3
R44118 vdd.n21944 vdd.n21930 9.3
R44119 vdd.n21941 vdd.n21932 9.3
R44120 vdd.n21940 vdd.n21939 9.3
R44121 vdd.n21937 vdd.n21936 9.3
R44122 vdd.n21948 vdd.n21929 9.3
R44123 vdd.n21950 vdd.n21949 9.3
R44124 vdd.n21743 vdd.n21742 9.3
R44125 vdd.n21742 vdd.n21741 9.3
R44126 vdd.n24524 vdd.n24520 9.3
R44127 vdd.n24553 vdd.n24552 9.3
R44128 vdd.n24972 vdd.n24971 9.3
R44129 vdd.n24906 vdd.n24905 9.3
R44130 vdd.n24896 vdd.n24895 9.3
R44131 vdd.n25008 vdd.n25007 9.3
R44132 vdd.n25022 vdd.n25021 9.3
R44133 vdd.n25032 vdd.n25031 9.3
R44134 vdd.n25046 vdd.n25045 9.3
R44135 vdd.n25044 vdd.n25043 9.3
R44136 vdd.n25042 vdd.n25041 9.3
R44137 vdd.n25039 vdd.n25038 9.3
R44138 vdd.n25035 vdd.n25034 9.3
R44139 vdd.n25037 vdd.n25036 9.3
R44140 vdd.n25030 vdd.n25029 9.3
R44141 vdd.n25028 vdd.n25027 9.3
R44142 vdd.n25019 vdd.n25018 9.3
R44143 vdd.n25017 vdd.n25016 9.3
R44144 vdd.n25015 vdd.n25014 9.3
R44145 vdd.n25010 vdd.n25009 9.3
R44146 vdd.n25012 vdd.n25011 9.3
R44147 vdd.n25005 vdd.n25004 9.3
R44148 vdd.n25003 vdd.n25002 9.3
R44149 vdd.n25001 vdd.n25000 9.3
R44150 vdd.n24996 vdd.n24995 9.3
R44151 vdd.n24998 vdd.n24997 9.3
R44152 vdd.n25050 vdd.n25049 9.3
R44153 vdd.n24915 vdd.n24914 9.3
R44154 vdd.n24574 vdd.n24573 9.3
R44155 vdd.n24581 vdd.n24580 9.3
R44156 vdd.n24588 vdd.n24587 9.3
R44157 vdd.n24595 vdd.n24594 9.3
R44158 vdd.n24605 vdd.n24604 9.3
R44159 vdd.n24612 vdd.n24611 9.3
R44160 vdd.n24619 vdd.n24618 9.3
R44161 vdd.n24617 vdd.n24616 9.3
R44162 vdd.n24614 vdd.n24613 9.3
R44163 vdd.n24610 vdd.n24609 9.3
R44164 vdd.n24607 vdd.n24606 9.3
R44165 vdd.n24603 vdd.n24602 9.3
R44166 vdd.n24597 vdd.n24596 9.3
R44167 vdd.n24593 vdd.n24592 9.3
R44168 vdd.n24591 vdd.n24590 9.3
R44169 vdd.n24586 vdd.n24585 9.3
R44170 vdd.n24584 vdd.n24583 9.3
R44171 vdd.n24579 vdd.n24578 9.3
R44172 vdd.n24577 vdd.n24576 9.3
R44173 vdd.n24572 vdd.n24571 9.3
R44174 vdd.n24624 vdd.n24623 9.3
R44175 vdd.n24629 vdd.n24628 9.3
R44176 vdd.n24631 vdd.n24630 9.3
R44177 vdd.n24681 vdd.n24680 9.3
R44178 vdd.n24680 vdd.n24679 9.3
R44179 vdd.n25139 vdd.n25138 9.3
R44180 vdd.n24683 vdd.n24682 9.3
R44181 vdd.n24685 vdd.n24684 9.3
R44182 vdd.n24693 vdd.n24692 9.3
R44183 vdd.n24692 vdd.n24691 9.3
R44184 vdd.n24695 vdd.n24694 9.3
R44185 vdd.n24697 vdd.n24696 9.3
R44186 vdd.n24705 vdd.n24704 9.3
R44187 vdd.n24704 vdd.n24703 9.3
R44188 vdd.n24707 vdd.n24706 9.3
R44189 vdd.n24709 vdd.n24708 9.3
R44190 vdd.n24717 vdd.n24716 9.3
R44191 vdd.n24716 vdd.n24715 9.3
R44192 vdd.n24514 vdd.n24513 9.3
R44193 vdd.n24983 vdd.n24982 9.3
R44194 vdd.n25148 vdd.n25147 9.3
R44195 vdd.n25147 vdd.n25146 9.3
R44196 vdd.n25150 vdd.n25149 9.3
R44197 vdd.n25152 vdd.n25151 9.3
R44198 vdd.n25160 vdd.n25159 9.3
R44199 vdd.n25159 vdd.n25158 9.3
R44200 vdd.n25176 vdd.n25175 9.3
R44201 vdd.n25175 vdd.n25174 9.3
R44202 vdd.n25178 vdd.n25177 9.3
R44203 vdd.n25180 vdd.n25179 9.3
R44204 vdd.n25188 vdd.n25187 9.3
R44205 vdd.n25187 vdd.n25186 9.3
R44206 vdd.n25190 vdd.n25189 9.3
R44207 vdd.n25192 vdd.n25191 9.3
R44208 vdd.n25200 vdd.n25199 9.3
R44209 vdd.n25199 vdd.n25198 9.3
R44210 vdd.n25202 vdd.n25201 9.3
R44211 vdd.n25204 vdd.n25203 9.3
R44212 vdd.n25212 vdd.n25211 9.3
R44213 vdd.n25211 vdd.n25210 9.3
R44214 vdd.n25214 vdd.n25213 9.3
R44215 vdd.n25216 vdd.n25215 9.3
R44216 vdd.n25224 vdd.n25223 9.3
R44217 vdd.n25223 vdd.n25222 9.3
R44218 vdd.n25226 vdd.n25225 9.3
R44219 vdd.n25228 vdd.n25227 9.3
R44220 vdd.n25236 vdd.n25235 9.3
R44221 vdd.n25235 vdd.n25234 9.3
R44222 vdd.n25238 vdd.n25237 9.3
R44223 vdd.n25240 vdd.n25239 9.3
R44224 vdd.n25248 vdd.n25247 9.3
R44225 vdd.n25247 vdd.n25246 9.3
R44226 vdd.n25250 vdd.n25249 9.3
R44227 vdd.n24832 vdd.n24831 9.3
R44228 vdd.n24830 vdd.n24829 9.3
R44229 vdd.n24829 vdd.n24828 9.3
R44230 vdd.n24822 vdd.n24821 9.3
R44231 vdd.n24820 vdd.n24819 9.3
R44232 vdd.n24818 vdd.n24817 9.3
R44233 vdd.n24817 vdd.n24816 9.3
R44234 vdd.n24810 vdd.n24809 9.3
R44235 vdd.n24808 vdd.n24807 9.3
R44236 vdd.n24806 vdd.n24805 9.3
R44237 vdd.n24805 vdd.n24804 9.3
R44238 vdd.n24798 vdd.n24797 9.3
R44239 vdd.n24796 vdd.n24795 9.3
R44240 vdd.n24794 vdd.n24793 9.3
R44241 vdd.n24793 vdd.n24792 9.3
R44242 vdd.n24786 vdd.n24785 9.3
R44243 vdd.n24784 vdd.n24783 9.3
R44244 vdd.n24782 vdd.n24781 9.3
R44245 vdd.n24781 vdd.n24780 9.3
R44246 vdd.n24774 vdd.n24773 9.3
R44247 vdd.n24772 vdd.n24771 9.3
R44248 vdd.n24770 vdd.n24769 9.3
R44249 vdd.n24769 vdd.n24768 9.3
R44250 vdd.n24762 vdd.n24761 9.3
R44251 vdd.n24760 vdd.n24759 9.3
R44252 vdd.n24758 vdd.n24757 9.3
R44253 vdd.n24757 vdd.n24756 9.3
R44254 vdd.n24744 vdd.n24743 9.3
R44255 vdd.n24743 vdd.n24742 9.3
R44256 vdd.n24734 vdd.n24733 9.3
R44257 vdd.n24732 vdd.n24731 9.3
R44258 vdd.n24730 vdd.n24729 9.3
R44259 vdd.n24729 vdd.n24728 9.3
R44260 vdd.n24721 vdd.n24720 9.3
R44261 vdd.n24719 vdd.n24718 9.3
R44262 vdd.n25137 vdd.n25136 9.3
R44263 vdd.n25135 vdd.n25134 9.3
R44264 vdd.n25134 vdd.n25133 9.3
R44265 vdd.n25127 vdd.n25126 9.3
R44266 vdd.n25125 vdd.n25124 9.3
R44267 vdd.n25123 vdd.n25122 9.3
R44268 vdd.n25122 vdd.n25121 9.3
R44269 vdd.n25115 vdd.n25114 9.3
R44270 vdd.n25113 vdd.n25112 9.3
R44271 vdd.n25111 vdd.n25110 9.3
R44272 vdd.n25110 vdd.n25109 9.3
R44273 vdd.n25103 vdd.n25102 9.3
R44274 vdd.n25101 vdd.n25100 9.3
R44275 vdd.n25099 vdd.n25098 9.3
R44276 vdd.n25098 vdd.n25097 9.3
R44277 vdd.t319 vdd.n9263 9.276
R44278 vdd.n13336 vdd.t284 9.175
R44279 vdd.n21543 vdd.n21540 9.148
R44280 vdd.n21493 vdd.n21490 9.148
R44281 vdd.n21284 vdd.n21281 9.148
R44282 vdd.n21234 vdd.n21231 9.148
R44283 vdd.n18918 vdd.n18915 9.148
R44284 vdd.n18868 vdd.n18865 9.148
R44285 vdd.n18659 vdd.n18656 9.148
R44286 vdd.n18609 vdd.n18606 9.148
R44287 vdd.n27655 vdd.n27651 9.114
R44288 vdd.n26077 vdd.n26073 9.114
R44289 vdd.n11865 vdd.n11837 9.02
R44290 vdd.n21956 vdd.n21928 9.02
R44291 vdd.n11715 vdd.n11690 9.019
R44292 vdd.n21765 vdd.n21764 9.019
R44293 vdd.n11715 vdd.n11691 9.019
R44294 vdd.n11846 vdd.n11837 9.019
R44295 vdd.n21937 vdd.n21928 9.019
R44296 vdd.n9442 vdd.n9441 8.986
R44297 vdd.n9609 vdd.n9608 8.986
R44298 vdd.n9801 vdd.n9800 8.986
R44299 vdd.n9969 vdd.n9968 8.986
R44300 vdd.n10244 vdd.n10243 8.986
R44301 vdd.n11184 vdd.t383 8.986
R44302 vdd.n27655 vdd.n27644 8.908
R44303 vdd.n26077 vdd.n26065 8.908
R44304 vdd.n24815 vdd.n24814 8.907
R44305 vdd.n25096 vdd.n25095 8.907
R44306 vdd.n27655 vdd.n27649 8.897
R44307 vdd.n26077 vdd.n26071 8.897
R44308 vdd.n11883 vdd.n11882 8.889
R44309 vdd.n21974 vdd.n21973 8.889
R44310 vdd.n27655 vdd.n27647 8.885
R44311 vdd.n26077 vdd.n26069 8.885
R44312 vdd.n10100 vdd.n10072 8.876
R44313 vdd.t102 vdd.n8317 8.869
R44314 vdd.n14547 vdd.t322 8.869
R44315 vdd.n33707 vdd.n33705 8.868
R44316 vdd.n33480 vdd.n33478 8.868
R44317 vdd.n34080 vdd.n34078 8.868
R44318 vdd.n33869 vdd.n33868 8.868
R44319 vdd.n34349 vdd.n34347 8.868
R44320 vdd.n35120 vdd.n35119 8.868
R44321 vdd.n35367 vdd.n35365 8.868
R44322 vdd.n35239 vdd.n35237 8.868
R44323 vdd.n34652 vdd.n34650 8.868
R44324 vdd.n34533 vdd.n34532 8.868
R44325 vdd.n34777 vdd.n34775 8.868
R44326 vdd.n791 vdd.n789 8.868
R44327 vdd.n965 vdd.n963 8.868
R44328 vdd.n224 vdd.n222 8.868
R44329 vdd.n3 vdd.n1 8.868
R44330 vdd.n6143 vdd.n6142 8.868
R44331 vdd.n6055 vdd.n6053 8.868
R44332 vdd.n5782 vdd.n5780 8.868
R44333 vdd.n5399 vdd.n5397 8.868
R44334 vdd.n5280 vdd.n5279 8.868
R44335 vdd.n5524 vdd.n5522 8.868
R44336 vdd.n4793 vdd.n4792 8.868
R44337 vdd.n4955 vdd.n4953 8.868
R44338 vdd.n4804 vdd.n4802 8.868
R44339 vdd.n4229 vdd.n4227 8.868
R44340 vdd.n4110 vdd.n4109 8.868
R44341 vdd.n4351 vdd.n4349 8.868
R44342 vdd.n27300 vdd.n27298 8.868
R44343 vdd.n27277 vdd.n27275 8.868
R44344 vdd.n27587 vdd.n27586 8.868
R44345 vdd.n25752 vdd.n25750 8.868
R44346 vdd.n25723 vdd.n25721 8.868
R44347 vdd.n26003 vdd.n26002 8.868
R44348 vdd.n25445 vdd.n25443 8.868
R44349 vdd.n24634 vdd.n24633 8.864
R44350 vdd.n36036 vdd.n36035 8.855
R44351 vdd.n36035 vdd.n36034 8.855
R44352 vdd.n36267 vdd.n36266 8.855
R44353 vdd.n36266 vdd.n36265 8.855
R44354 vdd.n36498 vdd.n36497 8.855
R44355 vdd.n36497 vdd.n36496 8.855
R44356 vdd.n36729 vdd.n36728 8.855
R44357 vdd.n36728 vdd.n36727 8.855
R44358 vdd.n36960 vdd.n36959 8.855
R44359 vdd.n36959 vdd.n36958 8.855
R44360 vdd.n37156 vdd.n37155 8.855
R44361 vdd.n37155 vdd.n37154 8.855
R44362 vdd.n35653 vdd.n35652 8.855
R44363 vdd.n35652 vdd.n35651 8.855
R44364 vdd.n37549 vdd.n37548 8.855
R44365 vdd.n37548 vdd.n37547 8.855
R44366 vdd.n38015 vdd.n38014 8.855
R44367 vdd.n38014 vdd.n38013 8.855
R44368 vdd.n37784 vdd.n37783 8.855
R44369 vdd.n37783 vdd.n37782 8.855
R44370 vdd.n28226 vdd.n28225 8.855
R44371 vdd.n28225 vdd.n28224 8.855
R44372 vdd.n28457 vdd.n28456 8.855
R44373 vdd.n28456 vdd.n28455 8.855
R44374 vdd.n28688 vdd.n28687 8.855
R44375 vdd.n28687 vdd.n28686 8.855
R44376 vdd.n28891 vdd.n28890 8.855
R44377 vdd.n28890 vdd.n28889 8.855
R44378 vdd.n32028 vdd.n32027 8.855
R44379 vdd.n30689 vdd.n30688 8.855
R44380 vdd.n30688 vdd.n30687 8.855
R44381 vdd.n2890 vdd.n2889 8.855
R44382 vdd.n3071 vdd.n3070 8.855
R44383 vdd.n3252 vdd.n3251 8.855
R44384 vdd.n3433 vdd.n3432 8.855
R44385 vdd.n3614 vdd.n3613 8.855
R44386 vdd.n3807 vdd.n3806 8.855
R44387 vdd.n2510 vdd.n2509 8.855
R44388 vdd.n1835 vdd.n1834 8.855
R44389 vdd.n1652 vdd.n1651 8.855
R44390 vdd.n1471 vdd.n1470 8.855
R44391 vdd.n1290 vdd.n1289 8.855
R44392 vdd.n26937 vdd.n26936 8.855
R44393 vdd.n27118 vdd.n27117 8.855
R44394 vdd.n26667 vdd.n26666 8.855
R44395 vdd.n32030 vdd.n32029 8.855
R44396 vdd.n32029 vdd.n32028 8.855
R44397 vdd.n32387 vdd.n32386 8.855
R44398 vdd.n14418 vdd.n14417 8.855
R44399 vdd.n14419 vdd.n14418 8.855
R44400 vdd.n14152 vdd.n14151 8.855
R44401 vdd.n14153 vdd.n14152 8.855
R44402 vdd.n13863 vdd.n13862 8.855
R44403 vdd.n13864 vdd.n13863 8.855
R44404 vdd.n13534 vdd.n8960 8.855
R44405 vdd.n8960 vdd.n8944 8.855
R44406 vdd.n13242 vdd.n9181 8.855
R44407 vdd.n9181 vdd.n9165 8.855
R44408 vdd.n13374 vdd.n13373 8.855
R44409 vdd.n13375 vdd.n13374 8.855
R44410 vdd.n13666 vdd.n13665 8.855
R44411 vdd.n13667 vdd.n13666 8.855
R44412 vdd.n13963 vdd.n13962 8.855
R44413 vdd.n13962 vdd.n13961 8.855
R44414 vdd.n14253 vdd.n14252 8.855
R44415 vdd.n14252 vdd.n14251 8.855
R44416 vdd.n18634 vdd.n18633 8.855
R44417 vdd.n18633 vdd.n18632 8.855
R44418 vdd.n18893 vdd.n18892 8.855
R44419 vdd.n18892 vdd.n18891 8.855
R44420 vdd.n21011 vdd.n21010 8.855
R44421 vdd.n21010 vdd.n21009 8.855
R44422 vdd.n21259 vdd.n21258 8.855
R44423 vdd.n21258 vdd.n21257 8.855
R44424 vdd.n21518 vdd.n21517 8.855
R44425 vdd.n21517 vdd.n21516 8.855
R44426 vdd.n19525 vdd.n19524 8.855
R44427 vdd.n19524 vdd.n19523 8.855
R44428 vdd.n19726 vdd.n19725 8.855
R44429 vdd.n19725 vdd.n19724 8.855
R44430 vdd.n20923 vdd.n20922 8.855
R44431 vdd.n20922 vdd.n20921 8.855
R44432 vdd.n20734 vdd.n20733 8.855
R44433 vdd.n20733 vdd.n20732 8.855
R44434 vdd.n25396 vdd.n25388 8.854
R44435 vdd.n25396 vdd.n25384 8.843
R44436 vdd.n11715 vdd.n11692 8.838
R44437 vdd.n11716 vdd.n11715 8.838
R44438 vdd.n11861 vdd.n11837 8.838
R44439 vdd.n11843 vdd.n11837 8.838
R44440 vdd.n21952 vdd.n21928 8.838
R44441 vdd.n21934 vdd.n21928 8.838
R44442 vdd.n953 vdd.n952 8.833
R44443 vdd.n25396 vdd.n25395 8.833
R44444 vdd.n27655 vdd.n27654 8.832
R44445 vdd.n26077 vdd.n26076 8.832
R44446 vdd.n25396 vdd.n25393 8.832
R44447 vdd.n10246 vdd.n10236 8.8
R44448 vdd.n16669 vdd.n16668 8.8
R44449 vdd.n19266 vdd.n19263 8.796
R44450 vdd.n19254 vdd.n19251 8.796
R44451 vdd.n19210 vdd.n19207 8.796
R44452 vdd.n19198 vdd.n19195 8.796
R44453 vdd.n19743 vdd.t144 8.796
R44454 vdd.n20940 vdd.t162 8.796
R44455 vdd.n19852 vdd.n19849 8.796
R44456 vdd.n19864 vdd.n19861 8.796
R44457 vdd.n19920 vdd.n19917 8.796
R44458 vdd.n19932 vdd.n19929 8.796
R44459 vdd.n20404 vdd.n20400 8.796
R44460 vdd.n20381 vdd.n20380 8.796
R44461 vdd.n20168 vdd.n20164 8.796
R44462 vdd.n20145 vdd.n20144 8.796
R44463 vdd.n14684 vdd.n8119 8.774
R44464 vdd.n14713 vdd.n14712 8.774
R44465 vdd.n14858 vdd.n8030 8.774
R44466 vdd.n14906 vdd.n8020 8.774
R44467 vdd.n11598 vdd.n11597 8.77
R44468 vdd.n24512 vdd.n24509 8.767
R44469 vdd.n10246 vdd.n10230 8.693
R44470 vdd.n16669 vdd.n16645 8.693
R44471 vdd.n9343 vdd.n9342 8.665
R44472 vdd.n9518 vdd.n9508 8.665
R44473 vdd.n9703 vdd.n9702 8.665
R44474 vdd.n9878 vdd.n9868 8.665
R44475 vdd.n10157 vdd.n10156 8.665
R44476 vdd.n15531 vdd.n15530 8.665
R44477 vdd.n15787 vdd.n15786 8.665
R44478 vdd.n16043 vdd.n16042 8.665
R44479 vdd.n16299 vdd.n16298 8.665
R44480 vdd.n16571 vdd.n16570 8.665
R44481 vdd.n13377 vdd.t335 8.564
R44482 vdd.n30285 vdd.n30284 8.537
R44483 vdd.n10491 vdd.n10490 8.533
R44484 vdd.n12585 vdd.n10122 8.533
R44485 vdd.n12599 vdd.n10097 8.533
R44486 vdd.n12602 vdd.n12601 8.533
R44487 vdd.n10137 vdd.n10090 8.533
R44488 vdd.n10285 vdd.n10281 8.533
R44489 vdd.n10458 vdd.n10457 8.533
R44490 vdd.n10294 vdd.n10292 8.533
R44491 vdd.n10445 vdd.n10295 8.533
R44492 vdd.n10438 vdd.n10437 8.533
R44493 vdd.n10427 vdd.n10426 8.533
R44494 vdd.n10421 vdd.n10311 8.533
R44495 vdd.n10413 vdd.n10412 8.533
R44496 vdd.n10328 vdd.n10324 8.533
R44497 vdd.n10398 vdd.n10333 8.533
R44498 vdd.n10347 vdd.n10338 8.533
R44499 vdd.n10384 vdd.n10383 8.533
R44500 vdd.n10375 vdd.n10351 8.533
R44501 vdd.n10360 vdd.n10358 8.533
R44502 vdd.n13078 vdd.n9293 8.533
R44503 vdd.n9303 vdd.n9300 8.533
R44504 vdd.n13064 vdd.n13063 8.533
R44505 vdd.n9312 vdd.n9310 8.533
R44506 vdd.n9337 vdd.n9336 8.533
R44507 vdd.n9348 vdd.n9347 8.533
R44508 vdd.n13040 vdd.n13039 8.533
R44509 vdd.n9373 vdd.n9352 8.533
R44510 vdd.n9381 vdd.n9380 8.533
R44511 vdd.n9390 vdd.n9389 8.533
R44512 vdd.n13018 vdd.n9394 8.533
R44513 vdd.n13010 vdd.n13009 8.533
R44514 vdd.n9427 vdd.n9405 8.533
R44515 vdd.n9445 vdd.n9444 8.533
R44516 vdd.n12991 vdd.n9418 8.533
R44517 vdd.n9449 vdd.n9423 8.533
R44518 vdd.n12977 vdd.n12976 8.533
R44519 vdd.n9459 vdd.n9457 8.533
R44520 vdd.n9488 vdd.n9487 8.533
R44521 vdd.n9490 vdd.n9481 8.533
R44522 vdd.n12953 vdd.n9478 8.533
R44523 vdd.n9513 vdd.n9510 8.533
R44524 vdd.n12939 vdd.n12938 8.533
R44525 vdd.n9532 vdd.n9531 8.533
R44526 vdd.n9545 vdd.n9544 8.533
R44527 vdd.n12923 vdd.n9549 8.533
R44528 vdd.n12915 vdd.n12914 8.533
R44529 vdd.n9584 vdd.n9560 8.533
R44530 vdd.n9591 vdd.n9590 8.533
R44531 vdd.n9600 vdd.n9599 8.533
R44532 vdd.n12893 vdd.n9604 8.533
R44533 vdd.n12885 vdd.n12884 8.533
R44534 vdd.n9638 vdd.n9637 8.533
R44535 vdd.n9640 vdd.n9628 8.533
R44536 vdd.n12870 vdd.n9625 8.533
R44537 vdd.n9663 vdd.n9660 8.533
R44538 vdd.n12856 vdd.n12855 8.533
R44539 vdd.n9673 vdd.n9671 8.533
R44540 vdd.n9697 vdd.n9696 8.533
R44541 vdd.n9708 vdd.n9707 8.533
R44542 vdd.n12832 vdd.n12831 8.533
R44543 vdd.n9733 vdd.n9712 8.533
R44544 vdd.n9741 vdd.n9740 8.533
R44545 vdd.n9750 vdd.n9749 8.533
R44546 vdd.n12810 vdd.n9754 8.533
R44547 vdd.n12802 vdd.n12801 8.533
R44548 vdd.n9787 vdd.n9765 8.533
R44549 vdd.n9804 vdd.n9803 8.533
R44550 vdd.n12783 vdd.n9779 8.533
R44551 vdd.n9808 vdd.n9783 8.533
R44552 vdd.n12769 vdd.n12768 8.533
R44553 vdd.n9819 vdd.n9817 8.533
R44554 vdd.n9848 vdd.n9847 8.533
R44555 vdd.n9850 vdd.n9841 8.533
R44556 vdd.n12745 vdd.n9838 8.533
R44557 vdd.n9873 vdd.n9870 8.533
R44558 vdd.n12731 vdd.n12730 8.533
R44559 vdd.n9893 vdd.n9892 8.533
R44560 vdd.n9905 vdd.n9904 8.533
R44561 vdd.n12715 vdd.n9909 8.533
R44562 vdd.n12707 vdd.n12706 8.533
R44563 vdd.n9944 vdd.n9919 8.533
R44564 vdd.n9951 vdd.n9950 8.533
R44565 vdd.n9960 vdd.n9959 8.533
R44566 vdd.n12685 vdd.n9964 8.533
R44567 vdd.n12677 vdd.n12676 8.533
R44568 vdd.n9998 vdd.n9997 8.533
R44569 vdd.n10000 vdd.n9988 8.533
R44570 vdd.n12662 vdd.n9985 8.533
R44571 vdd.n10023 vdd.n10020 8.533
R44572 vdd.n12648 vdd.n12647 8.533
R44573 vdd.n10033 vdd.n10031 8.533
R44574 vdd.n10151 vdd.n10150 8.533
R44575 vdd.n10186 vdd.n10086 8.533
R44576 vdd.n12523 vdd.n10521 8.533
R44577 vdd.n10546 vdd.n10545 8.533
R44578 vdd.n10557 vdd.n10556 8.533
R44579 vdd.n12510 vdd.n12509 8.533
R44580 vdd.n12499 vdd.n12498 8.533
R44581 vdd.n12493 vdd.n10568 8.533
R44582 vdd.n10594 vdd.n10593 8.533
R44583 vdd.n10591 vdd.n10587 8.533
R44584 vdd.n12475 vdd.n12474 8.533
R44585 vdd.n10609 vdd.n10607 8.533
R44586 vdd.n10636 vdd.n10635 8.533
R44587 vdd.n10643 vdd.n10642 8.533
R44588 vdd.n10651 vdd.n10626 8.533
R44589 vdd.n12446 vdd.n12445 8.533
R44590 vdd.n10660 vdd.n10658 8.533
R44591 vdd.n10693 vdd.n10692 8.533
R44592 vdd.n12422 vdd.n12421 8.533
R44593 vdd.n12411 vdd.n12410 8.533
R44594 vdd.n12405 vdd.n10703 8.533
R44595 vdd.n10731 vdd.n10730 8.533
R44596 vdd.n10742 vdd.n10741 8.533
R44597 vdd.n12391 vdd.n12390 8.533
R44598 vdd.n12380 vdd.n12379 8.533
R44599 vdd.n10760 vdd.n10759 8.533
R44600 vdd.n10787 vdd.n10786 8.533
R44601 vdd.n10794 vdd.n10793 8.533
R44602 vdd.n10802 vdd.n10777 8.533
R44603 vdd.n12357 vdd.n12356 8.533
R44604 vdd.n10811 vdd.n10809 8.533
R44605 vdd.n10835 vdd.n10834 8.533
R44606 vdd.n10837 vdd.n10831 8.533
R44607 vdd.n12328 vdd.n10853 8.533
R44608 vdd.n10878 vdd.n10877 8.533
R44609 vdd.n10889 vdd.n10888 8.533
R44610 vdd.n12314 vdd.n12313 8.533
R44611 vdd.n12303 vdd.n12302 8.533
R44612 vdd.n12297 vdd.n10900 8.533
R44613 vdd.n10931 vdd.n10930 8.533
R44614 vdd.n10942 vdd.n10941 8.533
R44615 vdd.n12283 vdd.n12282 8.533
R44616 vdd.n12275 vdd.n10924 8.533
R44617 vdd.n10974 vdd.n10973 8.533
R44618 vdd.n10981 vdd.n10980 8.533
R44619 vdd.n10989 vdd.n10963 8.533
R44620 vdd.n12256 vdd.n12255 8.533
R44621 vdd.n10998 vdd.n10996 8.533
R44622 vdd.n11022 vdd.n11021 8.533
R44623 vdd.n12231 vdd.n12230 8.533
R44624 vdd.n12220 vdd.n12219 8.533
R44625 vdd.n12214 vdd.n11040 8.533
R44626 vdd.n11068 vdd.n11067 8.533
R44627 vdd.n11079 vdd.n11078 8.533
R44628 vdd.n12200 vdd.n12199 8.533
R44629 vdd.n12189 vdd.n12188 8.533
R44630 vdd.n12183 vdd.n11090 8.533
R44631 vdd.n11115 vdd.n11092 8.533
R44632 vdd.n11123 vdd.n11109 8.533
R44633 vdd.n12166 vdd.n12165 8.533
R44634 vdd.n11132 vdd.n11130 8.533
R44635 vdd.n11159 vdd.n11158 8.533
R44636 vdd.n11166 vdd.n11165 8.533
R44637 vdd.n11173 vdd.n11149 8.533
R44638 vdd.n12137 vdd.n12136 8.533
R44639 vdd.n11203 vdd.n11202 8.533
R44640 vdd.n11214 vdd.n11213 8.533
R44641 vdd.n12112 vdd.n12111 8.533
R44642 vdd.n12101 vdd.n12100 8.533
R44643 vdd.n12095 vdd.n11225 8.533
R44644 vdd.n11252 vdd.n11251 8.533
R44645 vdd.n11263 vdd.n11262 8.533
R44646 vdd.n12081 vdd.n12080 8.533
R44647 vdd.n12070 vdd.n11268 8.533
R44648 vdd.n11296 vdd.n11295 8.533
R44649 vdd.n11303 vdd.n11302 8.533
R44650 vdd.n11311 vdd.n11285 8.533
R44651 vdd.n12051 vdd.n12050 8.533
R44652 vdd.n11320 vdd.n11318 8.533
R44653 vdd.n11344 vdd.n11343 8.533
R44654 vdd.n11346 vdd.n11340 8.533
R44655 vdd.n12022 vdd.n11362 8.533
R44656 vdd.n11387 vdd.n11386 8.533
R44657 vdd.n11398 vdd.n11397 8.533
R44658 vdd.n12008 vdd.n12007 8.533
R44659 vdd.n11997 vdd.n11996 8.533
R44660 vdd.n11991 vdd.n11409 8.533
R44661 vdd.n11475 vdd.n11474 8.533
R44662 vdd.n11486 vdd.n11485 8.533
R44663 vdd.n11977 vdd.n11976 8.533
R44664 vdd.n11969 vdd.n11433 8.533
R44665 vdd.n11506 vdd.n11505 8.533
R44666 vdd.n11949 vdd.n11948 8.533
R44667 vdd.n11937 vdd.n11936 8.533
R44668 vdd.n18387 vdd.n18386 8.533
R44669 vdd.n10555 vdd.n10536 8.489
R44670 vdd.n10644 vdd.n10631 8.489
R44671 vdd.n10712 vdd.n10706 8.489
R44672 vdd.n12355 vdd.n10806 8.489
R44673 vdd.n12316 vdd.n10869 8.489
R44674 vdd.n12262 vdd.n10961 8.489
R44675 vdd.n11065 vdd.n11044 8.489
R44676 vdd.n11139 vdd.n11136 8.489
R44677 vdd.n12102 vdd.n11220 8.489
R44678 vdd.n12049 vdd.n11315 8.489
R44679 vdd.n12010 vdd.n11378 8.489
R44680 vdd.n11956 vdd.n11446 8.489
R44681 vdd.n10406 vdd.n10321 8.489
R44682 vdd.n13075 vdd.n9292 8.489
R44683 vdd.n13015 vdd.n9398 8.489
R44684 vdd.n12964 vdd.n9462 8.489
R44685 vdd.n9580 vdd.n9563 8.489
R44686 vdd.n12867 vdd.n9624 8.489
R44687 vdd.n12807 vdd.n9758 8.489
R44688 vdd.n12756 vdd.n9822 8.489
R44689 vdd.n9940 vdd.n9921 8.489
R44690 vdd.n12659 vdd.n9984 8.489
R44691 vdd.n10109 vdd.n10108 8.489
R44692 vdd.n16894 vdd.n16893 8.489
R44693 vdd.n17050 vdd.n17049 8.489
R44694 vdd.n17166 vdd.n17165 8.489
R44695 vdd.n17322 vdd.n17321 8.489
R44696 vdd.n17438 vdd.n17437 8.489
R44697 vdd.n16829 vdd.n16828 8.489
R44698 vdd.n17696 vdd.n17695 8.489
R44699 vdd.n17852 vdd.n17851 8.489
R44700 vdd.n17967 vdd.n17966 8.489
R44701 vdd.n18123 vdd.n18122 8.489
R44702 vdd.n18238 vdd.n18237 8.489
R44703 vdd.n15020 vdd.n15019 8.489
R44704 vdd.n15382 vdd.n15378 8.489
R44705 vdd.n15462 vdd.n15452 8.489
R44706 vdd.n15627 vdd.n15620 8.489
R44707 vdd.n15718 vdd.n15708 8.489
R44708 vdd.n15883 vdd.n15876 8.489
R44709 vdd.n15974 vdd.n15964 8.489
R44710 vdd.n16139 vdd.n16132 8.489
R44711 vdd.n16230 vdd.n16220 8.489
R44712 vdd.n16395 vdd.n16388 8.489
R44713 vdd.n16486 vdd.n16476 8.489
R44714 vdd.n16623 vdd.n16622 8.489
R44715 vdd.n25396 vdd.n25377 8.465
R44716 vdd.n10600 vdd.n10599 8.45
R44717 vdd.n10599 vdd.n10598 8.45
R44718 vdd.n10751 vdd.n10750 8.45
R44719 vdd.n10750 vdd.n10749 8.45
R44720 vdd.n10919 vdd.n10916 8.45
R44721 vdd.n12286 vdd.n10916 8.45
R44722 vdd.n12181 vdd.n12180 8.45
R44723 vdd.n12180 vdd.n12179 8.45
R44724 vdd.n12076 vdd.n12075 8.45
R44725 vdd.n12075 vdd.n12074 8.45
R44726 vdd.n11428 vdd.n11425 8.45
R44727 vdd.n11980 vdd.n11425 8.45
R44728 vdd.n16978 vdd.n16977 8.45
R44729 vdd.n16977 vdd.n16976 8.45
R44730 vdd.n17250 vdd.n17249 8.45
R44731 vdd.n17249 vdd.n17248 8.45
R44732 vdd.n17522 vdd.n17521 8.45
R44733 vdd.n17521 vdd.n17520 8.45
R44734 vdd.n17780 vdd.n17779 8.45
R44735 vdd.n17779 vdd.n17778 8.45
R44736 vdd.n18051 vdd.n18050 8.45
R44737 vdd.n18050 vdd.n18049 8.45
R44738 vdd.n16817 vdd.n16816 8.45
R44739 vdd.n16816 vdd.n16815 8.45
R44740 vdd.n21616 vdd.n21615 8.444
R44741 vdd.n21430 vdd.n21429 8.444
R44742 vdd.n21349 vdd.n21348 8.444
R44743 vdd.n21183 vdd.t349 8.444
R44744 vdd.n21171 vdd.n21170 8.444
R44745 vdd.n21086 vdd.n21085 8.444
R44746 vdd.n19064 vdd.n19063 8.444
R44747 vdd.n18983 vdd.n18982 8.444
R44748 vdd.n18963 vdd.t281 8.444
R44749 vdd.n18805 vdd.n18804 8.444
R44750 vdd.n18724 vdd.n18723 8.444
R44751 vdd.n18546 vdd.n18545 8.444
R44752 vdd.n9342 vdd.n9328 8.344
R44753 vdd.n12994 vdd.n9414 8.344
R44754 vdd.n12936 vdd.n9518 8.344
R44755 vdd.n12935 vdd.n9519 8.344
R44756 vdd.n12887 vdd.n9610 8.344
R44757 vdd.n9702 vdd.n9688 8.344
R44758 vdd.n12835 vdd.n12834 8.344
R44759 vdd.n12786 vdd.n9775 8.344
R44760 vdd.n12728 vdd.n9878 8.344
R44761 vdd.n12727 vdd.n9879 8.344
R44762 vdd.n12679 vdd.n9970 8.344
R44763 vdd.n10156 vdd.n10155 8.344
R44764 vdd.n12627 vdd.n12626 8.344
R44765 vdd.n12588 vdd.n10118 8.344
R44766 vdd.n15530 vdd.n15527 8.344
R44767 vdd.n15786 vdd.n15783 8.344
R44768 vdd.n15807 vdd.n15806 8.344
R44769 vdd.n15200 vdd.n15199 8.344
R44770 vdd.n16042 vdd.n16039 8.344
R44771 vdd.n16063 vdd.n16062 8.344
R44772 vdd.n16298 vdd.n16295 8.344
R44773 vdd.n16319 vdd.n16318 8.344
R44774 vdd.n16570 vdd.n16564 8.344
R44775 vdd.n16563 vdd.n16561 8.344
R44776 vdd.n16662 vdd.n16661 8.344
R44777 vdd.n10682 vdd.n10681 8.296
R44778 vdd.n10681 vdd.n10680 8.296
R44779 vdd.n12333 vdd.n10828 8.296
R44780 vdd.n12333 vdd.n12332 8.296
R44781 vdd.n11030 vdd.n11018 8.296
R44782 vdd.n11031 vdd.n11030 8.296
R44783 vdd.n11181 vdd.n11179 8.296
R44784 vdd.n12125 vdd.n11181 8.296
R44785 vdd.n12027 vdd.n11337 8.296
R44786 vdd.n12027 vdd.n12026 8.296
R44787 vdd.n17126 vdd.n17110 8.296
R44788 vdd.n17398 vdd.n17382 8.296
R44789 vdd.n17656 vdd.n17640 8.296
R44790 vdd.n17927 vdd.n17911 8.296
R44791 vdd.n18199 vdd.n18183 8.296
R44792 vdd.n2682 vdd.n2681 8.282
R44793 vdd.n14265 vdd.t114 8.258
R44794 vdd.n19399 vdd.n19398 8.209
R44795 vdd.n19448 vdd.n19447 8.209
R44796 vdd.n19605 vdd.n19604 8.209
R44797 vdd.n19648 vdd.n19647 8.209
R44798 vdd.n20856 vdd.n20855 8.209
R44799 vdd.n20813 vdd.n20812 8.209
R44800 vdd.n20657 vdd.n20656 8.209
R44801 vdd.n20608 vdd.n20607 8.209
R44802 vdd.n20281 vdd.n20280 8.209
R44803 vdd.n20263 vdd.n20260 8.209
R44804 vdd.n14789 vdd.n8072 8.189
R44805 vdd.n14801 vdd.n14800 8.189
R44806 vdd.n33834 vdd.n33833 8.128
R44807 vdd.n809 vdd.n808 8.128
R44808 vdd.n11661 vdd.n9287 8.06
R44809 vdd.n21742 vdd.n15006 8.06
R44810 vdd.n10446 vdd.n10294 8.059
R44811 vdd.n10446 vdd.n10445 8.059
R44812 vdd.n9347 vdd.n9332 8.059
R44813 vdd.n13040 vdd.n9332 8.059
R44814 vdd.n12938 vdd.n9516 8.059
R44815 vdd.n9531 vdd.n9516 8.059
R44816 vdd.n9707 vdd.n9692 8.059
R44817 vdd.n12832 vdd.n9692 8.059
R44818 vdd.n12730 vdd.n9876 8.059
R44819 vdd.n9892 vdd.n9876 8.059
R44820 vdd.n11537 vdd.n11448 8.059
R44821 vdd.n15312 vdd.n15310 8.059
R44822 vdd.n15312 vdd.n15311 8.059
R44823 vdd.n15540 vdd.n15538 8.059
R44824 vdd.n15540 vdd.n15539 8.059
R44825 vdd.n15796 vdd.n15794 8.059
R44826 vdd.n15796 vdd.n15795 8.059
R44827 vdd.n16052 vdd.n16050 8.059
R44828 vdd.n16052 vdd.n16051 8.059
R44829 vdd.n16308 vdd.n16306 8.059
R44830 vdd.n16308 vdd.n16307 8.059
R44831 vdd.n9441 vdd.n9440 8.023
R44832 vdd.n12889 vdd.n9609 8.023
R44833 vdd.n9800 vdd.n9799 8.023
R44834 vdd.n12681 vdd.n9969 8.023
R44835 vdd.n10243 vdd.n10242 8.023
R44836 vdd.n15230 vdd.n15227 8.023
R44837 vdd.n15202 vdd.n15187 8.023
R44838 vdd.n15174 vdd.n15171 8.023
R44839 vdd.n15146 vdd.n15143 8.023
R44840 vdd.n16664 vdd.n16652 8.023
R44841 vdd.t328 vdd.n8874 7.952
R44842 vdd.n31021 vdd.n31020 7.905
R44843 vdd.n36017 vdd.n36013 7.862
R44844 vdd.n36059 vdd.n36055 7.862
R44845 vdd.n36248 vdd.n36244 7.862
R44846 vdd.n36290 vdd.n36286 7.862
R44847 vdd.n36479 vdd.n36475 7.862
R44848 vdd.n36521 vdd.n36517 7.862
R44849 vdd.n36710 vdd.n36706 7.862
R44850 vdd.n36752 vdd.n36748 7.862
R44851 vdd.n36941 vdd.n36937 7.862
R44852 vdd.n35685 vdd.n35684 7.862
R44853 vdd.n37149 vdd.n37145 7.862
R44854 vdd.n37177 vdd.n37173 7.862
R44855 vdd.n32990 vdd.n32986 7.862
R44856 vdd.n32976 vdd.n32972 7.862
R44857 vdd.n37524 vdd.n37520 7.862
R44858 vdd.n37570 vdd.n37566 7.862
R44859 vdd.n38038 vdd.n38034 7.862
R44860 vdd.n37996 vdd.n37992 7.862
R44861 vdd.n37807 vdd.n37803 7.862
R44862 vdd.n37765 vdd.n37761 7.862
R44863 vdd.n28207 vdd.n28203 7.862
R44864 vdd.n28249 vdd.n28245 7.862
R44865 vdd.n28438 vdd.n28434 7.862
R44866 vdd.n28480 vdd.n28476 7.862
R44867 vdd.n28669 vdd.n28665 7.862
R44868 vdd.n28711 vdd.n28707 7.862
R44869 vdd.n28114 vdd.n28110 7.862
R44870 vdd.n28088 vdd.n28084 7.862
R44871 vdd.n31628 vdd.n31627 7.862
R44872 vdd.n32066 vdd.n32065 7.862
R44873 vdd.n29722 vdd.n29718 7.862
R44874 vdd.n30190 vdd.n30186 7.862
R44875 vdd.n2875 vdd.n2874 7.862
R44876 vdd.n2907 vdd.n2906 7.862
R44877 vdd.n3056 vdd.n3055 7.862
R44878 vdd.n3088 vdd.n3087 7.862
R44879 vdd.n3237 vdd.n3236 7.862
R44880 vdd.n3269 vdd.n3268 7.862
R44881 vdd.n3418 vdd.n3417 7.862
R44882 vdd.n3450 vdd.n3449 7.862
R44883 vdd.n3599 vdd.n3598 7.862
R44884 vdd.n3644 vdd.n3640 7.862
R44885 vdd.n3919 vdd.n3918 7.862
R44886 vdd.n3853 vdd.n3852 7.862
R44887 vdd.n2419 vdd.n2418 7.862
R44888 vdd.n2478 vdd.n2477 7.862
R44889 vdd.n1864 vdd.n1863 7.862
R44890 vdd.n1797 vdd.n1796 7.862
R44891 vdd.n1669 vdd.n1668 7.862
R44892 vdd.n1637 vdd.n1636 7.862
R44893 vdd.n1488 vdd.n1487 7.862
R44894 vdd.n1456 vdd.n1455 7.862
R44895 vdd.n1307 vdd.n1306 7.862
R44896 vdd.n26773 vdd.n26772 7.862
R44897 vdd.n26922 vdd.n26921 7.862
R44898 vdd.n26954 vdd.n26953 7.862
R44899 vdd.n27103 vdd.n27102 7.862
R44900 vdd.n27135 vdd.n27134 7.862
R44901 vdd.n26618 vdd.n26617 7.862
R44902 vdd.n26346 vdd.n26345 7.862
R44903 vdd.n31630 vdd.n31623 7.862
R44904 vdd.n32068 vdd.n32061 7.862
R44905 vdd.n31474 vdd.n31473 7.862
R44906 vdd.n32505 vdd.n32504 7.862
R44907 vdd.n9124 vdd.n9068 7.862
R44908 vdd.n13392 vdd.n9053 7.862
R44909 vdd.n8903 vdd.n8848 7.862
R44910 vdd.n13684 vdd.n8833 7.862
R44911 vdd.n13914 vdd.n8659 7.862
R44912 vdd.n13978 vdd.n8602 7.862
R44913 vdd.n14204 vdd.n8439 7.862
R44914 vdd.n14268 vdd.n8380 7.862
R44915 vdd.n14694 vdd.n8126 7.862
R44916 vdd.n14740 vdd.n8107 7.862
R44917 vdd.n14868 vdd.n8036 7.862
R44918 vdd.n14893 vdd.n14885 7.862
R44919 vdd.n13220 vdd.n9202 7.862
R44920 vdd.n13305 vdd.n9139 7.862
R44921 vdd.n13512 vdd.n8980 7.862
R44922 vdd.n13597 vdd.n8917 7.862
R44923 vdd.n13811 vdd.n8748 7.862
R44924 vdd.n13878 vdd.n8702 7.862
R44925 vdd.n14098 vdd.n8534 7.862
R44926 vdd.n14167 vdd.n8479 7.862
R44927 vdd.n14393 vdd.n8306 7.862
R44928 vdd.n14450 vdd.n8263 7.862
R44929 vdd.n19280 vdd.n19274 7.862
R44930 vdd.n19244 vdd.n19238 7.862
R44931 vdd.n19224 vdd.n19218 7.862
R44932 vdd.n19187 vdd.n19181 7.862
R44933 vdd.n19841 vdd.n19835 7.862
R44934 vdd.n19878 vdd.n19872 7.862
R44935 vdd.n19910 vdd.n19904 7.862
R44936 vdd.n19946 vdd.n19940 7.862
R44937 vdd.n21545 vdd.n21539 7.862
R44938 vdd.n21495 vdd.n21489 7.862
R44939 vdd.n21286 vdd.n21280 7.862
R44940 vdd.n21236 vdd.n21230 7.862
R44941 vdd.n21027 vdd.n21023 7.862
R44942 vdd.n19128 vdd.n19123 7.862
R44943 vdd.n18920 vdd.n18914 7.862
R44944 vdd.n18870 vdd.n18864 7.862
R44945 vdd.n18661 vdd.n18655 7.862
R44946 vdd.n18611 vdd.n18605 7.862
R44947 vdd.n20415 vdd.n20414 7.862
R44948 vdd.n20357 vdd.n20356 7.862
R44949 vdd.n20179 vdd.n20178 7.862
R44950 vdd.n20121 vdd.n20120 7.862
R44951 vdd.n24766 vdd.n24765 7.862
R44952 vdd.n25144 vdd.n25143 7.862
R44953 vdd.n10443 vdd.t295 7.744
R44954 vdd.n15321 vdd.t263 7.744
R44955 vdd.n21559 vdd.n21556 7.74
R44956 vdd.n21477 vdd.n21474 7.74
R44957 vdd.n21218 vdd.n21215 7.74
R44958 vdd.n21041 vdd.n21038 7.74
R44959 vdd.n19111 vdd.n19108 7.74
R44960 vdd.n18934 vdd.n18931 7.74
R44961 vdd.n18675 vdd.n18672 7.74
R44962 vdd.n18593 vdd.n18590 7.74
R44963 vdd.t296 vdd.n13073 7.702
R44964 vdd.n13049 vdd.n9318 7.702
R44965 vdd.n13043 vdd.t225 7.702
R44966 vdd.n12948 vdd.n12947 7.702
R44967 vdd.n12841 vdd.n9680 7.702
R44968 vdd.n12740 vdd.n12739 7.702
R44969 vdd.n12633 vdd.t299 7.702
R44970 vdd.n12627 vdd.t372 7.702
R44971 vdd.n12132 vdd.t383 7.702
R44972 vdd.t249 vdd.n15460 7.702
R44973 vdd.t195 vdd.n15550 7.702
R44974 vdd.t14 vdd.n16563 7.702
R44975 vdd.n17904 vdd.t30 7.702
R44976 vdd.n11781 vdd.n11778 7.67
R44977 vdd.n11885 vdd.n11884 7.668
R44978 vdd.n21976 vdd.n21975 7.668
R44979 vdd.n14021 vdd.t124 7.646
R44980 vdd.t305 vdd.n8134 7.632
R44981 vdd.n19278 vdd.n19275 7.623
R44982 vdd.n19242 vdd.n19239 7.623
R44983 vdd.n19222 vdd.n19219 7.623
R44984 vdd.n19185 vdd.n19182 7.623
R44985 vdd.n19839 vdd.n19836 7.623
R44986 vdd.n19876 vdd.n19873 7.623
R44987 vdd.n19908 vdd.n19905 7.623
R44988 vdd.n19944 vdd.n19941 7.623
R44989 vdd.n20420 vdd.n20419 7.623
R44990 vdd.n20362 vdd.n20361 7.623
R44991 vdd.n20184 vdd.n20183 7.623
R44992 vdd.n20126 vdd.n20125 7.623
R44993 vdd.n14695 vdd.n8125 7.604
R44994 vdd.n14741 vdd.n8104 7.604
R44995 vdd.n14869 vdd.n8035 7.604
R44996 vdd.n14896 vdd.n14895 7.604
R44997 vdd.n10235 vdd.n10234 7.597
R44998 vdd.n11516 vdd.n11457 7.585
R44999 vdd.n24702 vdd.n24701 7.542
R45000 vdd.n25209 vdd.n25208 7.542
R45001 vdd.n24701 vdd.n24700 7.542
R45002 vdd.n25208 vdd.n25207 7.542
R45003 vdd.n11624 vdd.n11582 7.529
R45004 vdd.n21635 vdd.n21634 7.529
R45005 vdd.n11729 vdd.n11724 7.498
R45006 vdd.n11885 vdd.n11882 7.474
R45007 vdd.n21976 vdd.n21973 7.474
R45008 vdd.n12899 vdd.n12898 7.381
R45009 vdd.n12792 vdd.n9769 7.381
R45010 vdd.n12691 vdd.n12690 7.381
R45011 vdd.n12594 vdd.n10103 7.381
R45012 vdd.n15916 vdd.n15913 7.381
R45013 vdd.n16172 vdd.n16169 7.381
R45014 vdd.n16428 vdd.n16425 7.381
R45015 vdd.n16643 vdd.n16640 7.381
R45016 vdd.n11674 vdd.n11670 7.376
R45017 vdd.n362 vdd.n361 7.375
R45018 vdd.n13366 vdd.t120 7.34
R45019 vdd.t114 vdd.n8371 7.34
R45020 vdd.t322 vdd.n8183 7.34
R45021 vdd.n12504 vdd.n10563 7.276
R45022 vdd.n12462 vdd.n10612 7.276
R45023 vdd.n10736 vdd.n10727 7.276
R45024 vdd.n10799 vdd.n10782 7.276
R45025 vdd.n10908 vdd.n10897 7.276
R45026 vdd.n10969 vdd.n10953 7.276
R45027 vdd.n12202 vdd.n11058 7.276
R45028 vdd.n12160 vdd.n11127 7.276
R45029 vdd.n12092 vdd.n11229 7.276
R45030 vdd.n11308 vdd.n11290 7.276
R45031 vdd.n11417 vdd.n11406 7.276
R45032 vdd.n11523 vdd.n11438 7.276
R45033 vdd.n10469 vdd.n10273 7.276
R45034 vdd.n10317 vdd.n10314 7.276
R45035 vdd.n13062 vdd.n9307 7.276
R45036 vdd.n9387 vdd.n9361 7.276
R45037 vdd.n9500 vdd.n9482 7.276
R45038 vdd.n12916 vdd.n9553 7.276
R45039 vdd.n12854 vdd.n9667 7.276
R45040 vdd.n9747 vdd.n9721 7.276
R45041 vdd.n9860 vdd.n9842 7.276
R45042 vdd.n12708 vdd.n9913 7.276
R45043 vdd.n12646 vdd.n10027 7.276
R45044 vdd.n10192 vdd.n10063 7.276
R45045 vdd.n16932 vdd.n16926 7.276
R45046 vdd.n17024 vdd.n17018 7.276
R45047 vdd.n17204 vdd.n17198 7.276
R45048 vdd.n17296 vdd.n17290 7.276
R45049 vdd.n17476 vdd.n17470 7.276
R45050 vdd.n17568 vdd.n17562 7.276
R45051 vdd.n17734 vdd.n17728 7.276
R45052 vdd.n17826 vdd.n17820 7.276
R45053 vdd.n18005 vdd.n17999 7.276
R45054 vdd.n18097 vdd.n18091 7.276
R45055 vdd.n18273 vdd.n18268 7.276
R45056 vdd.n18345 vdd.n18340 7.276
R45057 vdd.n15270 vdd.n15269 7.276
R45058 vdd.n15349 vdd.n15348 7.276
R45059 vdd.n15489 vdd.n15488 7.276
R45060 vdd.n15586 vdd.n15585 7.276
R45061 vdd.n15745 vdd.n15744 7.276
R45062 vdd.n15842 vdd.n15841 7.276
R45063 vdd.n16001 vdd.n16000 7.276
R45064 vdd.n16098 vdd.n16097 7.276
R45065 vdd.n16257 vdd.n16256 7.276
R45066 vdd.n16354 vdd.n16353 7.276
R45067 vdd.n16513 vdd.n16512 7.276
R45068 vdd.n16727 vdd.n16726 7.276
R45069 vdd.n9320 vdd.n9319 7.06
R45070 vdd.n12956 vdd.n12955 7.06
R45071 vdd.n9678 vdd.n9669 7.06
R45072 vdd.n12748 vdd.n12747 7.06
R45073 vdd.n10038 vdd.n10029 7.06
R45074 vdd.n12278 vdd.t385 7.06
R45075 vdd.n17535 vdd.t4 7.06
R45076 vdd.n24098 vdd.n24097 7.058
R45077 vdd.n24072 vdd.n24071 7.058
R45078 vdd.n23866 vdd.n23865 7.058
R45079 vdd.n23840 vdd.n23839 7.058
R45080 vdd.n23634 vdd.n23633 7.058
R45081 vdd.n23152 vdd.n23151 7.058
R45082 vdd.n23178 vdd.n23177 7.058
R45083 vdd.n23384 vdd.n23383 7.058
R45084 vdd.n23410 vdd.n23409 7.058
R45085 vdd.n23616 vdd.n23615 7.058
R45086 vdd.n22573 vdd.n22572 7.058
R45087 vdd.n22599 vdd.n22598 7.058
R45088 vdd.n22805 vdd.n22804 7.058
R45089 vdd.n22831 vdd.n22830 7.058
R45090 vdd.n23037 vdd.n23036 7.058
R45091 vdd.n22189 vdd.n22188 7.058
R45092 vdd.n22047 vdd.n22046 7.058
R45093 vdd.n22168 vdd.n22167 7.058
R45094 vdd.n21592 vdd.n21591 7.037
R45095 vdd.n21446 vdd.n21445 7.037
R45096 vdd.n21333 vdd.n21332 7.037
R45097 vdd.t276 vdd.n21247 7.037
R45098 vdd.n21187 vdd.n21186 7.037
R45099 vdd.n21074 vdd.n21073 7.037
R45100 vdd.n19080 vdd.n19079 7.037
R45101 vdd.n18967 vdd.n18966 7.037
R45102 vdd.t344 vdd.n18899 7.037
R45103 vdd.n18821 vdd.n18820 7.037
R45104 vdd.n18708 vdd.n18707 7.037
R45105 vdd.n18562 vdd.n18561 7.037
R45106 vdd.n19383 vdd.n19382 7.037
R45107 vdd.n19464 vdd.n19463 7.037
R45108 vdd.n19664 vdd.n19663 7.037
R45109 vdd.n19791 vdd.n19790 7.037
R45110 vdd.n20988 vdd.n20987 7.037
R45111 vdd.n19890 vdd.n19889 7.037
R45112 vdd.n20673 vdd.n20672 7.037
R45113 vdd.n20592 vdd.n20591 7.037
R45114 vdd.n20472 vdd.n20471 7.037
R45115 vdd.n20297 vdd.n20296 7.037
R45116 vdd.n20247 vdd.n20244 7.037
R45117 vdd.n20061 vdd.n20060 7.037
R45118 vdd.t335 vdd.n13376 7.034
R45119 vdd.n14302 vdd.t287 7.034
R45120 vdd.n14773 vdd.n8083 7.019
R45121 vdd.n14828 vdd.n8054 7.019
R45122 vdd.n14942 vdd.n7987 7.019
R45123 vdd.n9099 vdd.t107 6.923
R45124 vdd.n9099 vdd.t121 6.923
R45125 vdd.n13417 vdd.t119 6.923
R45126 vdd.n13417 vdd.t117 6.923
R45127 vdd.n8940 vdd.t127 6.923
R45128 vdd.n8940 vdd.t137 6.923
R45129 vdd.n8831 vdd.t135 6.923
R45130 vdd.n8831 vdd.t129 6.923
R45131 vdd.n8661 vdd.t111 6.923
R45132 vdd.n8661 vdd.t109 6.923
R45133 vdd.n14043 vdd.t125 6.923
R45134 vdd.n14043 vdd.t123 6.923
R45135 vdd.n8464 vdd.t133 6.923
R45136 vdd.n8464 vdd.t131 6.923
R45137 vdd.n8352 vdd.t115 6.923
R45138 vdd.n8352 vdd.t103 6.923
R45139 vdd.n13784 vdd.t105 6.923
R45140 vdd.n13784 vdd.t113 6.923
R45141 vdd.n19283 vdd.t153 6.923
R45142 vdd.n19283 vdd.t141 6.923
R45143 vdd.n19234 vdd.t171 6.923
R45144 vdd.n19234 vdd.t165 6.923
R45145 vdd.n19227 vdd.t155 6.923
R45146 vdd.n19227 vdd.t159 6.923
R45147 vdd.n19190 vdd.t143 6.923
R45148 vdd.n19190 vdd.t145 6.923
R45149 vdd.n19844 vdd.t163 6.923
R45150 vdd.n19844 vdd.t147 6.923
R45151 vdd.n19881 vdd.t149 6.923
R45152 vdd.n19881 vdd.t173 6.923
R45153 vdd.n19899 vdd.t175 6.923
R45154 vdd.n19899 vdd.t167 6.923
R45155 vdd.n19949 vdd.t151 6.923
R45156 vdd.n19949 vdd.t157 6.923
R45157 vdd.n19828 vdd.t169 6.923
R45158 vdd.n19828 vdd.t161 6.923
R45159 vdd.n24521 vdd.t239 6.923
R45160 vdd.n24538 vdd.t202 6.923
R45161 vdd.n24538 vdd.t338 6.923
R45162 vdd.n24960 vdd.t343 6.923
R45163 vdd.n24960 vdd.t342 6.923
R45164 vdd.n24887 vdd.t340 6.923
R45165 vdd.n24887 vdd.t236 6.923
R45166 vdd.n25023 vdd.t237 6.923
R45167 vdd.n25023 vdd.t206 6.923
R45168 vdd.n24922 vdd.t207 6.923
R45169 vdd.n24633 vdd.t240 6.923
R45170 vdd.n24633 vdd.t201 6.923
R45171 vdd.n10235 vdd.n10227 6.874
R45172 vdd.n13136 vdd.n13135 6.776
R45173 vdd.n21686 vdd.n21685 6.776
R45174 vdd.n9406 vdd.n9401 6.739
R45175 vdd.n9595 vdd.n9594 6.739
R45176 vdd.n9766 vdd.n9761 6.739
R45177 vdd.n9955 vdd.n9954 6.739
R45178 vdd.n10112 vdd.n10102 6.739
R45179 vdd.t291 vdd.n11376 6.739
R45180 vdd.n15643 vdd.n15640 6.739
R45181 vdd.n15899 vdd.n15896 6.739
R45182 vdd.n16155 vdd.n16152 6.739
R45183 vdd.n16411 vdd.n16408 6.739
R45184 vdd.n16632 vdd.n16628 6.739
R45185 vdd.n8664 vdd.t331 6.728
R45186 vdd.n11468 vdd.n10260 6.639
R45187 vdd.n16797 vdd.n16796 6.639
R45188 vdd.n34204 vdd.n34203 6.622
R45189 vdd.n35288 vdd.n35287 6.622
R45190 vdd.n34704 vdd.n34703 6.622
R45191 vdd.n5905 vdd.n5904 6.622
R45192 vdd.n5451 vdd.n5450 6.622
R45193 vdd.n4278 vdd.n4277 6.622
R45194 vdd.n27340 vdd.n27339 6.622
R45195 vdd.n25792 vdd.n25791 6.622
R45196 vdd.n11740 vdd.n11739 6.586
R45197 vdd.n11824 vdd.n11823 6.586
R45198 vdd.n21816 vdd.n21815 6.586
R45199 vdd.n21915 vdd.n21914 6.586
R45200 vdd.n19334 vdd.n19331 6.45
R45201 vdd.n19510 vdd.n19507 6.45
R45202 vdd.n19540 vdd.n19537 6.45
R45203 vdd.n19635 vdd.t154 6.45
R45204 vdd.n19696 vdd.t158 6.45
R45205 vdd.n19711 vdd.n19708 6.45
R45206 vdd.n19742 vdd.n19739 6.45
R45207 vdd.n20939 vdd.n20936 6.45
R45208 vdd.n20908 vdd.n20905 6.45
R45209 vdd.n20893 vdd.t148 6.45
R45210 vdd.n20843 vdd.t172 6.45
R45211 vdd.n20749 vdd.n20746 6.45
R45212 vdd.n20719 vdd.n20716 6.45
R45213 vdd.n20543 vdd.n20540 6.45
R45214 vdd.n20436 vdd.n20435 6.45
R45215 vdd.n20346 vdd.n20345 6.45
R45216 vdd.n20200 vdd.n20199 6.45
R45217 vdd.n20110 vdd.n20109 6.45
R45218 vdd.n14674 vdd.n14673 6.434
R45219 vdd.n14731 vdd.n14730 6.434
R45220 vdd.n14846 vdd.n14845 6.434
R45221 vdd.n14913 vdd.n8016 6.434
R45222 vdd.n13720 vdd.t128 6.423
R45223 vdd.n13061 vdd.n9308 6.418
R45224 vdd.n9498 vdd.n9497 6.418
R45225 vdd.n12853 vdd.n9668 6.418
R45226 vdd.n9858 vdd.n9857 6.418
R45227 vdd.n12645 vdd.n10028 6.418
R45228 vdd.n12624 vdd.n12623 6.4
R45229 vdd.n21575 vdd.n21572 6.333
R45230 vdd.n21461 vdd.n21458 6.333
R45231 vdd.n21316 vdd.n21313 6.333
R45232 vdd.n21300 vdd.t278 6.333
R45233 vdd.n21202 vdd.n21199 6.333
R45234 vdd.n21057 vdd.n21054 6.333
R45235 vdd.n19095 vdd.n19092 6.333
R45236 vdd.n18950 vdd.n18947 6.333
R45237 vdd.n18852 vdd.t346 6.333
R45238 vdd.n18836 vdd.n18833 6.333
R45239 vdd.n18691 vdd.n18688 6.333
R45240 vdd.n18577 vdd.n18574 6.333
R45241 vdd.n10478 vdd.n10271 6.273
R45242 vdd.n15258 vdd.n15257 6.273
R45243 vdd.n33823 vdd.n33822 6.259
R45244 vdd.n34190 vdd.n34189 6.259
R45245 vdd.n35300 vdd.n35299 6.259
R45246 vdd.n34716 vdd.n34715 6.259
R45247 vdd.n839 vdd.n838 6.259
R45248 vdd.n348 vdd.n347 6.259
R45249 vdd.n5891 vdd.n5890 6.259
R45250 vdd.n5463 vdd.n5462 6.259
R45251 vdd.n4893 vdd.n4892 6.259
R45252 vdd.n4290 vdd.n4289 6.259
R45253 vdd.n27328 vdd.n27327 6.259
R45254 vdd.n25780 vdd.n25779 6.259
R45255 vdd.n33714 vdd.n33712 6.246
R45256 vdd.n34087 vdd.n34085 6.246
R45257 vdd.n35248 vdd.n35246 6.246
R45258 vdd.n34661 vdd.n34659 6.246
R45259 vdd.n904 vdd.n902 6.246
R45260 vdd.n231 vdd.n229 6.246
R45261 vdd.n5789 vdd.n5787 6.246
R45262 vdd.n5408 vdd.n5406 6.246
R45263 vdd.n4813 vdd.n4811 6.246
R45264 vdd.n4238 vdd.n4236 6.246
R45265 vdd.n27294 vdd.n27292 6.246
R45266 vdd.n25746 vdd.n25744 6.246
R45267 vdd.n25638 vdd.n25637 6.211
R45268 vdd.n13213 vdd.n9173 6.208
R45269 vdd.n13254 vdd.n13253 6.208
R45270 vdd.n13506 vdd.n8953 6.208
R45271 vdd.n13545 vdd.n13544 6.208
R45272 vdd.n13787 vdd.n8734 6.208
R45273 vdd.n13830 vdd.n13829 6.208
R45274 vdd.n14115 vdd.n8516 6.208
R45275 vdd.n14110 vdd.n8518 6.208
R45276 vdd.n14399 vdd.n8299 6.208
R45277 vdd.n14403 vdd.n8277 6.208
R45278 vdd.n14792 vdd.n8067 6.208
R45279 vdd.n14797 vdd.n8066 6.208
R45280 vdd.n13382 vdd.n9058 6.208
R45281 vdd.n13386 vdd.n9024 6.208
R45282 vdd.n13674 vdd.n8838 6.208
R45283 vdd.n13678 vdd.n8804 6.208
R45284 vdd.n13950 vdd.n8597 6.208
R45285 vdd.n14001 vdd.n14000 6.208
R45286 vdd.n14240 vdd.n8375 6.208
R45287 vdd.n14292 vdd.n14291 6.208
R45288 vdd.n14605 vdd.n8177 6.208
R45289 vdd.n14610 vdd.n8176 6.208
R45290 vdd.n19173 vdd.n19172 6.208
R45291 vdd.n22153 vdd.n22142 6.143
R45292 vdd.n22164 vdd.n22154 6.143
R45293 vdd.n22185 vdd.n22175 6.143
R45294 vdd.n22268 vdd.n22257 6.143
R45295 vdd.n22279 vdd.n22269 6.143
R45296 vdd.n13647 vdd.t134 6.117
R45297 vdd.n8631 vdd.t108 6.117
R45298 vdd.n14233 vdd.t315 6.117
R45299 vdd.n27769 vdd.n27768 6.114
R45300 vdd.n11625 vdd.n11624 6.098
R45301 vdd.n21636 vdd.n21635 6.098
R45302 vdd.n13014 vdd.n9400 6.097
R45303 vdd.n12905 vdd.n9564 6.097
R45304 vdd.n12806 vdd.n9760 6.097
R45305 vdd.n10107 vdd.n10106 6.097
R45306 vdd.t368 vdd.n10574 6.097
R45307 vdd.n15626 vdd.n15623 6.097
R45308 vdd.n15882 vdd.n15879 6.097
R45309 vdd.n16138 vdd.n16135 6.097
R45310 vdd.n16624 vdd.n16620 6.097
R45311 vdd.n33811 vdd.n33810 6.088
R45312 vdd.n33655 vdd.n33654 6.088
R45313 vdd.n34175 vdd.n34174 6.088
R45314 vdd.n34306 vdd.n34305 6.088
R45315 vdd.n35320 vdd.n35319 6.088
R45316 vdd.n35572 vdd.n35571 6.088
R45317 vdd.n34725 vdd.n34724 6.088
R45318 vdd.n34901 vdd.n34900 6.088
R45319 vdd.n819 vdd.n818 6.088
R45320 vdd.n1071 vdd.n1070 6.088
R45321 vdd.n336 vdd.n335 6.088
R45322 vdd.n154 vdd.n153 6.088
R45323 vdd.n5878 vdd.n5877 6.088
R45324 vdd.n5944 vdd.n5943 6.088
R45325 vdd.n5472 vdd.n5471 6.088
R45326 vdd.n5648 vdd.n5647 6.088
R45327 vdd.n4914 vdd.n4913 6.088
R45328 vdd.n4632 vdd.n4631 6.088
R45329 vdd.n4299 vdd.n4298 6.088
R45330 vdd.n4475 vdd.n4474 6.088
R45331 vdd.n27317 vdd.n27316 6.088
R45332 vdd.n27440 vdd.n27439 6.088
R45333 vdd.n25769 vdd.n25768 6.088
R45334 vdd.n25886 vdd.n25885 6.088
R45335 vdd.n25648 vdd.n25647 6.088
R45336 vdd.n3662 vdd.n3661 6.088
R45337 vdd.n3668 vdd.n3667 6.088
R45338 vdd.n10537 vdd.n10524 6.063
R45339 vdd.n12452 vdd.n10624 6.063
R45340 vdd.n12412 vdd.n10699 6.063
R45341 vdd.n10814 vdd.n10808 6.063
R45342 vdd.n10887 vdd.n10874 6.063
R45343 vdd.n12254 vdd.n10993 6.063
R45344 vdd.n11049 vdd.n11043 6.063
R45345 vdd.n11167 vdd.n11154 6.063
R45346 vdd.n12114 vdd.n11194 6.063
R45347 vdd.n11323 vdd.n11317 6.063
R45348 vdd.n11396 vdd.n11383 6.063
R45349 vdd.n11947 vdd.n11548 6.063
R45350 vdd.n10402 vdd.n10327 6.063
R45351 vdd.n10367 vdd.n9291 6.063
R45352 vdd.n13003 vdd.n9402 6.063
R45353 vdd.n12971 vdd.n9453 6.063
R45354 vdd.n9597 vdd.n9578 6.063
R45355 vdd.n9650 vdd.n9623 6.063
R45356 vdd.n12795 vdd.n9762 6.063
R45357 vdd.n12763 vdd.n9812 6.063
R45358 vdd.n9957 vdd.n9937 6.063
R45359 vdd.n10010 vdd.n9983 6.063
R45360 vdd.n12596 vdd.n10099 6.063
R45361 vdd.n12568 vdd.n10270 6.063
R45362 vdd.n16878 vdd.n16877 6.063
R45363 vdd.n17066 vdd.n17065 6.063
R45364 vdd.n17150 vdd.n17149 6.063
R45365 vdd.n17338 vdd.n17337 6.063
R45366 vdd.n17422 vdd.n17421 6.063
R45367 vdd.n16823 vdd.n16822 6.063
R45368 vdd.n17680 vdd.n17679 6.063
R45369 vdd.n17868 vdd.n17867 6.063
R45370 vdd.n17951 vdd.n17950 6.063
R45371 vdd.n18139 vdd.n18138 6.063
R45372 vdd.n18223 vdd.n18222 6.063
R45373 vdd.n18397 vdd.n18396 6.063
R45374 vdd.n15396 vdd.n15392 6.063
R45375 vdd.n15442 vdd.n15438 6.063
R45376 vdd.n15644 vdd.n15637 6.063
R45377 vdd.n15698 vdd.n15691 6.063
R45378 vdd.n15900 vdd.n15893 6.063
R45379 vdd.n15954 vdd.n15947 6.063
R45380 vdd.n16156 vdd.n16149 6.063
R45381 vdd.n16210 vdd.n16203 6.063
R45382 vdd.n16412 vdd.n16405 6.063
R45383 vdd.n16466 vdd.n16459 6.063
R45384 vdd.n16631 vdd.n16630 6.063
R45385 vdd.n15117 vdd.n15071 6.063
R45386 vdd.n34430 vdd.n34429 6.023
R45387 vdd.n35388 vdd.n35387 6.023
R45388 vdd.n34860 vdd.n34859 6.023
R45389 vdd.n6081 vdd.n6080 6.023
R45390 vdd.n5607 vdd.n5606 6.023
R45391 vdd.n4722 vdd.n4721 6.023
R45392 vdd.n4434 vdd.n4433 6.023
R45393 vdd.n30300 vdd.n30292 6.023
R45394 vdd.n30568 vdd.n30561 6.023
R45395 vdd.n35913 vdd.n35906 6.023
R45396 vdd.n35934 vdd.n35926 6.023
R45397 vdd.n36144 vdd.n36137 6.023
R45398 vdd.n36165 vdd.n36157 6.023
R45399 vdd.n36375 vdd.n36368 6.023
R45400 vdd.n36396 vdd.n36388 6.023
R45401 vdd.n36606 vdd.n36599 6.023
R45402 vdd.n36627 vdd.n36619 6.023
R45403 vdd.n36837 vdd.n36830 6.023
R45404 vdd.n36858 vdd.n36850 6.023
R45405 vdd.n33268 vdd.n33261 6.023
R45406 vdd.n33250 vdd.n33242 6.023
R45407 vdd.n33074 vdd.n33067 6.023
R45408 vdd.n37260 vdd.n37252 6.023
R45409 vdd.n37446 vdd.n37438 6.023
R45410 vdd.n32914 vdd.n32907 6.023
R45411 vdd.n38125 vdd.n38118 6.023
R45412 vdd.n38136 vdd.n38128 6.023
R45413 vdd.n37913 vdd.n37905 6.023
R45414 vdd.n37892 vdd.n37885 6.023
R45415 vdd.n37682 vdd.n37674 6.023
R45416 vdd.n37661 vdd.n37654 6.023
R45417 vdd.n28334 vdd.n28327 6.023
R45418 vdd.n28355 vdd.n28347 6.023
R45419 vdd.n28565 vdd.n28558 6.023
R45420 vdd.n28586 vdd.n28578 6.023
R45421 vdd.n28796 vdd.n28789 6.023
R45422 vdd.n28153 vdd.n28145 6.023
R45423 vdd.n27768 vdd.n27760 6.023
R45424 vdd.n29694 vdd.n29686 6.023
R45425 vdd.n1739 vdd.n1735 6.023
R45426 vdd.n1746 vdd.n1742 6.023
R45427 vdd.n1572 vdd.n1568 6.023
R45428 vdd.n1555 vdd.n1551 6.023
R45429 vdd.n1391 vdd.n1387 6.023
R45430 vdd.n1374 vdd.n1370 6.023
R45431 vdd.n26840 vdd.n26836 6.023
R45432 vdd.n26857 vdd.n26853 6.023
R45433 vdd.n27021 vdd.n27017 6.023
R45434 vdd.n27038 vdd.n27034 6.023
R45435 vdd.n27202 vdd.n27198 6.023
R45436 vdd.n26745 vdd.n26741 6.023
R45437 vdd.n1979 vdd.n1975 6.023
R45438 vdd.n2793 vdd.n2789 6.023
R45439 vdd.n2810 vdd.n2806 6.023
R45440 vdd.n2974 vdd.n2970 6.023
R45441 vdd.n2991 vdd.n2987 6.023
R45442 vdd.n3155 vdd.n3151 6.023
R45443 vdd.n3172 vdd.n3168 6.023
R45444 vdd.n3336 vdd.n3332 6.023
R45445 vdd.n3353 vdd.n3349 6.023
R45446 vdd.n3517 vdd.n3513 6.023
R45447 vdd.n3534 vdd.n3530 6.023
R45448 vdd.n31893 vdd.n31883 6.023
R45449 vdd.n13214 vdd.n13213 6.023
R45450 vdd.n13253 vdd.n9175 6.023
R45451 vdd.n13507 vdd.n13506 6.023
R45452 vdd.n13544 vdd.n8955 6.023
R45453 vdd.n13788 vdd.n13787 6.023
R45454 vdd.n13829 vdd.n8736 6.023
R45455 vdd.n14116 vdd.n14115 6.023
R45456 vdd.n14110 vdd.n8521 6.023
R45457 vdd.n14399 vdd.n14398 6.023
R45458 vdd.n14428 vdd.n8277 6.023
R45459 vdd.n14785 vdd.n14784 6.023
R45460 vdd.n14783 vdd.n8078 6.023
R45461 vdd.n13143 vdd.n9248 6.023
R45462 vdd.n13382 vdd.n13381 6.023
R45463 vdd.n13436 vdd.n9024 6.023
R45464 vdd.n13674 vdd.n13673 6.023
R45465 vdd.n13728 vdd.n8804 6.023
R45466 vdd.n13952 vdd.n13950 6.023
R45467 vdd.n14000 vdd.n13995 6.023
R45468 vdd.n14242 vdd.n14240 6.023
R45469 vdd.n14291 vdd.n14286 6.023
R45470 vdd.n14605 vdd.n8179 6.023
R45471 vdd.n14612 vdd.n14610 6.023
R45472 vdd.n22144 vdd.n22143 6.023
R45473 vdd.n22156 vdd.n22155 6.023
R45474 vdd.n24194 vdd.n24193 6.023
R45475 vdd.n23972 vdd.n23971 6.023
R45476 vdd.n23962 vdd.n23961 6.023
R45477 vdd.n23740 vdd.n23739 6.023
R45478 vdd.n23730 vdd.n23729 6.023
R45479 vdd.n23052 vdd.n23051 6.023
R45480 vdd.n23274 vdd.n23273 6.023
R45481 vdd.n23284 vdd.n23283 6.023
R45482 vdd.n23506 vdd.n23505 6.023
R45483 vdd.n23516 vdd.n23515 6.023
R45484 vdd.n22473 vdd.n22472 6.023
R45485 vdd.n22695 vdd.n22694 6.023
R45486 vdd.n22705 vdd.n22704 6.023
R45487 vdd.n22927 vdd.n22926 6.023
R45488 vdd.n22937 vdd.n22936 6.023
R45489 vdd.n22177 vdd.n22176 6.023
R45490 vdd.n22259 vdd.n22258 6.023
R45491 vdd.n22271 vdd.n22270 6.023
R45492 vdd.n19420 vdd.n19408 6.023
R45493 vdd.n19434 vdd.n19425 6.023
R45494 vdd.n19623 vdd.n19611 6.023
R45495 vdd.n19637 vdd.n19628 6.023
R45496 vdd.n19825 vdd.n19813 6.023
R45497 vdd.n19172 vdd.n19163 6.023
R45498 vdd.n20845 vdd.n20833 6.023
R45499 vdd.n20828 vdd.n20819 6.023
R45500 vdd.n20643 vdd.n20631 6.023
R45501 vdd.n20626 vdd.n20617 6.023
R45502 vdd.n21675 vdd.n21655 6.023
R45503 vdd.n21400 vdd.n21388 6.023
R45504 vdd.n21383 vdd.n21374 6.023
R45505 vdd.n21141 vdd.n21129 6.023
R45506 vdd.n21124 vdd.n21115 6.023
R45507 vdd.n19034 vdd.n19022 6.023
R45508 vdd.n19017 vdd.n19008 6.023
R45509 vdd.n18775 vdd.n18763 6.023
R45510 vdd.n18758 vdd.n18749 6.023
R45511 vdd.n18516 vdd.n18504 6.023
R45512 vdd.n18499 vdd.n18463 6.023
R45513 vdd.n19991 vdd.n19990 6.023
R45514 vdd.n20003 vdd.n20002 6.023
R45515 vdd.n24410 vdd.n24409 6.023
R45516 vdd.n24978 vdd.n24977 6.023
R45517 vdd.n13369 vdd.n9065 6.009
R45518 vdd.n13400 vdd.n13399 6.009
R45519 vdd.n13661 vdd.n8845 6.009
R45520 vdd.n13693 vdd.n13692 6.009
R45521 vdd.n8668 vdd.n8667 6.009
R45522 vdd.n13981 vdd.n8609 6.009
R45523 vdd.n8445 vdd.n8444 6.009
R45524 vdd.n14271 vdd.n8387 6.009
R45525 vdd.n14681 vdd.n8117 6.009
R45526 vdd.n14710 vdd.n8115 6.009
R45527 vdd.n14855 vdd.n14854 6.009
R45528 vdd.n8026 vdd.n8024 6.009
R45529 vdd.n24890 vdd.n24889 5.966
R45530 vdd.n24541 vdd.n24540 5.965
R45531 vdd.n24963 vdd.n24962 5.965
R45532 vdd.n24925 vdd.n24924 5.965
R45533 vdd.n10081 vdd.n10054 5.925
R45534 vdd.n35894 vdd.n35893 5.896
R45535 vdd.n35943 vdd.n35942 5.896
R45536 vdd.n36125 vdd.n36124 5.896
R45537 vdd.n36174 vdd.n36173 5.896
R45538 vdd.n36356 vdd.n36355 5.896
R45539 vdd.n36405 vdd.n36404 5.896
R45540 vdd.n36587 vdd.n36586 5.896
R45541 vdd.n36636 vdd.n36635 5.896
R45542 vdd.n36818 vdd.n36817 5.896
R45543 vdd.n36867 vdd.n36866 5.896
R45544 vdd.n37053 vdd.n37052 5.896
R45545 vdd.n37092 vdd.n37091 5.896
R45546 vdd.n37226 vdd.n37225 5.896
R45547 vdd.n33054 vdd.n33053 5.896
R45548 vdd.n32924 vdd.n32923 5.896
R45549 vdd.n37465 vdd.n37464 5.896
R45550 vdd.n38147 vdd.n38146 5.896
R45551 vdd.n38104 vdd.n38103 5.896
R45552 vdd.n37922 vdd.n37921 5.896
R45553 vdd.n37873 vdd.n37872 5.896
R45554 vdd.n37691 vdd.n37690 5.896
R45555 vdd.n37642 vdd.n37641 5.896
R45556 vdd.n28315 vdd.n28314 5.896
R45557 vdd.n28364 vdd.n28363 5.896
R45558 vdd.n28546 vdd.n28545 5.896
R45559 vdd.n28595 vdd.n28594 5.896
R45560 vdd.n28777 vdd.n28776 5.896
R45561 vdd.n28160 vdd.n28159 5.896
R45562 vdd.n31844 vdd.n31843 5.896
R45563 vdd.n29025 vdd.n29024 5.896
R45564 vdd.n29867 vdd.n29866 5.896
R45565 vdd.n29833 vdd.n29832 5.896
R45566 vdd.n31092 vdd.n31091 5.896
R45567 vdd.n30542 vdd.n30541 5.896
R45568 vdd.n2780 vdd.n2779 5.896
R45569 vdd.n2819 vdd.n2818 5.896
R45570 vdd.n2961 vdd.n2960 5.896
R45571 vdd.n3000 vdd.n2999 5.896
R45572 vdd.n3142 vdd.n3141 5.896
R45573 vdd.n3181 vdd.n3180 5.896
R45574 vdd.n3323 vdd.n3322 5.896
R45575 vdd.n3362 vdd.n3361 5.896
R45576 vdd.n3504 vdd.n3503 5.896
R45577 vdd.n3543 vdd.n3542 5.896
R45578 vdd.n3689 vdd.n3688 5.896
R45579 vdd.n3994 vdd.n3993 5.896
R45580 vdd.n2153 vdd.n2152 5.896
R45581 vdd.n2319 vdd.n2318 5.896
R45582 vdd.n2565 vdd.n2564 5.896
R45583 vdd.n2070 vdd.n2069 5.896
R45584 vdd.n1756 vdd.n1755 5.896
R45585 vdd.n1723 vdd.n1722 5.896
R45586 vdd.n1581 vdd.n1580 5.896
R45587 vdd.n1542 vdd.n1541 5.896
R45588 vdd.n1400 vdd.n1399 5.896
R45589 vdd.n1361 vdd.n1360 5.896
R45590 vdd.n26827 vdd.n26826 5.896
R45591 vdd.n26866 vdd.n26865 5.896
R45592 vdd.n27008 vdd.n27007 5.896
R45593 vdd.n27047 vdd.n27046 5.896
R45594 vdd.n27189 vdd.n27188 5.896
R45595 vdd.n26735 vdd.n26734 5.896
R45596 vdd.n31840 vdd.n31839 5.896
R45597 vdd.n31909 vdd.n31908 5.896
R45598 vdd.n32201 vdd.n32200 5.896
R45599 vdd.n32281 vdd.n32280 5.896
R45600 vdd.n31088 vdd.n31087 5.896
R45601 vdd.n31266 vdd.n31265 5.896
R45602 vdd.n13178 vdd.n9208 5.896
R45603 vdd.n13267 vdd.n9160 5.896
R45604 vdd.n13473 vdd.n8987 5.896
R45605 vdd.n13559 vdd.n8938 5.896
R45606 vdd.n13779 vdd.n8772 5.896
R45607 vdd.n13841 vdd.n8720 5.896
R45608 vdd.n14071 vdd.n8553 5.896
R45609 vdd.n14130 vdd.n8499 5.896
R45610 vdd.n14359 vdd.n8335 5.896
R45611 vdd.n8284 vdd.n8242 5.896
R45612 vdd.n8088 vdd.n8070 5.896
R45613 vdd.n14803 vdd.n8063 5.896
R45614 vdd.n13134 vdd.n9238 5.896
R45615 vdd.n9088 vdd.n9077 5.896
R45616 vdd.n9031 vdd.n9015 5.896
R45617 vdd.n8868 vdd.n8857 5.896
R45618 vdd.n8811 vdd.n8795 5.896
R45619 vdd.n13944 vdd.n8630 5.896
R45620 vdd.n14020 vdd.n8582 5.896
R45621 vdd.n14234 vdd.n8409 5.896
R45622 vdd.n14309 vdd.n8363 5.896
R45623 vdd.n14550 vdd.n14539 5.896
R45624 vdd.n19394 vdd.n19393 5.896
R45625 vdd.n19443 vdd.n19442 5.896
R45626 vdd.n19600 vdd.n19599 5.896
R45627 vdd.n19643 vdd.n19642 5.896
R45628 vdd.n19802 vdd.n19801 5.896
R45629 vdd.n19158 vdd.n19157 5.896
R45630 vdd.n20851 vdd.n20850 5.896
R45631 vdd.n20808 vdd.n20807 5.896
R45632 vdd.n20652 vdd.n20651 5.896
R45633 vdd.n20603 vdd.n20602 5.896
R45634 vdd.n21605 vdd.n21604 5.896
R45635 vdd.n21409 vdd.n21408 5.896
R45636 vdd.n21360 vdd.n21359 5.896
R45637 vdd.n21150 vdd.n21149 5.896
R45638 vdd.n21101 vdd.n21100 5.896
R45639 vdd.n19043 vdd.n19042 5.896
R45640 vdd.n18994 vdd.n18993 5.896
R45641 vdd.n18784 vdd.n18783 5.896
R45642 vdd.n18735 vdd.n18734 5.896
R45643 vdd.n18525 vdd.n18524 5.896
R45644 vdd.n20283 vdd.n20277 5.896
R45645 vdd.n20265 vdd.n20259 5.896
R45646 vdd.n25246 vdd.n25245 5.896
R45647 vdd.n30302 vdd.n30301 5.882
R45648 vdd.n22174 vdd.n22173 5.88
R45649 vdd.n22195 vdd.n22194 5.88
R45650 vdd.n22053 vdd.n22052 5.88
R45651 vdd.n4885 vdd.n4884 5.869
R45652 vdd.n19367 vdd.n19366 5.864
R45653 vdd.n19480 vdd.n19479 5.864
R45654 vdd.n19573 vdd.n19572 5.864
R45655 vdd.n19680 vdd.n19679 5.864
R45656 vdd.n19775 vdd.n19774 5.864
R45657 vdd.n20972 vdd.n20971 5.864
R45658 vdd.n20877 vdd.n20876 5.864
R45659 vdd.n20781 vdd.n20780 5.864
R45660 vdd.n20689 vdd.n20688 5.864
R45661 vdd.n20576 vdd.n20575 5.864
R45662 vdd.n19978 vdd.n19977 5.864
R45663 vdd.n20313 vdd.n20312 5.864
R45664 vdd.n20231 vdd.n20228 5.864
R45665 vdd.n20077 vdd.n20076 5.864
R45666 vdd.n33679 vdd.n33678 5.862
R45667 vdd.n1144 vdd.n1143 5.862
R45668 vdd.n178 vdd.n177 5.855
R45669 vdd.n14760 vdd.n14759 5.849
R45670 vdd.n14818 vdd.n14817 5.849
R45671 vdd.n14931 vdd.n14930 5.849
R45672 vdd.n25432 vdd.n25431 5.834
R45673 vdd.n13391 vdd.t118 5.811
R45674 vdd.n8836 vdd.t327 5.811
R45675 vdd.t286 vdd.n8599 5.811
R45676 vdd.n8174 vdd.n8173 5.811
R45677 vdd.n13501 vdd.n8984 5.803
R45678 vdd.n13541 vdd.n8942 5.803
R45679 vdd.n13781 vdd.n8769 5.803
R45680 vdd.n13826 vdd.n8726 5.803
R45681 vdd.n14076 vdd.n8555 5.803
R45682 vdd.n8519 vdd.n8505 5.803
R45683 vdd.n13073 vdd.n13072 5.777
R45684 vdd.n13000 vdd.t294 5.777
R45685 vdd.n12962 vdd.n9466 5.777
R45686 vdd.n12865 vdd.n12864 5.777
R45687 vdd.n12754 vdd.n9826 5.777
R45688 vdd.n12709 vdd.t303 5.777
R45689 vdd.n9923 vdd.t303 5.777
R45690 vdd.n12657 vdd.n12656 5.777
R45691 vdd.n10155 vdd.t372 5.777
R45692 vdd.n12566 vdd.t381 5.777
R45693 vdd.n11047 vdd.t309 5.777
R45694 vdd.t266 vdd.n15657 5.777
R45695 vdd.n16374 vdd.t260 5.777
R45696 vdd.n16564 vdd.t14 5.777
R45697 vdd.n15115 vdd.t0 5.777
R45698 vdd.n17685 vdd.t271 5.777
R45699 vdd.n24714 vdd.n24713 5.715
R45700 vdd.n25197 vdd.n25196 5.715
R45701 vdd.n24713 vdd.n24712 5.715
R45702 vdd.n25196 vdd.n25195 5.715
R45703 vdd.n25534 vdd.n25533 5.697
R45704 vdd.n30302 vdd.n30300 5.693
R45705 vdd.n10165 vdd.n10146 5.688
R45706 vdd.n12624 vdd.n10050 5.688
R45707 vdd.n16761 vdd.n16760 5.688
R45708 vdd.n10264 vdd.n10261 5.655
R45709 vdd.n15065 vdd.n15064 5.655
R45710 vdd.n24199 vdd.n24198 5.654
R45711 vdd.n23977 vdd.n23976 5.654
R45712 vdd.n23967 vdd.n23966 5.654
R45713 vdd.n23745 vdd.n23744 5.654
R45714 vdd.n23735 vdd.n23734 5.654
R45715 vdd.n23057 vdd.n23056 5.654
R45716 vdd.n23279 vdd.n23278 5.654
R45717 vdd.n23289 vdd.n23288 5.654
R45718 vdd.n23511 vdd.n23510 5.654
R45719 vdd.n23521 vdd.n23520 5.654
R45720 vdd.n22478 vdd.n22477 5.654
R45721 vdd.n22700 vdd.n22699 5.654
R45722 vdd.n22710 vdd.n22709 5.654
R45723 vdd.n22932 vdd.n22931 5.654
R45724 vdd.n22942 vdd.n22941 5.654
R45725 vdd.n22182 vdd.n22181 5.654
R45726 vdd.n22265 vdd.n22264 5.654
R45727 vdd.n22276 vdd.n22275 5.654
R45728 vdd.n22150 vdd.n22149 5.654
R45729 vdd.n22161 vdd.n22160 5.654
R45730 vdd.n31542 vdd.n31541 5.647
R45731 vdd.n31551 vdd.n31550 5.647
R45732 vdd.n31030 vdd.n31029 5.647
R45733 vdd.n31284 vdd.n31283 5.647
R45734 vdd.n36025 vdd.n36024 5.647
R45735 vdd.n36039 vdd.n36038 5.647
R45736 vdd.n36256 vdd.n36255 5.647
R45737 vdd.n36270 vdd.n36269 5.647
R45738 vdd.n36487 vdd.n36486 5.647
R45739 vdd.n36501 vdd.n36500 5.647
R45740 vdd.n36718 vdd.n36717 5.647
R45741 vdd.n36732 vdd.n36731 5.647
R45742 vdd.n36949 vdd.n36948 5.647
R45743 vdd.n36963 vdd.n36962 5.647
R45744 vdd.n33141 vdd.n33140 5.647
R45745 vdd.n35635 vdd.n35634 5.647
R45746 vdd.n37317 vdd.n37316 5.647
R45747 vdd.n37347 vdd.n37346 5.647
R45748 vdd.n35662 vdd.n35661 5.647
R45749 vdd.n32824 vdd.n32823 5.647
R45750 vdd.n38018 vdd.n38017 5.647
R45751 vdd.n38004 vdd.n38003 5.647
R45752 vdd.n37787 vdd.n37786 5.647
R45753 vdd.n37773 vdd.n37772 5.647
R45754 vdd.n28215 vdd.n28214 5.647
R45755 vdd.n28229 vdd.n28228 5.647
R45756 vdd.n28446 vdd.n28445 5.647
R45757 vdd.n28460 vdd.n28459 5.647
R45758 vdd.n28677 vdd.n28676 5.647
R45759 vdd.n28691 vdd.n28690 5.647
R45760 vdd.n27987 vdd.n27977 5.647
R45761 vdd.n27979 vdd.n27978 5.647
R45762 vdd.n27875 vdd.n27874 5.647
R45763 vdd.n1655 vdd.n1654 5.647
R45764 vdd.n1645 vdd.n1644 5.647
R45765 vdd.n1474 vdd.n1473 5.647
R45766 vdd.n1464 vdd.n1463 5.647
R45767 vdd.n1293 vdd.n1292 5.647
R45768 vdd.n26759 vdd.n26758 5.647
R45769 vdd.n26930 vdd.n26929 5.647
R45770 vdd.n26940 vdd.n26939 5.647
R45771 vdd.n27111 vdd.n27110 5.647
R45772 vdd.n27121 vdd.n27120 5.647
R45773 vdd.n2066 vdd.n2065 5.647
R45774 vdd.n2124 vdd.n2123 5.647
R45775 vdd.n2139 vdd.n2138 5.647
R45776 vdd.n3727 vdd.n3726 5.647
R45777 vdd.n2689 vdd.n2688 5.647
R45778 vdd.n2883 vdd.n2882 5.647
R45779 vdd.n2893 vdd.n2892 5.647
R45780 vdd.n3064 vdd.n3063 5.647
R45781 vdd.n3074 vdd.n3073 5.647
R45782 vdd.n3245 vdd.n3244 5.647
R45783 vdd.n3255 vdd.n3254 5.647
R45784 vdd.n3426 vdd.n3425 5.647
R45785 vdd.n3436 vdd.n3435 5.647
R45786 vdd.n3607 vdd.n3606 5.647
R45787 vdd.n3617 vdd.n3616 5.647
R45788 vdd.n31682 vdd.n31681 5.647
R45789 vdd.n31683 vdd.n31682 5.647
R45790 vdd.n13357 vdd.n9064 5.647
R45791 vdd.n13402 vdd.n9049 5.647
R45792 vdd.n13649 vdd.n8844 5.647
R45793 vdd.n13695 vdd.n8828 5.647
R45794 vdd.n13965 vdd.n13964 5.647
R45795 vdd.n8626 vdd.n8625 5.647
R45796 vdd.n14255 vdd.n14254 5.647
R45797 vdd.n8404 vdd.n8403 5.647
R45798 vdd.n14682 vdd.n14681 5.647
R45799 vdd.n14710 vdd.n8111 5.647
R45800 vdd.n14855 vdd.n14853 5.647
R45801 vdd.n14904 vdd.n8024 5.647
R45802 vdd.n9199 vdd.n9182 5.647
R45803 vdd.n13243 vdd.n13241 5.647
R45804 vdd.n13278 vdd.n9155 5.647
R45805 vdd.n13283 vdd.n9153 5.647
R45806 vdd.n8977 vdd.n8961 5.647
R45807 vdd.n13535 vdd.n13533 5.647
R45808 vdd.n13570 vdd.n8934 5.647
R45809 vdd.n13575 vdd.n8932 5.647
R45810 vdd.n13816 vdd.n8741 5.647
R45811 vdd.n13818 vdd.n8715 5.647
R45812 vdd.n13858 vdd.n8716 5.647
R45813 vdd.n13874 vdd.n8705 5.647
R45814 vdd.n14103 vdd.n8528 5.647
R45815 vdd.n14104 vdd.n8493 5.647
R45816 vdd.n14147 vdd.n8494 5.647
R45817 vdd.n14163 vdd.n8482 5.647
R45818 vdd.n14389 vdd.n8293 5.647
R45819 vdd.n8294 vdd.n8290 5.647
R45820 vdd.n14413 vdd.n8291 5.647
R45821 vdd.n14443 vdd.n8267 5.647
R45822 vdd.n11737 vdd.n11726 5.647
R45823 vdd.n11737 vdd.n11736 5.647
R45824 vdd.n11697 vdd.n11687 5.647
R45825 vdd.n11709 vdd.n11708 5.647
R45826 vdd.n11821 vdd.n11815 5.647
R45827 vdd.n11830 vdd.n11815 5.647
R45828 vdd.n11860 vdd.n11859 5.647
R45829 vdd.n11852 vdd.n11841 5.647
R45830 vdd.n22173 vdd.n22166 5.647
R45831 vdd.n24103 vdd.n24096 5.647
R45832 vdd.n24077 vdd.n24070 5.647
R45833 vdd.n23871 vdd.n23864 5.647
R45834 vdd.n23845 vdd.n23838 5.647
R45835 vdd.n23639 vdd.n23632 5.647
R45836 vdd.n23157 vdd.n23150 5.647
R45837 vdd.n23183 vdd.n23176 5.647
R45838 vdd.n23389 vdd.n23382 5.647
R45839 vdd.n23415 vdd.n23408 5.647
R45840 vdd.n23621 vdd.n23614 5.647
R45841 vdd.n22578 vdd.n22571 5.647
R45842 vdd.n22604 vdd.n22597 5.647
R45843 vdd.n22810 vdd.n22803 5.647
R45844 vdd.n22836 vdd.n22829 5.647
R45845 vdd.n23042 vdd.n23035 5.647
R45846 vdd.n22194 vdd.n22187 5.647
R45847 vdd.n22052 vdd.n22045 5.647
R45848 vdd.n19260 vdd.n19259 5.647
R45849 vdd.n19248 vdd.n19247 5.647
R45850 vdd.n19204 vdd.n19203 5.647
R45851 vdd.n19192 vdd.n19191 5.647
R45852 vdd.n19846 vdd.n19845 5.647
R45853 vdd.n19858 vdd.n19857 5.647
R45854 vdd.n19914 vdd.n19913 5.647
R45855 vdd.n19926 vdd.n19925 5.647
R45856 vdd.n21521 vdd.n21520 5.647
R45857 vdd.n21503 vdd.n21502 5.647
R45858 vdd.n21262 vdd.n21261 5.647
R45859 vdd.n21244 vdd.n21243 5.647
R45860 vdd.n18896 vdd.n18895 5.647
R45861 vdd.n18878 vdd.n18877 5.647
R45862 vdd.n18637 vdd.n18636 5.647
R45863 vdd.n18619 vdd.n18618 5.647
R45864 vdd.n20406 vdd.n20394 5.647
R45865 vdd.n20383 vdd.n20371 5.647
R45866 vdd.n20170 vdd.n20158 5.647
R45867 vdd.n20147 vdd.n20135 5.647
R45868 vdd.n21819 vdd.n21814 5.647
R45869 vdd.n21912 vdd.n21906 5.647
R45870 vdd.n21921 vdd.n21906 5.647
R45871 vdd.n21951 vdd.n21950 5.647
R45872 vdd.n21943 vdd.n21932 5.647
R45873 vdd.n24743 vdd.n24736 5.647
R45874 vdd.n24757 vdd.n24752 5.647
R45875 vdd.n25175 vdd.n25168 5.647
R45876 vdd.n25159 vdd.n25154 5.647
R45877 vdd.n33288 vdd.n33287 5.643
R45878 vdd.n598 vdd.n597 5.643
R45879 vdd.n506 vdd.n505 5.643
R45880 vdd.n21576 vdd.n21575 5.629
R45881 vdd.n21458 vdd.t282 5.629
R45882 vdd.n21462 vdd.n21461 5.629
R45883 vdd.n21317 vdd.n21316 5.629
R45884 vdd.n21203 vdd.n21202 5.629
R45885 vdd.n21058 vdd.n21057 5.629
R45886 vdd.n19096 vdd.n19095 5.629
R45887 vdd.n18951 vdd.n18950 5.629
R45888 vdd.n18837 vdd.n18836 5.629
R45889 vdd.n18692 vdd.n18691 5.629
R45890 vdd.n18688 vdd.t350 5.629
R45891 vdd.n18578 vdd.n18577 5.629
R45892 vdd.n13344 vdd.n9098 5.591
R45893 vdd.n13395 vdd.n13394 5.591
R45894 vdd.n13636 vdd.n8878 5.591
R45895 vdd.n13687 vdd.n13686 5.591
R45896 vdd.n13912 vdd.n13911 5.591
R45897 vdd.n8607 vdd.n8604 5.591
R45898 vdd.n14202 vdd.n14201 5.591
R45899 vdd.n8385 vdd.n8382 5.591
R45900 vdd.n33668 vdd.n33667 5.506
R45901 vdd.n1061 vdd.n1060 5.506
R45902 vdd.t134 vdd.n13646 5.505
R45903 vdd.t315 vdd.n8399 5.505
R45904 vdd.n25381 vdd.n25380 5.484
R45905 vdd.n34102 vdd.n34101 5.461
R45906 vdd.n35481 vdd.n35480 5.461
R45907 vdd.n34960 vdd.n34959 5.461
R45908 vdd.n5810 vdd.n5809 5.461
R45909 vdd.n5707 vdd.n5706 5.461
R45910 vdd.n4534 vdd.n4533 5.461
R45911 vdd.n27383 vdd.n27382 5.461
R45912 vdd.n25826 vdd.n25825 5.461
R45913 vdd.n13024 vdd.n13023 5.456
R45914 vdd.n9561 vdd.n9556 5.456
R45915 vdd.n12816 vdd.n12815 5.456
R45916 vdd.n9923 vdd.n9922 5.456
R45917 vdd.n9938 vdd.t353 5.456
R45918 vdd.n12607 vdd.n12606 5.456
R45919 vdd.n10598 vdd.n10597 5.456
R45920 vdd.n10757 vdd.n10749 5.456
R45921 vdd.n12286 vdd.n12285 5.456
R45922 vdd.n12179 vdd.n11096 5.456
R45923 vdd.n12074 vdd.n12073 5.456
R45924 vdd.n11980 vdd.n11979 5.456
R45925 vdd.n11526 vdd.t374 5.456
R45926 vdd.n11599 vdd.n11564 5.456
R45927 vdd.n15609 vdd.n15606 5.456
R45928 vdd.n15865 vdd.n15862 5.456
R45929 vdd.n16121 vdd.n16118 5.456
R45930 vdd.n16377 vdd.n16374 5.456
R45931 vdd.n16394 vdd.t16 5.456
R45932 vdd.n16616 vdd.n16614 5.456
R45933 vdd.n16976 vdd.n16973 5.456
R45934 vdd.n17248 vdd.n17245 5.456
R45935 vdd.n17520 vdd.n17517 5.456
R45936 vdd.n17778 vdd.n17775 5.456
R45937 vdd.n18049 vdd.n18046 5.456
R45938 vdd.n16815 vdd.n16813 5.456
R45939 vdd.n18363 vdd.t23 5.456
R45940 vdd.n21704 vdd.n15016 5.456
R45941 vdd.n24827 vdd.n24826 5.449
R45942 vdd.n25025 vdd.n25024 5.418
R45943 vdd.n24599 vdd.n24598 5.418
R45944 vdd.n25386 vdd.n25385 5.395
R45945 vdd.n28092 vdd.n28091 5.375
R45946 vdd.n22238 vdd.n22237 5.343
R45947 vdd.n22114 vdd.n22113 5.343
R45948 vdd.n33988 vdd.n33987 5.335
R45949 vdd.n35150 vdd.n35149 5.335
R45950 vdd.n34565 vdd.n34564 5.335
R45951 vdd.n6276 vdd.n6275 5.335
R45952 vdd.n5312 vdd.n5311 5.335
R45953 vdd.n5145 vdd.n5144 5.335
R45954 vdd.n4143 vdd.n4142 5.335
R45955 vdd.n27615 vdd.n27614 5.335
R45956 vdd.n26036 vdd.n26035 5.335
R45957 vdd.n33344 vdd.n33343 5.327
R45958 vdd.n610 vdd.n609 5.327
R45959 vdd.n515 vdd.n514 5.327
R45960 vdd.n33397 vdd.n33396 5.32
R45961 vdd.n716 vdd.n715 5.32
R45962 vdd.n447 vdd.n446 5.32
R45963 vdd.n33895 vdd.n33894 5.313
R45964 vdd.n35089 vdd.n35088 5.313
R45965 vdd.n34502 vdd.n34501 5.313
R45966 vdd.n6169 vdd.n6168 5.313
R45967 vdd.n5249 vdd.n5248 5.313
R45968 vdd.n4977 vdd.n4976 5.313
R45969 vdd.n4079 vdd.n4078 5.313
R45970 vdd.n27552 vdd.n27551 5.313
R45971 vdd.n25989 vdd.n25988 5.313
R45972 vdd.n34373 vdd.n34372 5.305
R45973 vdd.n35396 vdd.n35395 5.305
R45974 vdd.n34799 vdd.n34798 5.305
R45975 vdd.n6087 vdd.n6086 5.305
R45976 vdd.n5546 vdd.n5545 5.305
R45977 vdd.n4762 vdd.n4761 5.305
R45978 vdd.n4373 vdd.n4372 5.305
R45979 vdd.n27267 vdd.n27266 5.305
R45980 vdd.n25922 vdd.n25921 5.305
R45981 vdd.n25424 vdd.n25423 5.279
R45982 vdd.n19350 vdd.n19347 5.277
R45983 vdd.n19495 vdd.n19492 5.277
R45984 vdd.n19556 vdd.n19553 5.277
R45985 vdd.t164 vdd.n19588 5.277
R45986 vdd.n19695 vdd.n19692 5.277
R45987 vdd.n19758 vdd.n19755 5.277
R45988 vdd.n20955 vdd.n20952 5.277
R45989 vdd.n20892 vdd.n20889 5.277
R45990 vdd.t174 vdd.n20796 5.277
R45991 vdd.n20765 vdd.n20762 5.277
R45992 vdd.n20704 vdd.n20701 5.277
R45993 vdd.n20559 vdd.n20556 5.277
R45994 vdd.n20451 vdd.n20450 5.277
R45995 vdd.n20330 vdd.n20329 5.277
R45996 vdd.n20216 vdd.n20215 5.277
R45997 vdd.n20094 vdd.n20093 5.277
R45998 vdd.n33510 vdd.n33509 5.27
R45999 vdd.n1034 vdd.n1033 5.27
R46000 vdd.n31268 vdd.n31264 5.27
R46001 vdd.n30547 vdd.n30540 5.27
R46002 vdd.n35899 vdd.n35892 5.27
R46003 vdd.n35948 vdd.n35941 5.27
R46004 vdd.n36130 vdd.n36123 5.27
R46005 vdd.n36179 vdd.n36172 5.27
R46006 vdd.n36361 vdd.n36354 5.27
R46007 vdd.n36410 vdd.n36403 5.27
R46008 vdd.n36592 vdd.n36585 5.27
R46009 vdd.n36641 vdd.n36634 5.27
R46010 vdd.n36823 vdd.n36816 5.27
R46011 vdd.n36872 vdd.n36865 5.27
R46012 vdd.n37058 vdd.n37051 5.27
R46013 vdd.n37097 vdd.n37090 5.27
R46014 vdd.n37228 vdd.n37224 5.27
R46015 vdd.n33059 vdd.n33052 5.27
R46016 vdd.n32929 vdd.n32922 5.27
R46017 vdd.n37470 vdd.n37463 5.27
R46018 vdd.n38152 vdd.n38145 5.27
R46019 vdd.n38109 vdd.n38102 5.27
R46020 vdd.n37927 vdd.n37920 5.27
R46021 vdd.n37878 vdd.n37871 5.27
R46022 vdd.n37696 vdd.n37689 5.27
R46023 vdd.n37647 vdd.n37640 5.27
R46024 vdd.n28320 vdd.n28313 5.27
R46025 vdd.n28369 vdd.n28362 5.27
R46026 vdd.n28551 vdd.n28544 5.27
R46027 vdd.n28600 vdd.n28593 5.27
R46028 vdd.n28782 vdd.n28775 5.27
R46029 vdd.n28165 vdd.n28158 5.27
R46030 vdd.n29872 vdd.n29865 5.27
R46031 vdd.n29838 vdd.n29831 5.27
R46032 vdd.n1758 vdd.n1754 5.27
R46033 vdd.n1725 vdd.n1721 5.27
R46034 vdd.n1583 vdd.n1579 5.27
R46035 vdd.n1544 vdd.n1540 5.27
R46036 vdd.n1402 vdd.n1398 5.27
R46037 vdd.n1363 vdd.n1359 5.27
R46038 vdd.n26829 vdd.n26825 5.27
R46039 vdd.n26868 vdd.n26864 5.27
R46040 vdd.n27010 vdd.n27006 5.27
R46041 vdd.n27049 vdd.n27045 5.27
R46042 vdd.n27191 vdd.n27187 5.27
R46043 vdd.n26737 vdd.n26733 5.27
R46044 vdd.n2067 vdd.n2066 5.27
R46045 vdd.n2782 vdd.n2778 5.27
R46046 vdd.n2821 vdd.n2817 5.27
R46047 vdd.n2963 vdd.n2959 5.27
R46048 vdd.n3002 vdd.n2998 5.27
R46049 vdd.n3144 vdd.n3140 5.27
R46050 vdd.n3183 vdd.n3179 5.27
R46051 vdd.n3325 vdd.n3321 5.27
R46052 vdd.n3364 vdd.n3360 5.27
R46053 vdd.n3506 vdd.n3502 5.27
R46054 vdd.n3545 vdd.n3541 5.27
R46055 vdd.n13207 vdd.n9206 5.27
R46056 vdd.n13208 vdd.n13207 5.27
R46057 vdd.n13249 vdd.n9163 5.27
R46058 vdd.n13268 vdd.n9163 5.27
R46059 vdd.n13501 vdd.n8986 5.27
R46060 vdd.n13560 vdd.n8942 5.27
R46061 vdd.n13781 vdd.n13780 5.27
R46062 vdd.n13842 vdd.n8726 5.27
R46063 vdd.n14076 vdd.n8554 5.27
R46064 vdd.n14131 vdd.n8505 5.27
R46065 vdd.n14357 vdd.n14356 5.27
R46066 vdd.n14356 vdd.n8338 5.27
R46067 vdd.n14422 vdd.n8278 5.27
R46068 vdd.n14422 vdd.n8283 5.27
R46069 vdd.n14769 vdd.n8090 5.27
R46070 vdd.n14791 vdd.n8069 5.27
R46071 vdd.n14798 vdd.n8061 5.27
R46072 vdd.n14806 vdd.n14805 5.27
R46073 vdd.n9086 vdd.n9085 5.27
R46074 vdd.n9085 vdd.n9080 5.27
R46075 vdd.n13430 vdd.n9025 5.27
R46076 vdd.n13430 vdd.n9030 5.27
R46077 vdd.n8866 vdd.n8865 5.27
R46078 vdd.n8865 vdd.n8860 5.27
R46079 vdd.n13722 vdd.n8805 5.27
R46080 vdd.n13722 vdd.n8810 5.27
R46081 vdd.n13958 vdd.n8634 5.27
R46082 vdd.n13958 vdd.n8635 5.27
R46083 vdd.n14014 vdd.n8586 5.27
R46084 vdd.n14014 vdd.n8583 5.27
R46085 vdd.n14248 vdd.n8412 5.27
R46086 vdd.n14248 vdd.n8413 5.27
R46087 vdd.n14304 vdd.n8366 5.27
R46088 vdd.n14304 vdd.n8364 5.27
R46089 vdd.n14545 vdd.n14538 5.27
R46090 vdd.n14545 vdd.n14544 5.27
R46091 vdd.n24285 vdd.n24284 5.27
R46092 vdd.n24180 vdd.n24179 5.27
R46093 vdd.n23986 vdd.n23985 5.27
R46094 vdd.n23948 vdd.n23947 5.27
R46095 vdd.n23754 vdd.n23753 5.27
R46096 vdd.n23716 vdd.n23715 5.27
R46097 vdd.n23066 vdd.n23065 5.27
R46098 vdd.n23260 vdd.n23259 5.27
R46099 vdd.n23298 vdd.n23297 5.27
R46100 vdd.n23492 vdd.n23491 5.27
R46101 vdd.n23530 vdd.n23529 5.27
R46102 vdd.n22487 vdd.n22486 5.27
R46103 vdd.n22681 vdd.n22680 5.27
R46104 vdd.n22719 vdd.n22718 5.27
R46105 vdd.n22913 vdd.n22912 5.27
R46106 vdd.n22951 vdd.n22950 5.27
R46107 vdd.n22457 vdd.n22456 5.27
R46108 vdd.n22313 vdd.n22312 5.27
R46109 vdd.n19401 vdd.n19392 5.27
R46110 vdd.n19450 vdd.n19441 5.27
R46111 vdd.n19607 vdd.n19598 5.27
R46112 vdd.n19650 vdd.n19641 5.27
R46113 vdd.n19809 vdd.n19800 5.27
R46114 vdd.n20997 vdd.n19160 5.27
R46115 vdd.n20858 vdd.n20849 5.27
R46116 vdd.n20815 vdd.n20806 5.27
R46117 vdd.n20659 vdd.n20650 5.27
R46118 vdd.n20610 vdd.n20601 5.27
R46119 vdd.n21416 vdd.n21407 5.27
R46120 vdd.n21367 vdd.n21358 5.27
R46121 vdd.n21157 vdd.n21148 5.27
R46122 vdd.n21108 vdd.n21099 5.27
R46123 vdd.n19050 vdd.n19041 5.27
R46124 vdd.n19001 vdd.n18992 5.27
R46125 vdd.n18791 vdd.n18782 5.27
R46126 vdd.n18742 vdd.n18733 5.27
R46127 vdd.n18532 vdd.n18523 5.27
R46128 vdd.n20275 vdd.n20274 5.27
R46129 vdd.n20257 vdd.n20256 5.27
R46130 vdd.n24824 vdd.n24823 5.27
R46131 vdd.n25242 vdd.n25241 5.27
R46132 vdd.n25566 vdd.n25565 5.266
R46133 vdd.n14672 vdd.n8134 5.264
R46134 vdd.n14748 vdd.n8100 5.264
R46135 vdd.n14834 vdd.n8044 5.264
R46136 vdd.n14926 vdd.n8009 5.264
R46137 vdd.t118 vdd.n9020 5.199
R46138 vdd.n8601 vdd.t286 5.199
R46139 vdd.n10387 vdd.n10339 5.135
R46140 vdd.n10381 vdd.n10380 5.135
R46141 vdd.n13081 vdd.n13080 5.135
R46142 vdd.n12993 vdd.n9415 5.135
R46143 vdd.n9464 vdd.n9455 5.135
R46144 vdd.n12888 vdd.n12887 5.135
R46145 vdd.n12881 vdd.n9614 5.135
R46146 vdd.n12873 vdd.n12872 5.135
R46147 vdd.n9798 vdd.n9775 5.135
R46148 vdd.n12785 vdd.n9776 5.135
R46149 vdd.n9824 vdd.n9815 5.135
R46150 vdd.n12680 vdd.n12679 5.135
R46151 vdd.n12673 vdd.n9974 5.135
R46152 vdd.n12665 vdd.n12664 5.135
R46153 vdd.n10241 vdd.n10118 5.135
R46154 vdd.n12587 vdd.n10119 5.135
R46155 vdd.n12432 vdd.n10665 5.135
R46156 vdd.n10689 vdd.n10688 5.135
R46157 vdd.n10845 vdd.n10824 5.135
R46158 vdd.n10860 vdd.n10825 5.135
R46159 vdd.n12240 vdd.n11004 5.135
R46160 vdd.n12234 vdd.n11011 5.135
R46161 vdd.n12133 vdd.n12132 5.135
R46162 vdd.n12122 vdd.n12121 5.135
R46163 vdd.n11354 vdd.n11333 5.135
R46164 vdd.n11369 vdd.n11334 5.135
R46165 vdd.n15251 vdd.n15250 5.135
R46166 vdd.n15240 vdd.n15239 5.135
R46167 vdd.n15456 vdd.n15455 5.135
R46168 vdd.n15215 vdd.n15214 5.135
R46169 vdd.n15712 vdd.n15711 5.135
R46170 vdd.n15201 vdd.n15200 5.135
R46171 vdd.n15196 vdd.n15195 5.135
R46172 vdd.n15968 vdd.n15967 5.135
R46173 vdd.n15173 vdd.n15172 5.135
R46174 vdd.n15159 vdd.n15158 5.135
R46175 vdd.n16224 vdd.n16223 5.135
R46176 vdd.n15145 vdd.n15144 5.135
R46177 vdd.n15131 vdd.n15130 5.135
R46178 vdd.n16480 vdd.n16479 5.135
R46179 vdd.n16663 vdd.n16662 5.135
R46180 vdd.n16658 vdd.n16657 5.135
R46181 vdd.n17103 vdd.n17102 5.135
R46182 vdd.n17123 vdd.n17122 5.135
R46183 vdd.n17375 vdd.n17374 5.135
R46184 vdd.n17395 vdd.n17394 5.135
R46185 vdd.n17633 vdd.n17632 5.135
R46186 vdd.n17653 vdd.n17652 5.135
R46187 vdd.n17904 vdd.n17903 5.135
R46188 vdd.n17924 vdd.n17923 5.135
R46189 vdd.n18176 vdd.n18175 5.135
R46190 vdd.n18196 vdd.n18195 5.135
R46191 vdd.n11628 vdd.n9276 5.117
R46192 vdd.n13110 vdd.n9276 5.117
R46193 vdd.n13145 vdd.n9244 5.117
R46194 vdd.n13217 vdd.n13216 5.117
R46195 vdd.n33464 vdd.n33463 5.081
R46196 vdd.n783 vdd.n782 5.081
R46197 vdd.n478 vdd.n477 5.081
R46198 vdd.n33877 vdd.n33876 5.081
R46199 vdd.n35102 vdd.n35101 5.081
R46200 vdd.n34515 vdd.n34514 5.081
R46201 vdd.n6151 vdd.n6150 5.081
R46202 vdd.n5262 vdd.n5261 5.081
R46203 vdd.n4960 vdd.n4959 5.081
R46204 vdd.n4092 vdd.n4091 5.081
R46205 vdd.n27572 vdd.n27571 5.081
R46206 vdd.n25685 vdd.n25684 5.081
R46207 vdd.n29033 vdd.n29032 5.079
R46208 vdd.n12570 vdd.n10257 4.991
R46209 vdd.n15120 vdd.n15119 4.991
R46210 vdd.n10169 vdd.n10146 4.977
R46211 vdd.n16767 vdd.n16765 4.977
R46212 vdd.n25583 vdd.n25582 4.951
R46213 vdd.n21591 vdd.n21588 4.925
R46214 vdd.n21445 vdd.n21442 4.925
R46215 vdd.n21332 vdd.n21329 4.925
R46216 vdd.n21186 vdd.n21183 4.925
R46217 vdd.n21073 vdd.n21070 4.925
R46218 vdd.n21025 vdd.t280 4.925
R46219 vdd.n19126 vdd.t347 4.925
R46220 vdd.n19079 vdd.n19076 4.925
R46221 vdd.n18966 vdd.n18963 4.925
R46222 vdd.n18820 vdd.n18817 4.925
R46223 vdd.n18707 vdd.n18704 4.925
R46224 vdd.n18561 vdd.n18558 4.925
R46225 vdd.n36011 vdd.n36010 4.894
R46226 vdd.n36053 vdd.n36052 4.894
R46227 vdd.n36242 vdd.n36241 4.894
R46228 vdd.n36284 vdd.n36283 4.894
R46229 vdd.n36473 vdd.n36472 4.894
R46230 vdd.n36515 vdd.n36514 4.894
R46231 vdd.n36704 vdd.n36703 4.894
R46232 vdd.n36746 vdd.n36745 4.894
R46233 vdd.n36935 vdd.n36934 4.894
R46234 vdd.n35682 vdd.n35681 4.894
R46235 vdd.n37143 vdd.n37142 4.894
R46236 vdd.n37171 vdd.n37170 4.894
R46237 vdd.n32984 vdd.n32983 4.894
R46238 vdd.n32970 vdd.n32969 4.894
R46239 vdd.n37518 vdd.n37517 4.894
R46240 vdd.n37564 vdd.n37563 4.894
R46241 vdd.n38032 vdd.n38031 4.894
R46242 vdd.n37990 vdd.n37989 4.894
R46243 vdd.n37801 vdd.n37800 4.894
R46244 vdd.n37759 vdd.n37758 4.894
R46245 vdd.n28201 vdd.n28200 4.894
R46246 vdd.n28243 vdd.n28242 4.894
R46247 vdd.n28432 vdd.n28431 4.894
R46248 vdd.n28474 vdd.n28473 4.894
R46249 vdd.n28663 vdd.n28662 4.894
R46250 vdd.n28705 vdd.n28704 4.894
R46251 vdd.n28117 vdd.n28116 4.894
R46252 vdd.n28082 vdd.n28081 4.894
R46253 vdd.n29716 vdd.n29715 4.894
R46254 vdd.n1666 vdd.n1665 4.894
R46255 vdd.n1634 vdd.n1633 4.894
R46256 vdd.n1485 vdd.n1484 4.894
R46257 vdd.n1453 vdd.n1452 4.894
R46258 vdd.n1304 vdd.n1303 4.894
R46259 vdd.n26770 vdd.n26769 4.894
R46260 vdd.n26919 vdd.n26918 4.894
R46261 vdd.n26951 vdd.n26950 4.894
R46262 vdd.n27100 vdd.n27099 4.894
R46263 vdd.n27132 vdd.n27131 4.894
R46264 vdd.n2872 vdd.n2871 4.894
R46265 vdd.n2904 vdd.n2903 4.894
R46266 vdd.n3053 vdd.n3052 4.894
R46267 vdd.n3085 vdd.n3084 4.894
R46268 vdd.n3234 vdd.n3233 4.894
R46269 vdd.n3266 vdd.n3265 4.894
R46270 vdd.n3415 vdd.n3414 4.894
R46271 vdd.n3447 vdd.n3446 4.894
R46272 vdd.n3596 vdd.n3595 4.894
R46273 vdd.n3638 vdd.n3637 4.894
R46274 vdd.n13368 vdd.n9067 4.894
R46275 vdd.n9052 vdd.n9051 4.894
R46276 vdd.n13660 vdd.n8847 4.894
R46277 vdd.n8832 vdd.n8830 4.894
R46278 vdd.n8666 vdd.n8660 4.894
R46279 vdd.n13980 vdd.n8611 4.894
R46280 vdd.n8443 vdd.n8440 4.894
R46281 vdd.n14270 vdd.n8389 4.894
R46282 vdd.n14693 vdd.n14692 4.894
R46283 vdd.n14692 vdd.n8129 4.894
R46284 vdd.n14718 vdd.n8108 4.894
R46285 vdd.n14739 vdd.n8108 4.894
R46286 vdd.n14867 vdd.n14866 4.894
R46287 vdd.n14866 vdd.n8039 4.894
R46288 vdd.n14898 vdd.n8025 4.894
R46289 vdd.n14898 vdd.n14884 4.894
R46290 vdd.n13225 vdd.n9195 4.894
R46291 vdd.n9201 vdd.n9200 4.894
R46292 vdd.n13284 vdd.n9137 4.894
R46293 vdd.n13308 vdd.n13307 4.894
R46294 vdd.n13517 vdd.n8973 4.894
R46295 vdd.n8979 vdd.n8978 4.894
R46296 vdd.n13576 vdd.n8915 4.894
R46297 vdd.n13600 vdd.n13599 4.894
R46298 vdd.n8761 vdd.n8743 4.894
R46299 vdd.n8746 vdd.n8744 4.894
R46300 vdd.n13873 vdd.n8703 4.894
R46301 vdd.n13882 vdd.n8701 4.894
R46302 vdd.n8548 vdd.n8530 4.894
R46303 vdd.n8532 vdd.n8531 4.894
R46304 vdd.n14162 vdd.n8480 4.894
R46305 vdd.n14171 vdd.n8478 4.894
R46306 vdd.n14385 vdd.n8307 4.894
R46307 vdd.n14388 vdd.n8308 4.894
R46308 vdd.n14442 vdd.n8264 4.894
R46309 vdd.n14445 vdd.n8265 4.894
R46310 vdd.n11690 vdd.n11685 4.894
R46311 vdd.n11704 vdd.n11691 4.894
R46312 vdd.n11820 vdd.n11817 4.894
R46313 vdd.n11865 vdd.n11864 4.894
R46314 vdd.n11847 vdd.n11846 4.894
R46315 vdd.n24219 vdd.n24212 4.894
R46316 vdd.n24117 vdd.n24110 4.894
R46317 vdd.n24063 vdd.n24056 4.894
R46318 vdd.n23885 vdd.n23878 4.894
R46319 vdd.n23831 vdd.n23824 4.894
R46320 vdd.n23653 vdd.n23646 4.894
R46321 vdd.n23143 vdd.n23136 4.894
R46322 vdd.n23197 vdd.n23190 4.894
R46323 vdd.n23375 vdd.n23368 4.894
R46324 vdd.n23429 vdd.n23422 4.894
R46325 vdd.n23607 vdd.n23600 4.894
R46326 vdd.n22564 vdd.n22557 4.894
R46327 vdd.n22618 vdd.n22611 4.894
R46328 vdd.n22796 vdd.n22789 4.894
R46329 vdd.n22850 vdd.n22843 4.894
R46330 vdd.n23028 vdd.n23021 4.894
R46331 vdd.n22391 vdd.n22384 4.894
R46332 vdd.n22361 vdd.n22352 4.894
R46333 vdd.n24336 vdd.n24329 4.894
R46334 vdd.n22090 vdd.n22081 4.894
R46335 vdd.n19272 vdd.n19271 4.894
R46336 vdd.n19236 vdd.n19235 4.894
R46337 vdd.n19216 vdd.n19215 4.894
R46338 vdd.n19179 vdd.n19178 4.894
R46339 vdd.n19833 vdd.n19832 4.894
R46340 vdd.n19870 vdd.n19869 4.894
R46341 vdd.n19902 vdd.n19901 4.894
R46342 vdd.n19938 vdd.n19937 4.894
R46343 vdd.n21537 vdd.n21536 4.894
R46344 vdd.n21487 vdd.n21486 4.894
R46345 vdd.n21278 vdd.n21277 4.894
R46346 vdd.n21228 vdd.n21227 4.894
R46347 vdd.n21021 vdd.n21020 4.894
R46348 vdd.n19121 vdd.n19120 4.894
R46349 vdd.n18912 vdd.n18911 4.894
R46350 vdd.n18862 vdd.n18861 4.894
R46351 vdd.n18653 vdd.n18652 4.894
R46352 vdd.n18603 vdd.n18602 4.894
R46353 vdd.n20422 vdd.n20413 4.894
R46354 vdd.n20364 vdd.n20355 4.894
R46355 vdd.n20186 vdd.n20177 4.894
R46356 vdd.n20128 vdd.n20119 4.894
R46357 vdd.n21911 vdd.n21908 4.894
R46358 vdd.n21956 vdd.n21955 4.894
R46359 vdd.n21938 vdd.n21937 4.894
R46360 vdd.n24729 vdd.n24724 4.894
R46361 vdd.n24769 vdd.n24764 4.894
R46362 vdd.n25187 vdd.n25182 4.894
R46363 vdd.n25147 vdd.n25142 4.894
R46364 vdd.n13438 vdd.n9020 4.893
R46365 vdd.n13510 vdd.n13509 4.893
R46366 vdd.n13730 vdd.n8800 4.893
R46367 vdd.n8766 vdd.n8749 4.893
R46368 vdd.n13935 vdd.t331 4.893
R46369 vdd.n13993 vdd.n8599 4.893
R46370 vdd.n14284 vdd.n8377 4.893
R46371 vdd.n14396 vdd.n14395 4.893
R46372 vdd.n14603 vdd.n14566 4.893
R46373 vdd.n14614 vdd.n8172 4.893
R46374 vdd.n32013 vdd.n31617 4.86
R46375 vdd.n26706 vdd.n26705 4.86
R46376 vdd.n10576 vdd.n10565 4.851
R46377 vdd.n12469 vdd.n10604 4.851
R46378 vdd.n12393 vdd.n10721 4.851
R46379 vdd.n10783 vdd.n10765 4.851
R46380 vdd.n12294 vdd.n10904 4.851
R46381 vdd.n12272 vdd.n10923 4.851
R46382 vdd.n12194 vdd.n11085 4.851
R46383 vdd.n12172 vdd.n11108 4.851
R46384 vdd.n11257 vdd.n11248 4.851
R46385 vdd.n11291 vdd.n11275 4.851
R46386 vdd.n11988 vdd.n11413 4.851
R46387 vdd.n11966 vdd.n11432 4.851
R46388 vdd.n10464 vdd.n10278 4.851
R46389 vdd.n10428 vdd.n10306 4.851
R46390 vdd.n9315 vdd.n9309 4.851
R46391 vdd.n9382 vdd.n9369 4.851
R46392 vdd.n12954 vdd.n9477 4.851
R46393 vdd.n9552 vdd.n9527 4.851
R46394 vdd.n9676 vdd.n9670 4.851
R46395 vdd.n9742 vdd.n9729 4.851
R46396 vdd.n12746 vdd.n9837 4.851
R46397 vdd.n9912 vdd.n9888 4.851
R46398 vdd.n10036 vdd.n10030 4.851
R46399 vdd.n10187 vdd.n10141 4.851
R46400 vdd.n16948 vdd.n16942 4.851
R46401 vdd.n17008 vdd.n17002 4.851
R46402 vdd.n17220 vdd.n17214 4.851
R46403 vdd.n17280 vdd.n17274 4.851
R46404 vdd.n17492 vdd.n17486 4.851
R46405 vdd.n17552 vdd.n17546 4.851
R46406 vdd.n17750 vdd.n17744 4.851
R46407 vdd.n17810 vdd.n17804 4.851
R46408 vdd.n18021 vdd.n18015 4.851
R46409 vdd.n18081 vdd.n18075 4.851
R46410 vdd.n18288 vdd.n18283 4.851
R46411 vdd.n18328 vdd.n18323 4.851
R46412 vdd.n15284 vdd.n15283 4.851
R46413 vdd.n15335 vdd.n15334 4.851
R46414 vdd.n15506 vdd.n15505 4.851
R46415 vdd.n15569 vdd.n15568 4.851
R46416 vdd.n15762 vdd.n15761 4.851
R46417 vdd.n15825 vdd.n15824 4.851
R46418 vdd.n16018 vdd.n16017 4.851
R46419 vdd.n16081 vdd.n16080 4.851
R46420 vdd.n16274 vdd.n16273 4.851
R46421 vdd.n16337 vdd.n16336 4.851
R46422 vdd.n16530 vdd.n16529 4.851
R46423 vdd.n16714 vdd.n16713 4.851
R46424 vdd.n10454 vdd.n10453 4.84
R46425 vdd.n10442 vdd.n10441 4.84
R46426 vdd.n15303 vdd.n15301 4.84
R46427 vdd.n15324 vdd.n15323 4.84
R46428 vdd.n9343 vdd.n9341 4.814
R46429 vdd.n13032 vdd.n9354 4.814
R46430 vdd.n9385 vdd.n9384 4.814
R46431 vdd.n12946 vdd.n9508 4.814
R46432 vdd.n9541 vdd.n9539 4.814
R46433 vdd.n12842 vdd.t355 4.814
R46434 vdd.n9703 vdd.n9701 4.814
R46435 vdd.n12824 vdd.n9714 4.814
R46436 vdd.n9745 vdd.n9744 4.814
R46437 vdd.n12738 vdd.n9868 4.814
R46438 vdd.n9901 vdd.n9900 4.814
R46439 vdd.n12711 vdd.n9915 4.814
R46440 vdd.n10157 vdd.n10154 4.814
R46441 vdd.n12615 vdd.n10056 4.814
R46442 vdd.n10190 vdd.n10189 4.814
R46443 vdd.n12488 vdd.n10574 4.814
R46444 vdd.n12482 vdd.n10583 4.814
R46445 vdd.n12383 vdd.n12382 4.814
R46446 vdd.n10763 vdd.n10762 4.814
R46447 vdd.t379 vdd.n12342 4.814
R46448 vdd.n10938 vdd.n10915 4.814
R46449 vdd.n12279 vdd.n10917 4.814
R46450 vdd.n11099 vdd.n11095 4.814
R46451 vdd.n11118 vdd.n11117 4.814
R46452 vdd.n12084 vdd.n11241 4.814
R46453 vdd.n11482 vdd.n11424 4.814
R46454 vdd.n11973 vdd.n11426 4.814
R46455 vdd.n15531 vdd.n15526 4.814
R46456 vdd.n15558 vdd.n15557 4.814
R46457 vdd.n15592 vdd.n15589 4.814
R46458 vdd.n15787 vdd.n15782 4.814
R46459 vdd.n15814 vdd.n15813 4.814
R46460 vdd.n16024 vdd.t18 4.814
R46461 vdd.n16043 vdd.n16038 4.814
R46462 vdd.n16070 vdd.n16069 4.814
R46463 vdd.n16104 vdd.n16101 4.814
R46464 vdd.n16299 vdd.n16294 4.814
R46465 vdd.n16326 vdd.n16325 4.814
R46466 vdd.n16360 vdd.n16357 4.814
R46467 vdd.n16571 vdd.n16548 4.814
R46468 vdd.n16558 vdd.n16556 4.814
R46469 vdd.n16610 vdd.n16609 4.814
R46470 vdd.n16962 vdd.n16959 4.814
R46471 vdd.n16990 vdd.n16987 4.814
R46472 vdd.n17234 vdd.n17231 4.814
R46473 vdd.n17262 vdd.n17259 4.814
R46474 vdd.n17355 vdd.t25 4.814
R46475 vdd.n17506 vdd.n17503 4.814
R46476 vdd.n17534 vdd.n17531 4.814
R46477 vdd.n17764 vdd.n17761 4.814
R46478 vdd.n17792 vdd.n17789 4.814
R46479 vdd.n18035 vdd.n18032 4.814
R46480 vdd.n18301 vdd.n18299 4.814
R46481 vdd.n15033 vdd.n15031 4.814
R46482 vdd.n24908 vdd.n24893 4.812
R46483 vdd.n24529 vdd.n24526 4.811
R46484 vdd.n35848 vdd.n35706 4.804
R46485 vdd.n1820 vdd.n1819 4.802
R46486 vdd.n24554 vdd.n24535 4.79
R46487 vdd.n2743 vdd.n2735 4.772
R46488 vdd.n24932 vdd.n24912 4.767
R46489 vdd.n167 vdd.n166 4.753
R46490 vdd.n34319 vdd.n34318 4.746
R46491 vdd.n35585 vdd.n35584 4.746
R46492 vdd.n34891 vdd.n34890 4.746
R46493 vdd.n5934 vdd.n5933 4.746
R46494 vdd.n5638 vdd.n5637 4.746
R46495 vdd.n4625 vdd.n4624 4.746
R46496 vdd.n4465 vdd.n4464 4.746
R46497 vdd.n27451 vdd.n27450 4.746
R46498 vdd.n25897 vdd.n25896 4.746
R46499 vdd.n12618 vdd.n12617 4.74
R46500 vdd.n16751 vdd.n16750 4.74
R46501 vdd.n31149 vdd.n31141 4.739
R46502 vdd.n33979 vdd.n33978 4.738
R46503 vdd.n35141 vdd.n35140 4.738
R46504 vdd.n34554 vdd.n34553 4.738
R46505 vdd.n6264 vdd.n6263 4.738
R46506 vdd.n5301 vdd.n5300 4.738
R46507 vdd.n5158 vdd.n5157 4.738
R46508 vdd.n4131 vdd.n4130 4.738
R46509 vdd.n27257 vdd.n27256 4.738
R46510 vdd.n26025 vdd.n26024 4.738
R46511 vdd.n33355 vdd.n33354 4.731
R46512 vdd.n673 vdd.n672 4.731
R46513 vdd.n565 vdd.n564 4.731
R46514 vdd.n24976 vdd.n24975 4.723
R46515 vdd.n25054 vdd.n25053 4.723
R46516 vdd.n24635 vdd.n24634 4.723
R46517 vdd.n24994 vdd.n24993 4.722
R46518 vdd.n24570 vdd.n24569 4.722
R46519 vdd.n30507 vdd.n30332 4.707
R46520 vdd.n34356 vdd.n34355 4.704
R46521 vdd.n35372 vdd.n35371 4.704
R46522 vdd.n34782 vdd.n34781 4.704
R46523 vdd.n6062 vdd.n6061 4.704
R46524 vdd.n5529 vdd.n5528 4.704
R46525 vdd.n4775 vdd.n4774 4.704
R46526 vdd.n4356 vdd.n4355 4.704
R46527 vdd.n27479 vdd.n27478 4.704
R46528 vdd.n25717 vdd.n25716 4.704
R46529 vdd.n25379 vdd.n25378 4.704
R46530 vdd.n17 vdd.n16 4.703
R46531 vdd.n25413 vdd.n25410 4.703
R46532 vdd.n31548 vdd.n31547 4.702
R46533 vdd.n1960 vdd.n1959 4.702
R46534 vdd.n11616 vdd.n11615 4.702
R46535 vdd.n21630 vdd.n21629 4.702
R46536 vdd.n14609 vdd.n8169 4.7
R46537 vdd.n18500 vdd.n18461 4.7
R46538 vdd.n19351 vdd.n19350 4.691
R46539 vdd.n19496 vdd.n19495 4.691
R46540 vdd.n19557 vdd.n19556 4.691
R46541 vdd.n19696 vdd.n19695 4.691
R46542 vdd.n19759 vdd.n19758 4.691
R46543 vdd.n20956 vdd.n20955 4.691
R46544 vdd.n20893 vdd.n20892 4.691
R46545 vdd.n20766 vdd.n20765 4.691
R46546 vdd.n20705 vdd.n20704 4.691
R46547 vdd.n20560 vdd.n20559 4.691
R46548 vdd.n20450 vdd.n20448 4.691
R46549 vdd.n20329 vdd.n20328 4.691
R46550 vdd.n20215 vdd.n20212 4.691
R46551 vdd.n20093 vdd.n20092 4.691
R46552 vdd.n11606 vdd.n11576 4.69
R46553 vdd.n21644 vdd.n21643 4.69
R46554 vdd.n14748 vdd.n8094 4.679
R46555 vdd.n14834 vdd.n8050 4.679
R46556 vdd.n14927 vdd.n14926 4.679
R46557 vdd.n25556 vdd.n25432 4.658
R46558 vdd.n32388 vdd.n32387 4.651
R46559 vdd.n3879 vdd.n3807 4.651
R46560 vdd.n33835 vdd.n33834 4.65
R46561 vdd.n33534 vdd.n33533 4.65
R46562 vdd.n33457 vdd.n33456 4.65
R46563 vdd.n33405 vdd.n33404 4.65
R46564 vdd.n34307 vdd.n34306 4.65
R46565 vdd.n34396 vdd.n34395 4.65
R46566 vdd.n34066 vdd.n34065 4.65
R46567 vdd.n35227 vdd.n35226 4.65
R46568 vdd.n35412 vdd.n35411 4.65
R46569 vdd.n35573 vdd.n35572 4.65
R46570 vdd.n34902 vdd.n34901 4.65
R46571 vdd.n34816 vdd.n34815 4.65
R46572 vdd.n34640 vdd.n34639 4.65
R46573 vdd.n810 vdd.n809 4.65
R46574 vdd.n646 vdd.n645 4.65
R46575 vdd.n776 vdd.n775 4.65
R46576 vdd.n726 vdd.n725 4.65
R46577 vdd.n201 vdd.n200 4.65
R46578 vdd.n437 vdd.n436 4.65
R46579 vdd.n471 vdd.n470 4.65
R46580 vdd.n6350 vdd.n6349 4.65
R46581 vdd.n6109 vdd.n6108 4.65
R46582 vdd.n5945 vdd.n5944 4.65
R46583 vdd.n5649 vdd.n5648 4.65
R46584 vdd.n5563 vdd.n5562 4.65
R46585 vdd.n5387 vdd.n5386 4.65
R46586 vdd.n4633 vdd.n4632 4.65
R46587 vdd.n4739 vdd.n4738 4.65
R46588 vdd.n5181 vdd.n5180 4.65
R46589 vdd.n4896 vdd.n4893 4.65
R46590 vdd.n4476 vdd.n4475 4.65
R46591 vdd.n4389 vdd.n4388 4.65
R46592 vdd.n4217 vdd.n4216 4.65
R46593 vdd.n33275 vdd.n33273 4.65
R46594 vdd.n37213 vdd.n37211 4.65
R46595 vdd.n32944 vdd.n32939 4.65
R46596 vdd.n38172 vdd.n38170 4.65
R46597 vdd.n33275 vdd.n33274 4.65
R46598 vdd.n37213 vdd.n37212 4.65
R46599 vdd.n32944 vdd.n32938 4.65
R46600 vdd.n38172 vdd.n38171 4.65
R46601 vdd.n31167 vdd.n31130 4.65
R46602 vdd.n31175 vdd.n31168 4.65
R46603 vdd.n28054 vdd.n28053 4.65
R46604 vdd.n27894 vdd.n27893 4.65
R46605 vdd.n28026 vdd.n28024 4.65
R46606 vdd.n29781 vdd.n29779 4.65
R46607 vdd.n28026 vdd.n28025 4.65
R46608 vdd.n29781 vdd.n29780 4.65
R46609 vdd.n30524 vdd.n30522 4.65
R46610 vdd.n30524 vdd.n30523 4.65
R46611 vdd.n27441 vdd.n27440 4.65
R46612 vdd.n27508 vdd.n27507 4.65
R46613 vdd.n27597 vdd.n27596 4.65
R46614 vdd.n25887 vdd.n25886 4.65
R46615 vdd.n25945 vdd.n25944 4.65
R46616 vdd.n26013 vdd.n26012 4.65
R46617 vdd.n25451 vdd.n25450 4.65
R46618 vdd.n25614 vdd.n25613 4.65
R46619 vdd.n25649 vdd.n25648 4.65
R46620 vdd.n3679 vdd.n3677 4.65
R46621 vdd.n2256 vdd.n2254 4.65
R46622 vdd.n2648 vdd.n2646 4.65
R46623 vdd.n3679 vdd.n3678 4.65
R46624 vdd.n2256 vdd.n2255 4.65
R46625 vdd.n2648 vdd.n2647 4.65
R46626 vdd.n36037 vdd.n36036 4.65
R46627 vdd.n36268 vdd.n36267 4.65
R46628 vdd.n36499 vdd.n36498 4.65
R46629 vdd.n36730 vdd.n36729 4.65
R46630 vdd.n36961 vdd.n36960 4.65
R46631 vdd.n37157 vdd.n37156 4.65
R46632 vdd.n35654 vdd.n35653 4.65
R46633 vdd.n37550 vdd.n37549 4.65
R46634 vdd.n38016 vdd.n38015 4.65
R46635 vdd.n37785 vdd.n37784 4.65
R46636 vdd.n28227 vdd.n28226 4.65
R46637 vdd.n28458 vdd.n28457 4.65
R46638 vdd.n28689 vdd.n28688 4.65
R46639 vdd.n28991 vdd.n28990 4.65
R46640 vdd.n30690 vdd.n30689 4.65
R46641 vdd.n2891 vdd.n2890 4.65
R46642 vdd.n3072 vdd.n3071 4.65
R46643 vdd.n3253 vdd.n3252 4.65
R46644 vdd.n3434 vdd.n3433 4.65
R46645 vdd.n3615 vdd.n3614 4.65
R46646 vdd.n2511 vdd.n2510 4.65
R46647 vdd.n1836 vdd.n1835 4.65
R46648 vdd.n1653 vdd.n1652 4.65
R46649 vdd.n1472 vdd.n1471 4.65
R46650 vdd.n1291 vdd.n1290 4.65
R46651 vdd.n26938 vdd.n26937 4.65
R46652 vdd.n27119 vdd.n27118 4.65
R46653 vdd.n27229 vdd.n27227 4.65
R46654 vdd.n31942 vdd.n31940 4.65
R46655 vdd.n32303 vdd.n32301 4.65
R46656 vdd.n27229 vdd.n27228 4.65
R46657 vdd.n31942 vdd.n31941 4.65
R46658 vdd.n32303 vdd.n32302 4.65
R46659 vdd.n26668 vdd.n26667 4.65
R46660 vdd.n32031 vdd.n32030 4.65
R46661 vdd.n10542 vdd.n10541 4.65
R46662 vdd.n10548 vdd.n10538 4.65
R46663 vdd.n10559 vdd.n10558 4.65
R46664 vdd.n12507 vdd.n10533 4.65
R46665 vdd.n12497 vdd.n12496 4.65
R46666 vdd.n12492 vdd.n10567 4.65
R46667 vdd.n10590 vdd.n10589 4.65
R46668 vdd.n12477 vdd.n10588 4.65
R46669 vdd.n12467 vdd.n12466 4.65
R46670 vdd.n10611 vdd.n10608 4.65
R46671 vdd.n10640 vdd.n10633 4.65
R46672 vdd.n10650 vdd.n10628 4.65
R46673 vdd.n12448 vdd.n10627 4.65
R46674 vdd.n12438 vdd.n12437 4.65
R46675 vdd.n10662 vdd.n10659 4.65
R46676 vdd.n10695 vdd.n10694 4.65
R46677 vdd.n12419 vdd.n10676 4.65
R46678 vdd.n12409 vdd.n12408 4.65
R46679 vdd.n12404 vdd.n10702 4.65
R46680 vdd.n10733 vdd.n10729 4.65
R46681 vdd.n10744 vdd.n10743 4.65
R46682 vdd.n12388 vdd.n10724 4.65
R46683 vdd.n12378 vdd.n12377 4.65
R46684 vdd.n10754 vdd.n10752 4.65
R46685 vdd.n10791 vdd.n10784 4.65
R46686 vdd.n10801 vdd.n10779 4.65
R46687 vdd.n12359 vdd.n10778 4.65
R46688 vdd.n12349 vdd.n12348 4.65
R46689 vdd.n10813 vdd.n10810 4.65
R46690 vdd.n10839 vdd.n10833 4.65
R46691 vdd.n10850 vdd.n10849 4.65
R46692 vdd.n12327 vdd.n10852 4.65
R46693 vdd.n10880 vdd.n10876 4.65
R46694 vdd.n10891 vdd.n10890 4.65
R46695 vdd.n12311 vdd.n10871 4.65
R46696 vdd.n12301 vdd.n12300 4.65
R46697 vdd.n12296 vdd.n10899 4.65
R46698 vdd.n10933 vdd.n10929 4.65
R46699 vdd.n10944 vdd.n10943 4.65
R46700 vdd.n10948 vdd.n10947 4.65
R46701 vdd.n10971 vdd.n10925 4.65
R46702 vdd.n10978 vdd.n10970 4.65
R46703 vdd.n10988 vdd.n10965 4.65
R46704 vdd.n12258 vdd.n10964 4.65
R46705 vdd.n12248 vdd.n12247 4.65
R46706 vdd.n11000 vdd.n10997 4.65
R46707 vdd.n11024 vdd.n11020 4.65
R46708 vdd.n12228 vdd.n11016 4.65
R46709 vdd.n12218 vdd.n12217 4.65
R46710 vdd.n12213 vdd.n11039 4.65
R46711 vdd.n11070 vdd.n11066 4.65
R46712 vdd.n11081 vdd.n11080 4.65
R46713 vdd.n12197 vdd.n11061 4.65
R46714 vdd.n12187 vdd.n12186 4.65
R46715 vdd.n12182 vdd.n11089 4.65
R46716 vdd.n11122 vdd.n11111 4.65
R46717 vdd.n12168 vdd.n11110 4.65
R46718 vdd.n12158 vdd.n12157 4.65
R46719 vdd.n11134 vdd.n11131 4.65
R46720 vdd.n11163 vdd.n11156 4.65
R46721 vdd.n11172 vdd.n11151 4.65
R46722 vdd.n12139 vdd.n11150 4.65
R46723 vdd.n12129 vdd.n12128 4.65
R46724 vdd.n11205 vdd.n11201 4.65
R46725 vdd.n11216 vdd.n11215 4.65
R46726 vdd.n12109 vdd.n11196 4.65
R46727 vdd.n12099 vdd.n12098 4.65
R46728 vdd.n12094 vdd.n11224 4.65
R46729 vdd.n11254 vdd.n11250 4.65
R46730 vdd.n11265 vdd.n11264 4.65
R46731 vdd.n12078 vdd.n11245 4.65
R46732 vdd.n11293 vdd.n11271 4.65
R46733 vdd.n11300 vdd.n11292 4.65
R46734 vdd.n11310 vdd.n11287 4.65
R46735 vdd.n12053 vdd.n11286 4.65
R46736 vdd.n12043 vdd.n12042 4.65
R46737 vdd.n11322 vdd.n11319 4.65
R46738 vdd.n11348 vdd.n11342 4.65
R46739 vdd.n11359 vdd.n11358 4.65
R46740 vdd.n12021 vdd.n11361 4.65
R46741 vdd.n11389 vdd.n11385 4.65
R46742 vdd.n11400 vdd.n11399 4.65
R46743 vdd.n12005 vdd.n11380 4.65
R46744 vdd.n11995 vdd.n11994 4.65
R46745 vdd.n11990 vdd.n11408 4.65
R46746 vdd.n11477 vdd.n11473 4.65
R46747 vdd.n11507 vdd.n11506 4.65
R46748 vdd.n11535 vdd.n11534 4.65
R46749 vdd.n14417 vdd.n14416 4.65
R46750 vdd.n14151 vdd.n14150 4.65
R46751 vdd.n13862 vdd.n13861 4.65
R46752 vdd.n13534 vdd.n8933 4.65
R46753 vdd.n13242 vdd.n9154 4.65
R46754 vdd.n9876 vdd.n9875 4.65
R46755 vdd.n9710 vdd.n9692 4.65
R46756 vdd.n9516 vdd.n9515 4.65
R46757 vdd.n9350 vdd.n9332 4.65
R46758 vdd.n10447 vdd.n10446 4.65
R46759 vdd.n10035 vdd.n10032 4.65
R46760 vdd.n12640 vdd.n12639 4.65
R46761 vdd.n12650 vdd.n10021 4.65
R46762 vdd.n10022 vdd.n9986 4.65
R46763 vdd.n10014 vdd.n10013 4.65
R46764 vdd.n10002 vdd.n9993 4.65
R46765 vdd.n9962 vdd.n9933 4.65
R46766 vdd.n9948 vdd.n9942 4.65
R46767 vdd.n9945 vdd.n9943 4.65
R46768 vdd.n12704 vdd.n9917 4.65
R46769 vdd.n12714 vdd.n9908 4.65
R46770 vdd.n9907 vdd.n9889 4.65
R46771 vdd.n9896 vdd.n9895 4.65
R46772 vdd.n12733 vdd.n9871 4.65
R46773 vdd.n9872 vdd.n9839 4.65
R46774 vdd.n9864 vdd.n9863 4.65
R46775 vdd.n9852 vdd.n9846 4.65
R46776 vdd.n9821 vdd.n9818 4.65
R46777 vdd.n12761 vdd.n12760 4.65
R46778 vdd.n12771 vdd.n9784 4.65
R46779 vdd.n9789 vdd.n9788 4.65
R46780 vdd.n12799 vdd.n9763 4.65
R46781 vdd.n12809 vdd.n9753 4.65
R46782 vdd.n9752 vdd.n9723 4.65
R46783 vdd.n9738 vdd.n9731 4.65
R46784 vdd.n9734 vdd.n9732 4.65
R46785 vdd.n12829 vdd.n9693 4.65
R46786 vdd.n9706 vdd.n9694 4.65
R46787 vdd.n9675 vdd.n9672 4.65
R46788 vdd.n12848 vdd.n12847 4.65
R46789 vdd.n12858 vdd.n9661 4.65
R46790 vdd.n9662 vdd.n9626 4.65
R46791 vdd.n9654 vdd.n9653 4.65
R46792 vdd.n9642 vdd.n9633 4.65
R46793 vdd.n9602 vdd.n9574 4.65
R46794 vdd.n9588 vdd.n9582 4.65
R46795 vdd.n9585 vdd.n9583 4.65
R46796 vdd.n12912 vdd.n9558 4.65
R46797 vdd.n12922 vdd.n9548 4.65
R46798 vdd.n9547 vdd.n9528 4.65
R46799 vdd.n9535 vdd.n9534 4.65
R46800 vdd.n12941 vdd.n9511 4.65
R46801 vdd.n9512 vdd.n9479 4.65
R46802 vdd.n9504 vdd.n9503 4.65
R46803 vdd.n9492 vdd.n9486 4.65
R46804 vdd.n9461 vdd.n9458 4.65
R46805 vdd.n12969 vdd.n12968 4.65
R46806 vdd.n12979 vdd.n9424 4.65
R46807 vdd.n9429 vdd.n9428 4.65
R46808 vdd.n13007 vdd.n9403 4.65
R46809 vdd.n13017 vdd.n9393 4.65
R46810 vdd.n9392 vdd.n9363 4.65
R46811 vdd.n9378 vdd.n9371 4.65
R46812 vdd.n9374 vdd.n9372 4.65
R46813 vdd.n13037 vdd.n9333 4.65
R46814 vdd.n9346 vdd.n9334 4.65
R46815 vdd.n9314 vdd.n9311 4.65
R46816 vdd.n13056 vdd.n13055 4.65
R46817 vdd.n13066 vdd.n9301 4.65
R46818 vdd.n9302 vdd.n9294 4.65
R46819 vdd.n10363 vdd.n10359 4.65
R46820 vdd.n10354 vdd.n10352 4.65
R46821 vdd.n10397 vdd.n10332 4.65
R46822 vdd.n10331 vdd.n10329 4.65
R46823 vdd.n10410 vdd.n10322 4.65
R46824 vdd.n10420 vdd.n10310 4.65
R46825 vdd.n10425 vdd.n10424 4.65
R46826 vdd.n10435 vdd.n10300 4.65
R46827 vdd.n10302 vdd.n10301 4.65
R46828 vdd.n10450 vdd.n10449 4.65
R46829 vdd.n10460 vdd.n10282 4.65
R46830 vdd.n10284 vdd.n10283 4.65
R46831 vdd.n11713 vdd.n11712 4.65
R46832 vdd.n11856 vdd.n11855 4.65
R46833 vdd.n9285 vdd.n9284 4.65
R46834 vdd.n13087 vdd.n13086 4.65
R46835 vdd.n13373 vdd.n13372 4.65
R46836 vdd.n13665 vdd.n13664 4.65
R46837 vdd.n13963 vdd.n8627 4.65
R46838 vdd.n14253 vdd.n8405 4.65
R46839 vdd.n14974 vdd.n14973 4.65
R46840 vdd.n14707 vdd.n14706 4.65
R46841 vdd.n14880 vdd.n14879 4.65
R46842 vdd.n14575 vdd.n8151 4.65
R46843 vdd.n14494 vdd.n8212 4.65
R46844 vdd.n23858 vdd.n23857 4.65
R46845 vdd.n24090 vdd.n24089 4.65
R46846 vdd.n23402 vdd.n23401 4.65
R46847 vdd.n23170 vdd.n23169 4.65
R46848 vdd.n22823 vdd.n22822 4.65
R46849 vdd.n22591 vdd.n22590 4.65
R46850 vdd.n16887 vdd.n16886 4.65
R46851 vdd.n16903 vdd.n16902 4.65
R46852 vdd.n16919 vdd.n16918 4.65
R46853 vdd.n16935 vdd.n16934 4.65
R46854 vdd.n16951 vdd.n16950 4.65
R46855 vdd.n16967 vdd.n16966 4.65
R46856 vdd.n16980 vdd.n16979 4.65
R46857 vdd.n16996 vdd.n16995 4.65
R46858 vdd.n17012 vdd.n17011 4.65
R46859 vdd.n17028 vdd.n17027 4.65
R46860 vdd.n17044 vdd.n17043 4.65
R46861 vdd.n17060 vdd.n17059 4.65
R46862 vdd.n17076 vdd.n17075 4.65
R46863 vdd.n17092 vdd.n17091 4.65
R46864 vdd.n17108 vdd.n17107 4.65
R46865 vdd.n17143 vdd.n17142 4.65
R46866 vdd.n17159 vdd.n17158 4.65
R46867 vdd.n17175 vdd.n17174 4.65
R46868 vdd.n17191 vdd.n17190 4.65
R46869 vdd.n17207 vdd.n17206 4.65
R46870 vdd.n17223 vdd.n17222 4.65
R46871 vdd.n17239 vdd.n17238 4.65
R46872 vdd.n17252 vdd.n17251 4.65
R46873 vdd.n17268 vdd.n17267 4.65
R46874 vdd.n17284 vdd.n17283 4.65
R46875 vdd.n17300 vdd.n17299 4.65
R46876 vdd.n17316 vdd.n17315 4.65
R46877 vdd.n17332 vdd.n17331 4.65
R46878 vdd.n17348 vdd.n17347 4.65
R46879 vdd.n17364 vdd.n17363 4.65
R46880 vdd.n17380 vdd.n17379 4.65
R46881 vdd.n17415 vdd.n17414 4.65
R46882 vdd.n17431 vdd.n17430 4.65
R46883 vdd.n17447 vdd.n17446 4.65
R46884 vdd.n17463 vdd.n17462 4.65
R46885 vdd.n17479 vdd.n17478 4.65
R46886 vdd.n17495 vdd.n17494 4.65
R46887 vdd.n17511 vdd.n17510 4.65
R46888 vdd.n17524 vdd.n17523 4.65
R46889 vdd.n17540 vdd.n17539 4.65
R46890 vdd.n17556 vdd.n17555 4.65
R46891 vdd.n17572 vdd.n17571 4.65
R46892 vdd.n17588 vdd.n17587 4.65
R46893 vdd.n17593 vdd.n17592 4.65
R46894 vdd.n17606 vdd.n17605 4.65
R46895 vdd.n17622 vdd.n17621 4.65
R46896 vdd.n17638 vdd.n17637 4.65
R46897 vdd.n17673 vdd.n17672 4.65
R46898 vdd.n17689 vdd.n17688 4.65
R46899 vdd.n17705 vdd.n17704 4.65
R46900 vdd.n17721 vdd.n17720 4.65
R46901 vdd.n17737 vdd.n17736 4.65
R46902 vdd.n17753 vdd.n17752 4.65
R46903 vdd.n17769 vdd.n17768 4.65
R46904 vdd.n17782 vdd.n17781 4.65
R46905 vdd.n17798 vdd.n17797 4.65
R46906 vdd.n17814 vdd.n17813 4.65
R46907 vdd.n17830 vdd.n17829 4.65
R46908 vdd.n17846 vdd.n17845 4.65
R46909 vdd.n17862 vdd.n17861 4.65
R46910 vdd.n17877 vdd.n17876 4.65
R46911 vdd.n17893 vdd.n17892 4.65
R46912 vdd.n17909 vdd.n17908 4.65
R46913 vdd.n17944 vdd.n17943 4.65
R46914 vdd.n17960 vdd.n17959 4.65
R46915 vdd.n17976 vdd.n17975 4.65
R46916 vdd.n17992 vdd.n17991 4.65
R46917 vdd.n18008 vdd.n18007 4.65
R46918 vdd.n18024 vdd.n18023 4.65
R46919 vdd.n18040 vdd.n18039 4.65
R46920 vdd.n18053 vdd.n18052 4.65
R46921 vdd.n18069 vdd.n18068 4.65
R46922 vdd.n18085 vdd.n18084 4.65
R46923 vdd.n18101 vdd.n18100 4.65
R46924 vdd.n18117 vdd.n18116 4.65
R46925 vdd.n18133 vdd.n18132 4.65
R46926 vdd.n18149 vdd.n18148 4.65
R46927 vdd.n18165 vdd.n18164 4.65
R46928 vdd.n18181 vdd.n18180 4.65
R46929 vdd.n18216 vdd.n18215 4.65
R46930 vdd.n18231 vdd.n18230 4.65
R46931 vdd.n18246 vdd.n18245 4.65
R46932 vdd.n18261 vdd.n18260 4.65
R46933 vdd.n18276 vdd.n18275 4.65
R46934 vdd.n18291 vdd.n18290 4.65
R46935 vdd.n18306 vdd.n18305 4.65
R46936 vdd.n18333 vdd.n18332 4.65
R46937 vdd.n18372 vdd.n18371 4.65
R46938 vdd.n16309 vdd.n16308 4.65
R46939 vdd.n16053 vdd.n16052 4.65
R46940 vdd.n15797 vdd.n15796 4.65
R46941 vdd.n15541 vdd.n15540 4.65
R46942 vdd.n15313 vdd.n15312 4.65
R46943 vdd.n16541 vdd.n16540 4.65
R46944 vdd.n16524 vdd.n16523 4.65
R46945 vdd.n16507 vdd.n16506 4.65
R46946 vdd.n16490 vdd.n16489 4.65
R46947 vdd.n16470 vdd.n16469 4.65
R46948 vdd.n16453 vdd.n16452 4.65
R46949 vdd.n16432 vdd.n16431 4.65
R46950 vdd.n16415 vdd.n16414 4.65
R46951 vdd.n16398 vdd.n16397 4.65
R46952 vdd.n16381 vdd.n16380 4.65
R46953 vdd.n16364 vdd.n16363 4.65
R46954 vdd.n16347 vdd.n16346 4.65
R46955 vdd.n16330 vdd.n16329 4.65
R46956 vdd.n16304 vdd.n16303 4.65
R46957 vdd.n16285 vdd.n16284 4.65
R46958 vdd.n16268 vdd.n16267 4.65
R46959 vdd.n16251 vdd.n16250 4.65
R46960 vdd.n16234 vdd.n16233 4.65
R46961 vdd.n16214 vdd.n16213 4.65
R46962 vdd.n16197 vdd.n16196 4.65
R46963 vdd.n16176 vdd.n16175 4.65
R46964 vdd.n16159 vdd.n16158 4.65
R46965 vdd.n16142 vdd.n16141 4.65
R46966 vdd.n16125 vdd.n16124 4.65
R46967 vdd.n16108 vdd.n16107 4.65
R46968 vdd.n16091 vdd.n16090 4.65
R46969 vdd.n16074 vdd.n16073 4.65
R46970 vdd.n16048 vdd.n16047 4.65
R46971 vdd.n16029 vdd.n16028 4.65
R46972 vdd.n16012 vdd.n16011 4.65
R46973 vdd.n15995 vdd.n15994 4.65
R46974 vdd.n15978 vdd.n15977 4.65
R46975 vdd.n15958 vdd.n15957 4.65
R46976 vdd.n15941 vdd.n15940 4.65
R46977 vdd.n15920 vdd.n15919 4.65
R46978 vdd.n15903 vdd.n15902 4.65
R46979 vdd.n15886 vdd.n15885 4.65
R46980 vdd.n15869 vdd.n15868 4.65
R46981 vdd.n15852 vdd.n15851 4.65
R46982 vdd.n15835 vdd.n15834 4.65
R46983 vdd.n15818 vdd.n15817 4.65
R46984 vdd.n15792 vdd.n15791 4.65
R46985 vdd.n15773 vdd.n15772 4.65
R46986 vdd.n15756 vdd.n15755 4.65
R46987 vdd.n15739 vdd.n15738 4.65
R46988 vdd.n15722 vdd.n15721 4.65
R46989 vdd.n15702 vdd.n15701 4.65
R46990 vdd.n15685 vdd.n15684 4.65
R46991 vdd.n15664 vdd.n15663 4.65
R46992 vdd.n15647 vdd.n15646 4.65
R46993 vdd.n15630 vdd.n15629 4.65
R46994 vdd.n15613 vdd.n15612 4.65
R46995 vdd.n15596 vdd.n15595 4.65
R46996 vdd.n15579 vdd.n15578 4.65
R46997 vdd.n15562 vdd.n15561 4.65
R46998 vdd.n15536 vdd.n15535 4.65
R46999 vdd.n15517 vdd.n15516 4.65
R47000 vdd.n15500 vdd.n15499 4.65
R47001 vdd.n15483 vdd.n15482 4.65
R47002 vdd.n15466 vdd.n15465 4.65
R47003 vdd.n15446 vdd.n15445 4.65
R47004 vdd.n15432 vdd.n15431 4.65
R47005 vdd.n15414 vdd.n15413 4.65
R47006 vdd.n15399 vdd.n15398 4.65
R47007 vdd.n15385 vdd.n15384 4.65
R47008 vdd.n15371 vdd.n15370 4.65
R47009 vdd.n15357 vdd.n15356 4.65
R47010 vdd.n15342 vdd.n15341 4.65
R47011 vdd.n15328 vdd.n15327 4.65
R47012 vdd.n15308 vdd.n15307 4.65
R47013 vdd.n15292 vdd.n15291 4.65
R47014 vdd.n15278 vdd.n15277 4.65
R47015 vdd.n18635 vdd.n18634 4.65
R47016 vdd.n18894 vdd.n18893 4.65
R47017 vdd.n21012 vdd.n21011 4.65
R47018 vdd.n21260 vdd.n21259 4.65
R47019 vdd.n21519 vdd.n21518 4.65
R47020 vdd.n20026 vdd.n20025 4.65
R47021 vdd.n20391 vdd.n20390 4.65
R47022 vdd.n20155 vdd.n20154 4.65
R47023 vdd.n19987 vdd.n19986 4.65
R47024 vdd.n19969 vdd.n19968 4.65
R47025 vdd.n19526 vdd.n19525 4.65
R47026 vdd.n19727 vdd.n19726 4.65
R47027 vdd.n20924 vdd.n20923 4.65
R47028 vdd.n20735 vdd.n20734 4.65
R47029 vdd.n19299 vdd.n19298 4.65
R47030 vdd.n21789 vdd.n21788 4.65
R47031 vdd.n21947 vdd.n21946 4.65
R47032 vdd.n21746 vdd.n21745 4.65
R47033 vdd.n25026 vdd.n25025 4.65
R47034 vdd.n24600 vdd.n24599 4.65
R47035 vdd.n25165 vdd.n25164 4.65
R47036 vdd.n24749 vdd.n24748 4.65
R47037 vdd.n25091 vdd.n25090 4.65
R47038 vdd.n24673 vdd.n24672 4.65
R47039 vdd.n10246 vdd.n10224 4.65
R47040 vdd.n16670 vdd.n16669 4.65
R47041 vdd.n31158 vdd.n31157 4.648
R47042 vdd.n32528 vdd.n32408 4.621
R47043 vdd.n32077 vdd.n32071 4.61
R47044 vdd.n33643 vdd.n33642 4.596
R47045 vdd.n33331 vdd.n33330 4.596
R47046 vdd.n33404 vdd.n33403 4.596
R47047 vdd.n34294 vdd.n34293 4.596
R47048 vdd.n33995 vdd.n33994 4.596
R47049 vdd.n35157 vdd.n35156 4.596
R47050 vdd.n35560 vdd.n35559 4.596
R47051 vdd.n34910 vdd.n34909 4.596
R47052 vdd.n34575 vdd.n34574 4.596
R47053 vdd.n1080 vdd.n1079 4.596
R47054 vdd.n620 vdd.n619 4.596
R47055 vdd.n725 vdd.n724 4.596
R47056 vdd.n142 vdd.n141 4.596
R47057 vdd.n436 vdd.n435 4.596
R47058 vdd.n522 vdd.n521 4.596
R47059 vdd.n6286 vdd.n6285 4.596
R47060 vdd.n5953 vdd.n5952 4.596
R47061 vdd.n5657 vdd.n5656 4.596
R47062 vdd.n5322 vdd.n5321 4.596
R47063 vdd.n4639 vdd.n4638 4.596
R47064 vdd.n5131 vdd.n5130 4.596
R47065 vdd.n4484 vdd.n4483 4.596
R47066 vdd.n4153 vdd.n4152 4.596
R47067 vdd.n27431 vdd.n27430 4.596
R47068 vdd.n27628 vdd.n27627 4.596
R47069 vdd.n25877 vdd.n25876 4.596
R47070 vdd.n26049 vdd.n26048 4.596
R47071 vdd.n25656 vdd.n25655 4.596
R47072 vdd.n11545 vdd.n11451 4.592
R47073 vdd.n18383 vdd.n15026 4.592
R47074 vdd.n33907 vdd.n33906 4.589
R47075 vdd.n35076 vdd.n35075 4.589
R47076 vdd.n34489 vdd.n34488 4.589
R47077 vdd.n6181 vdd.n6180 4.589
R47078 vdd.n5236 vdd.n5235 4.589
R47079 vdd.n4986 vdd.n4985 4.589
R47080 vdd.n4066 vdd.n4065 4.589
R47081 vdd.n27541 vdd.n27540 4.589
R47082 vdd.n25978 vdd.n25977 4.589
R47083 vdd.n13276 vdd.n9157 4.587
R47084 vdd.n13359 vdd.n13355 4.587
R47085 vdd.n13651 vdd.n13647 4.587
R47086 vdd.n13703 vdd.t128 4.587
R47087 vdd.n13856 vdd.n8718 4.587
R47088 vdd.n13967 vdd.n8621 4.587
R47089 vdd.n14145 vdd.n8496 4.587
R47090 vdd.n14257 vdd.n8399 4.587
R47091 vdd.n14461 vdd.n8239 4.587
R47092 vdd.n34385 vdd.n34384 4.582
R47093 vdd.n35404 vdd.n35403 4.582
R47094 vdd.n34808 vdd.n34807 4.582
R47095 vdd.n6098 vdd.n6097 4.582
R47096 vdd.n5555 vdd.n5554 4.582
R47097 vdd.n4749 vdd.n4748 4.582
R47098 vdd.n4381 vdd.n4380 4.582
R47099 vdd.n27496 vdd.n27495 4.582
R47100 vdd.n25933 vdd.n25932 4.582
R47101 vdd.n11793 vdd.n11792 4.582
R47102 vdd.n21884 vdd.n21883 4.582
R47103 vdd.n44 vdd.n43 4.574
R47104 vdd.n33520 vdd.n33519 4.567
R47105 vdd.n1001 vdd.n1000 4.567
R47106 vdd.n11905 vdd.n11790 4.563
R47107 vdd.n21996 vdd.n21881 4.563
R47108 vdd.n4840 vdd.n4839 4.56
R47109 vdd.n11688 vdd.n11681 4.559
R47110 vdd.n21761 vdd.n21760 4.559
R47111 vdd.n11772 vdd.n11667 4.559
R47112 vdd.n11835 vdd.n11804 4.559
R47113 vdd.n21864 vdd.n21860 4.559
R47114 vdd.n21926 vdd.n21895 4.559
R47115 vdd.n33741 vdd.n33740 4.558
R47116 vdd.n33698 vdd.n33576 4.558
R47117 vdd.n33363 vdd.n33291 4.558
R47118 vdd.n33367 vdd.n33288 4.558
R47119 vdd.n34340 vdd.n34241 4.558
R47120 vdd.n34103 vdd.n34102 4.558
R47121 vdd.n35607 vdd.n35468 4.558
R47122 vdd.n35486 vdd.n35481 4.558
R47123 vdd.n35019 vdd.n34883 4.558
R47124 vdd.n34961 vdd.n34960 4.558
R47125 vdd.n921 vdd.n920 4.558
R47126 vdd.n1165 vdd.n1052 4.558
R47127 vdd.n682 vdd.n601 4.558
R47128 vdd.n687 vdd.n598 4.558
R47129 vdd.n577 vdd.n506 4.558
R47130 vdd.n573 vdd.n509 4.558
R47131 vdd.n6042 vdd.n5926 4.558
R47132 vdd.n5811 vdd.n5810 4.558
R47133 vdd.n5766 vdd.n5630 4.558
R47134 vdd.n5708 vdd.n5707 4.558
R47135 vdd.n4706 vdd.n4619 4.558
R47136 vdd.n4830 vdd.n4829 4.558
R47137 vdd.n4596 vdd.n4457 4.558
R47138 vdd.n4535 vdd.n4534 4.558
R47139 vdd.n32858 vdd.n32857 4.558
R47140 vdd.n33177 vdd.n33166 4.558
R47141 vdd.n37127 vdd.n37121 4.558
R47142 vdd.n33023 vdd.n33005 4.558
R47143 vdd.n37315 vdd.n37298 4.558
R47144 vdd.n37516 vdd.n37501 4.558
R47145 vdd.n32858 vdd.n32851 4.558
R47146 vdd.n37315 vdd.n37305 4.558
R47147 vdd.n33023 vdd.n33020 4.558
R47148 vdd.n33177 vdd.n33164 4.558
R47149 vdd.n37127 vdd.n37120 4.558
R47150 vdd.n37516 vdd.n37499 4.558
R47151 vdd.n37262 vdd.n37242 4.558
R47152 vdd.n33229 vdd.n33228 4.558
R47153 vdd.n37064 vdd.n37063 4.558
R47154 vdd.n33076 vdd.n33065 4.558
R47155 vdd.n37457 vdd.n37448 4.558
R47156 vdd.n32919 vdd.n32897 4.558
R47157 vdd.n28804 vdd.n28143 4.558
R47158 vdd.n28103 vdd.n28102 4.558
R47159 vdd.n28130 vdd.n28121 4.558
R47160 vdd.n27824 vdd.n27795 4.558
R47161 vdd.n29034 vdd.n29033 4.558
R47162 vdd.n27853 vdd.n27851 4.558
R47163 vdd.n29848 vdd.n29695 4.558
R47164 vdd.n28925 vdd.n28080 4.558
R47165 vdd.n28928 vdd.n28078 4.558
R47166 vdd.n27944 vdd.n27904 4.558
R47167 vdd.n27926 vdd.n27925 4.558
R47168 vdd.n30631 vdd.n30215 4.558
R47169 vdd.n30626 vdd.n30625 4.558
R47170 vdd.n30626 vdd.n30224 4.558
R47171 vdd.n30631 vdd.n30213 4.558
R47172 vdd.n27926 vdd.n27918 4.558
R47173 vdd.n27944 vdd.n27902 4.558
R47174 vdd.n28928 vdd.n28076 4.558
R47175 vdd.n28925 vdd.n28079 4.558
R47176 vdd.n30571 vdd.n30311 4.558
R47177 vdd.n27384 vdd.n27383 4.558
R47178 vdd.n27464 vdd.n27287 4.558
R47179 vdd.n25827 vdd.n25826 4.558
R47180 vdd.n25910 vdd.n25733 4.558
R47181 vdd.n25495 vdd.n25494 4.558
R47182 vdd.n25568 vdd.n25566 4.558
R47183 vdd.n25630 vdd.n25629 4.558
R47184 vdd.n3944 vdd.n3781 4.558
R47185 vdd.n3932 vdd.n3931 4.558
R47186 vdd.n2393 vdd.n2104 4.558
R47187 vdd.n2556 vdd.n2555 4.558
R47188 vdd.n1893 vdd.n1216 4.558
R47189 vdd.n1884 vdd.n1883 4.558
R47190 vdd.n3944 vdd.n3779 4.558
R47191 vdd.n3932 vdd.n3789 4.558
R47192 vdd.n2393 vdd.n2102 4.558
R47193 vdd.n2556 vdd.n2409 4.558
R47194 vdd.n1893 vdd.n1214 4.558
R47195 vdd.n1884 vdd.n1226 4.558
R47196 vdd.n2000 vdd.n1960 4.558
R47197 vdd.n1991 vdd.n1985 4.558
R47198 vdd.n2298 vdd.n2130 4.558
R47199 vdd.n2285 vdd.n2135 4.558
R47200 vdd.n4013 vdd.n3723 4.558
R47201 vdd.n3712 vdd.n2685 4.558
R47202 vdd.n31744 vdd.n31743 4.558
R47203 vdd.n31762 vdd.n31735 4.558
R47204 vdd.n32088 vdd.n31584 4.558
R47205 vdd.n32111 vdd.n31581 4.558
R47206 vdd.n32487 vdd.n32420 4.558
R47207 vdd.n32473 vdd.n32472 4.558
R47208 vdd.n31744 vdd.n31742 4.558
R47209 vdd.n31762 vdd.n31733 4.558
R47210 vdd.n32088 vdd.n31583 4.558
R47211 vdd.n32111 vdd.n31579 4.558
R47212 vdd.n32487 vdd.n32418 4.558
R47213 vdd.n32473 vdd.n32422 4.558
R47214 vdd.n31181 vdd.n31129 4.558
R47215 vdd.n31121 vdd.n31027 4.558
R47216 vdd.n32254 vdd.n31545 4.558
R47217 vdd.n32233 vdd.n31548 4.558
R47218 vdd.n31881 vdd.n31678 4.558
R47219 vdd.n31869 vdd.n31694 4.558
R47220 vdd.n13948 vdd.n8597 4.558
R47221 vdd.n14001 vdd.n8598 4.558
R47222 vdd.n14238 vdd.n8375 4.558
R47223 vdd.n14292 vdd.n8376 4.558
R47224 vdd.n14607 vdd.n8177 4.558
R47225 vdd.n14608 vdd.n8176 4.558
R47226 vdd.n11616 vdd.n11611 4.558
R47227 vdd.n13384 vdd.n9058 4.558
R47228 vdd.n13386 vdd.n13385 4.558
R47229 vdd.n13676 vdd.n8838 4.558
R47230 vdd.n13678 vdd.n13677 4.558
R47231 vdd.n13211 vdd.n9173 4.558
R47232 vdd.n13254 vdd.n9174 4.558
R47233 vdd.n13504 vdd.n8953 4.558
R47234 vdd.n13545 vdd.n8954 4.558
R47235 vdd.n13785 vdd.n8734 4.558
R47236 vdd.n13830 vdd.n8735 4.558
R47237 vdd.n14113 vdd.n8516 4.558
R47238 vdd.n14112 vdd.n8518 4.558
R47239 vdd.n14401 vdd.n8299 4.558
R47240 vdd.n14403 vdd.n14402 4.558
R47241 vdd.n14795 vdd.n8066 4.558
R47242 vdd.n14794 vdd.n8067 4.558
R47243 vdd.n19020 vdd.n18442 4.558
R47244 vdd.n19019 vdd.n18443 4.558
R47245 vdd.n18761 vdd.n18446 4.558
R47246 vdd.n18760 vdd.n18447 4.558
R47247 vdd.n18502 vdd.n18450 4.558
R47248 vdd.n18501 vdd.n18451 4.558
R47249 vdd.n21652 vdd.n21630 4.558
R47250 vdd.n21386 vdd.n18434 4.558
R47251 vdd.n21385 vdd.n18435 4.558
R47252 vdd.n21127 vdd.n18438 4.558
R47253 vdd.n21126 vdd.n18439 4.558
R47254 vdd.n20270 vdd.n20013 4.558
R47255 vdd.n20271 vdd.n20001 4.558
R47256 vdd.n20628 vdd.n19954 4.558
R47257 vdd.n20629 vdd.n19953 4.558
R47258 vdd.n20830 vdd.n19897 4.558
R47259 vdd.n20831 vdd.n19896 4.558
R47260 vdd.n19829 vdd.n19173 4.558
R47261 vdd.n19827 vdd.n19176 4.558
R47262 vdd.n19626 vdd.n19229 4.558
R47263 vdd.n19625 vdd.n19232 4.558
R47264 vdd.n19423 vdd.n19285 4.558
R47265 vdd.n19422 vdd.n19288 4.558
R47266 vdd.n24833 vdd.n24515 4.558
R47267 vdd.n25251 vdd.n24984 4.558
R47268 vdd.n3903 vdd.n3902 4.546
R47269 vdd.n25509 vdd.n25508 4.533
R47270 vdd.n31785 vdd.n31775 4.521
R47271 vdd.n25091 vdd.n24882 4.518
R47272 vdd.n34115 vdd.n34114 4.517
R47273 vdd.n35471 vdd.n35470 4.517
R47274 vdd.n34949 vdd.n34948 4.517
R47275 vdd.n5823 vdd.n5822 4.517
R47276 vdd.n5696 vdd.n5695 4.517
R47277 vdd.n4523 vdd.n4522 4.517
R47278 vdd.n30274 vdd.n30267 4.517
R47279 vdd.n30276 vdd.n30274 4.517
R47280 vdd.n31260 vdd.n31253 4.517
R47281 vdd.n30530 vdd.n30526 4.517
R47282 vdd.n35885 vdd.n35878 4.517
R47283 vdd.n35962 vdd.n35955 4.517
R47284 vdd.n36116 vdd.n36109 4.517
R47285 vdd.n36193 vdd.n36186 4.517
R47286 vdd.n36347 vdd.n36340 4.517
R47287 vdd.n36424 vdd.n36417 4.517
R47288 vdd.n36578 vdd.n36571 4.517
R47289 vdd.n36655 vdd.n36648 4.517
R47290 vdd.n36809 vdd.n36802 4.517
R47291 vdd.n36886 vdd.n36879 4.517
R47292 vdd.n33283 vdd.n33279 4.517
R47293 vdd.n33220 vdd.n33213 4.517
R47294 vdd.n37219 vdd.n37215 4.517
R47295 vdd.n37279 vdd.n37272 4.517
R47296 vdd.n37420 vdd.n37413 4.517
R47297 vdd.n37482 vdd.n37475 4.517
R47298 vdd.n38168 vdd.n38161 4.517
R47299 vdd.n38095 vdd.n38088 4.517
R47300 vdd.n37941 vdd.n37934 4.517
R47301 vdd.n37864 vdd.n37857 4.517
R47302 vdd.n37710 vdd.n37703 4.517
R47303 vdd.n37633 vdd.n37626 4.517
R47304 vdd.n28306 vdd.n28299 4.517
R47305 vdd.n28383 vdd.n28376 4.517
R47306 vdd.n28537 vdd.n28530 4.517
R47307 vdd.n28614 vdd.n28607 4.517
R47308 vdd.n28768 vdd.n28761 4.517
R47309 vdd.n28175 vdd.n28168 4.517
R47310 vdd.n28990 vdd.n28983 4.517
R47311 vdd.n27748 vdd.n27747 4.517
R47312 vdd.n27794 vdd.n27787 4.517
R47313 vdd.n27289 vdd.n27288 4.517
R47314 vdd.n25832 vdd.n25831 4.517
R47315 vdd.n1769 vdd.n1765 4.517
R47316 vdd.n1714 vdd.n1710 4.517
R47317 vdd.n1594 vdd.n1590 4.517
R47318 vdd.n1533 vdd.n1529 4.517
R47319 vdd.n1413 vdd.n1409 4.517
R47320 vdd.n1352 vdd.n1348 4.517
R47321 vdd.n26818 vdd.n26814 4.517
R47322 vdd.n26879 vdd.n26875 4.517
R47323 vdd.n26999 vdd.n26995 4.517
R47324 vdd.n27060 vdd.n27056 4.517
R47325 vdd.n27180 vdd.n27176 4.517
R47326 vdd.n2771 vdd.n2767 4.517
R47327 vdd.n2832 vdd.n2828 4.517
R47328 vdd.n2952 vdd.n2948 4.517
R47329 vdd.n3013 vdd.n3009 4.517
R47330 vdd.n3133 vdd.n3129 4.517
R47331 vdd.n3194 vdd.n3190 4.517
R47332 vdd.n3314 vdd.n3310 4.517
R47333 vdd.n3375 vdd.n3371 4.517
R47334 vdd.n3495 vdd.n3491 4.517
R47335 vdd.n3556 vdd.n3552 4.517
R47336 vdd.n13184 vdd.n9220 4.517
R47337 vdd.n13184 vdd.n13183 4.517
R47338 vdd.n13274 vdd.n9161 4.517
R47339 vdd.n13274 vdd.n9148 4.517
R47340 vdd.n13478 vdd.n9000 4.517
R47341 vdd.n13478 vdd.n13477 4.517
R47342 vdd.n13566 vdd.n8939 4.517
R47343 vdd.n13566 vdd.n8927 4.517
R47344 vdd.n13758 vdd.n8783 4.517
R47345 vdd.n13758 vdd.n13757 4.517
R47346 vdd.n13854 vdd.n8723 4.517
R47347 vdd.n13854 vdd.n8724 4.517
R47348 vdd.n14040 vdd.n8559 4.517
R47349 vdd.n8559 vdd.n8557 4.517
R47350 vdd.n14143 vdd.n8502 4.517
R47351 vdd.n14143 vdd.n8503 4.517
R47352 vdd.n14348 vdd.n14347 4.517
R47353 vdd.n14349 vdd.n14348 4.517
R47354 vdd.n14459 vdd.n8244 4.517
R47355 vdd.n14459 vdd.n8245 4.517
R47356 vdd.n14654 vdd.n8149 4.517
R47357 vdd.n14649 vdd.n8150 4.517
R47358 vdd.n14764 vdd.n14763 4.517
R47359 vdd.n14771 vdd.n14770 4.517
R47360 vdd.n14826 vdd.n8058 4.517
R47361 vdd.n14821 vdd.n8059 4.517
R47362 vdd.n14938 vdd.n8003 4.517
R47363 vdd.n14940 vdd.n7983 4.517
R47364 vdd.n13155 vdd.n9235 4.517
R47365 vdd.n13362 vdd.n13361 4.517
R47366 vdd.n13361 vdd.n9075 4.517
R47367 vdd.n13448 vdd.n9014 4.517
R47368 vdd.n13448 vdd.n9011 4.517
R47369 vdd.n13654 vdd.n13653 4.517
R47370 vdd.n13653 vdd.n8855 4.517
R47371 vdd.n13739 vdd.n8794 4.517
R47372 vdd.n13739 vdd.n8792 4.517
R47373 vdd.n13941 vdd.n8637 4.517
R47374 vdd.n13942 vdd.n13941 4.517
R47375 vdd.n8584 vdd.n8581 4.517
R47376 vdd.n14024 vdd.n8581 4.517
R47377 vdd.n14231 vdd.n8415 4.517
R47378 vdd.n14232 vdd.n14231 4.517
R47379 vdd.n14312 vdd.n8362 4.517
R47380 vdd.n14312 vdd.n8359 4.517
R47381 vdd.n14557 vdd.n14556 4.517
R47382 vdd.n14556 vdd.n8192 4.517
R47383 vdd.n24269 vdd.n24268 4.517
R47384 vdd.n24278 vdd.n24277 4.517
R47385 vdd.n24166 vdd.n24165 4.517
R47386 vdd.n24000 vdd.n23999 4.517
R47387 vdd.n23934 vdd.n23933 4.517
R47388 vdd.n23768 vdd.n23767 4.517
R47389 vdd.n23702 vdd.n23701 4.517
R47390 vdd.n23080 vdd.n23079 4.517
R47391 vdd.n23246 vdd.n23245 4.517
R47392 vdd.n23312 vdd.n23311 4.517
R47393 vdd.n23478 vdd.n23477 4.517
R47394 vdd.n23544 vdd.n23543 4.517
R47395 vdd.n22501 vdd.n22500 4.517
R47396 vdd.n22667 vdd.n22666 4.517
R47397 vdd.n22733 vdd.n22732 4.517
R47398 vdd.n22899 vdd.n22898 4.517
R47399 vdd.n22965 vdd.n22964 4.517
R47400 vdd.n22441 vdd.n22440 4.517
R47401 vdd.n22450 vdd.n22449 4.517
R47402 vdd.n22254 vdd.n22243 4.517
R47403 vdd.n22245 vdd.n22244 4.517
R47404 vdd.n22297 vdd.n22296 4.517
R47405 vdd.n22306 vdd.n22305 4.517
R47406 vdd.n22130 vdd.n22119 4.517
R47407 vdd.n22121 vdd.n22120 4.517
R47408 vdd.n19385 vdd.n19376 4.517
R47409 vdd.n19466 vdd.n19457 4.517
R47410 vdd.n19591 vdd.n19582 4.517
R47411 vdd.n19666 vdd.n19657 4.517
R47412 vdd.n19793 vdd.n19784 4.517
R47413 vdd.n20990 vdd.n20981 4.517
R47414 vdd.n19892 vdd.n19883 4.517
R47415 vdd.n20799 vdd.n20790 4.517
R47416 vdd.n20675 vdd.n20666 4.517
R47417 vdd.n20594 vdd.n20585 4.517
R47418 vdd.n21618 vdd.n21601 4.517
R47419 vdd.n21432 vdd.n21423 4.517
R47420 vdd.n21351 vdd.n21342 4.517
R47421 vdd.n21173 vdd.n21164 4.517
R47422 vdd.n21089 vdd.n21088 4.517
R47423 vdd.n19066 vdd.n19057 4.517
R47424 vdd.n18985 vdd.n18976 4.517
R47425 vdd.n18807 vdd.n18798 4.517
R47426 vdd.n18726 vdd.n18717 4.517
R47427 vdd.n18548 vdd.n18539 4.517
R47428 vdd.n19982 vdd.n19981 4.517
R47429 vdd.n19985 vdd.n19984 4.517
R47430 vdd.n20291 vdd.n20290 4.517
R47431 vdd.n20241 vdd.n20240 4.517
R47432 vdd.n20028 vdd.n20027 4.517
R47433 vdd.n24675 vdd.n24674 4.517
R47434 vdd.n24812 vdd.n24811 4.517
R47435 vdd.n25230 vdd.n25229 4.517
R47436 vdd.n25093 vdd.n25092 4.517
R47437 vdd.n10180 vdd.n10092 4.51
R47438 vdd.n11684 vdd.n11683 4.505
R47439 vdd.n11867 vdd.n11866 4.505
R47440 vdd.n21958 vdd.n21957 4.505
R47441 vdd.n11917 vdd.n11787 4.503
R47442 vdd.n11760 vdd.n11679 4.503
R47443 vdd.n11899 vdd.n11795 4.503
R47444 vdd.n21990 vdd.n21886 4.503
R47445 vdd.n11767 vdd.n11669 4.503
R47446 vdd.n11789 vdd.n11788 4.502
R47447 vdd.n21880 vdd.n21879 4.502
R47448 vdd.n11666 vdd.n11665 4.501
R47449 vdd.n11875 vdd.n11806 4.501
R47450 vdd.n21966 vdd.n21897 4.501
R47451 vdd.n27331 vdd.n27330 4.5
R47452 vdd.n27343 vdd.n27342 4.5
R47453 vdd.n27351 vdd.n27350 4.5
R47454 vdd.n27357 vdd.n27356 4.5
R47455 vdd.n27301 vdd.n27300 4.5
R47456 vdd.n27295 vdd.n27294 4.5
R47457 vdd.n27372 vdd.n27371 4.5
R47458 vdd.n27380 vdd.n27379 4.5
R47459 vdd.n27398 vdd.n27397 4.5
R47460 vdd.n27443 vdd.n27442 4.5
R47461 vdd.n27454 vdd.n27453 4.5
R47462 vdd.n27463 vdd.n27462 4.5
R47463 vdd.n27278 vdd.n27277 4.5
R47464 vdd.n27475 vdd.n27474 4.5
R47465 vdd.n27270 vdd.n27269 4.5
R47466 vdd.n27499 vdd.n27498 4.5
R47467 vdd.n27544 vdd.n27543 4.5
R47468 vdd.n27555 vdd.n27554 4.5
R47469 vdd.n27567 vdd.n27566 4.5
R47470 vdd.n27579 vdd.n27578 4.5
R47471 vdd.n27588 vdd.n27587 4.5
R47472 vdd.n27600 vdd.n27599 4.5
R47473 vdd.n27260 vdd.n27259 4.5
R47474 vdd.n27618 vdd.n27617 4.5
R47475 vdd.n25783 vdd.n25782 4.5
R47476 vdd.n25795 vdd.n25794 4.5
R47477 vdd.n25803 vdd.n25802 4.5
R47478 vdd.n25809 vdd.n25808 4.5
R47479 vdd.n25753 vdd.n25752 4.5
R47480 vdd.n25747 vdd.n25746 4.5
R47481 vdd.n25740 vdd.n25739 4.5
R47482 vdd.n25823 vdd.n25822 4.5
R47483 vdd.n25844 vdd.n25843 4.5
R47484 vdd.n25889 vdd.n25888 4.5
R47485 vdd.n25900 vdd.n25899 4.5
R47486 vdd.n25909 vdd.n25908 4.5
R47487 vdd.n25724 vdd.n25723 4.5
R47488 vdd.n25713 vdd.n25712 4.5
R47489 vdd.n25925 vdd.n25924 4.5
R47490 vdd.n25936 vdd.n25935 4.5
R47491 vdd.n25981 vdd.n25980 4.5
R47492 vdd.n25992 vdd.n25991 4.5
R47493 vdd.n25703 vdd.n25702 4.5
R47494 vdd.n25692 vdd.n25691 4.5
R47495 vdd.n26004 vdd.n26003 4.5
R47496 vdd.n26016 vdd.n26015 4.5
R47497 vdd.n26028 vdd.n26027 4.5
R47498 vdd.n26039 vdd.n26038 4.5
R47499 vdd.n25446 vdd.n25445 4.5
R47500 vdd.n25488 vdd.n25487 4.5
R47501 vdd.n25505 vdd.n25504 4.5
R47502 vdd.n25513 vdd.n25511 4.5
R47503 vdd.n25523 vdd.n25522 4.5
R47504 vdd.n25530 vdd.n25529 4.5
R47505 vdd.n25441 vdd.n25440 4.5
R47506 vdd.n25543 vdd.n25542 4.5
R47507 vdd.n25579 vdd.n25578 4.5
R47508 vdd.n25597 vdd.n25596 4.5
R47509 vdd.n25607 vdd.n25606 4.5
R47510 vdd.n25621 vdd.n25620 4.5
R47511 vdd.n25414 vdd.n25413 4.5
R47512 vdd.n25403 vdd.n25402 4.5
R47513 vdd.n25670 vdd.n25669 4.5
R47514 vdd.n30553 vdd.n30552 4.5
R47515 vdd.n30575 vdd.n30574 4.5
R47516 vdd.n30277 vdd.n30276 4.5
R47517 vdd.n30247 vdd.n30246 4.5
R47518 vdd.n30254 vdd.n30253 4.5
R47519 vdd.n30201 vdd.n30200 4.5
R47520 vdd.n30194 vdd.n30193 4.5
R47521 vdd.n30692 vdd.n30691 4.5
R47522 vdd.n29713 vdd.n29712 4.5
R47523 vdd.n29767 vdd.n29766 4.5
R47524 vdd.n30012 vdd.n30011 4.5
R47525 vdd.n29828 vdd.n29827 4.5
R47526 vdd.n29846 vdd.n29845 4.5
R47527 vdd.n29946 vdd.n29945 4.5
R47528 vdd.n29861 vdd.n29860 4.5
R47529 vdd.n29882 vdd.n29881 4.5
R47530 vdd.n27917 vdd.n27916 4.5
R47531 vdd.n27940 vdd.n27939 4.5
R47532 vdd.n27802 vdd.n27801 4.5
R47533 vdd.n27822 vdd.n27821 4.5
R47534 vdd.n27815 vdd.n27814 4.5
R47535 vdd.n27753 vdd.n27752 4.5
R47536 vdd.n28976 vdd.n28975 4.5
R47537 vdd.n28067 vdd.n28066 4.5
R47538 vdd.n28072 vdd.n28071 4.5
R47539 vdd.n28125 vdd.n28124 4.5
R47540 vdd.n28817 vdd.n28816 4.5
R47541 vdd.n28803 vdd.n28181 4.5
R47542 vdd.n33838 vdd.n33837 4.5
R47543 vdd.n33850 vdd.n33849 4.5
R47544 vdd.n33787 vdd.n33786 4.5
R47545 vdd.n33778 vdd.n33777 4.5
R47546 vdd.n33708 vdd.n33707 4.5
R47547 vdd.n33715 vdd.n33714 4.5
R47548 vdd.n33725 vdd.n33724 4.5
R47549 vdd.n33736 vdd.n33735 4.5
R47550 vdd.n33744 vdd.n33743 4.5
R47551 vdd.n33671 vdd.n33670 4.5
R47552 vdd.n33684 vdd.n33683 4.5
R47553 vdd.n33695 vdd.n33694 4.5
R47554 vdd.n33481 vdd.n33480 4.5
R47555 vdd.n33490 vdd.n33489 4.5
R47556 vdd.n33501 vdd.n33500 4.5
R47557 vdd.n33523 vdd.n33522 4.5
R47558 vdd.n33347 vdd.n33346 4.5
R47559 vdd.n33360 vdd.n33359 4.5
R47560 vdd.n33371 vdd.n33370 4.5
R47561 vdd.n33469 vdd.n33468 4.5
R47562 vdd.n33451 vdd.n33450 4.5
R47563 vdd.n33400 vdd.n33399 4.5
R47564 vdd.n34193 vdd.n34192 4.5
R47565 vdd.n34207 vdd.n34206 4.5
R47566 vdd.n34219 vdd.n34218 4.5
R47567 vdd.n34230 vdd.n34229 4.5
R47568 vdd.n34081 vdd.n34080 4.5
R47569 vdd.n34088 vdd.n34087 4.5
R47570 vdd.n34097 vdd.n34096 4.5
R47571 vdd.n34106 vdd.n34105 4.5
R47572 vdd.n34122 vdd.n34121 4.5
R47573 vdd.n34309 vdd.n34308 4.5
R47574 vdd.n34322 vdd.n34321 4.5
R47575 vdd.n34337 vdd.n34336 4.5
R47576 vdd.n34350 vdd.n34349 4.5
R47577 vdd.n34363 vdd.n34362 4.5
R47578 vdd.n34376 vdd.n34375 4.5
R47579 vdd.n34388 vdd.n34387 4.5
R47580 vdd.n33910 vdd.n33909 4.5
R47581 vdd.n33898 vdd.n33897 4.5
R47582 vdd.n33956 vdd.n33955 4.5
R47583 vdd.n33884 vdd.n33883 4.5
R47584 vdd.n33870 vdd.n33869 4.5
R47585 vdd.n34060 vdd.n34059 4.5
R47586 vdd.n33982 vdd.n33981 4.5
R47587 vdd.n33991 vdd.n33990 4.5
R47588 vdd.n35303 vdd.n35302 4.5
R47589 vdd.n35291 vdd.n35290 4.5
R47590 vdd.n35339 vdd.n35338 4.5
R47591 vdd.n35351 vdd.n35350 4.5
R47592 vdd.n35240 vdd.n35239 4.5
R47593 vdd.n35249 vdd.n35248 4.5
R47594 vdd.n35258 vdd.n35257 4.5
R47595 vdd.n35485 vdd.n35484 4.5
R47596 vdd.n35509 vdd.n35508 4.5
R47597 vdd.n35575 vdd.n35574 4.5
R47598 vdd.n35588 vdd.n35587 4.5
R47599 vdd.n35603 vdd.n35602 4.5
R47600 vdd.n35368 vdd.n35367 4.5
R47601 vdd.n35379 vdd.n35378 4.5
R47602 vdd.n35399 vdd.n35398 4.5
R47603 vdd.n35407 vdd.n35406 4.5
R47604 vdd.n35079 vdd.n35078 4.5
R47605 vdd.n35092 vdd.n35091 4.5
R47606 vdd.n35042 vdd.n35041 4.5
R47607 vdd.n35109 vdd.n35108 4.5
R47608 vdd.n35121 vdd.n35120 4.5
R47609 vdd.n35221 vdd.n35220 4.5
R47610 vdd.n35144 vdd.n35143 4.5
R47611 vdd.n35153 vdd.n35152 4.5
R47612 vdd.n34719 vdd.n34718 4.5
R47613 vdd.n34707 vdd.n34706 4.5
R47614 vdd.n34755 vdd.n34754 4.5
R47615 vdd.n34767 vdd.n34766 4.5
R47616 vdd.n34653 vdd.n34652 4.5
R47617 vdd.n34662 vdd.n34661 4.5
R47618 vdd.n34674 vdd.n34673 4.5
R47619 vdd.n34957 vdd.n34956 4.5
R47620 vdd.n34976 vdd.n34975 4.5
R47621 vdd.n34904 vdd.n34903 4.5
R47622 vdd.n34894 vdd.n34893 4.5
R47623 vdd.n35015 vdd.n35014 4.5
R47624 vdd.n34778 vdd.n34777 4.5
R47625 vdd.n34789 vdd.n34788 4.5
R47626 vdd.n34802 vdd.n34801 4.5
R47627 vdd.n34811 vdd.n34810 4.5
R47628 vdd.n34492 vdd.n34491 4.5
R47629 vdd.n34505 vdd.n34504 4.5
R47630 vdd.n34458 vdd.n34457 4.5
R47631 vdd.n34522 vdd.n34521 4.5
R47632 vdd.n34534 vdd.n34533 4.5
R47633 vdd.n34634 vdd.n34633 4.5
R47634 vdd.n34557 vdd.n34556 4.5
R47635 vdd.n34568 vdd.n34567 4.5
R47636 vdd.n799 vdd.n798 4.5
R47637 vdd.n851 vdd.n850 4.5
R47638 vdd.n863 vdd.n862 4.5
R47639 vdd.n873 vdd.n872 4.5
R47640 vdd.n792 vdd.n791 4.5
R47641 vdd.n905 vdd.n904 4.5
R47642 vdd.n889 vdd.n888 4.5
R47643 vdd.n937 vdd.n936 4.5
R47644 vdd.n918 vdd.n917 4.5
R47645 vdd.n1064 vdd.n1063 4.5
R47646 vdd.n1149 vdd.n1148 4.5
R47647 vdd.n1161 vdd.n1160 4.5
R47648 vdd.n966 vdd.n965 4.5
R47649 vdd.n977 vdd.n976 4.5
R47650 vdd.n991 vdd.n990 4.5
R47651 vdd.n1004 vdd.n1003 4.5
R47652 vdd.n613 vdd.n612 4.5
R47653 vdd.n678 vdd.n677 4.5
R47654 vdd.n593 vdd.n592 4.5
R47655 vdd.n709 vdd.n708 4.5
R47656 vdd.n770 vdd.n769 4.5
R47657 vdd.n719 vdd.n718 4.5
R47658 vdd.n365 vdd.n364 4.5
R47659 vdd.n377 vdd.n376 4.5
R47660 vdd.n316 vdd.n315 4.5
R47661 vdd.n219 vdd.n218 4.5
R47662 vdd.n225 vdd.n224 4.5
R47663 vdd.n232 vdd.n231 4.5
R47664 vdd.n243 vdd.n242 4.5
R47665 vdd.n254 vdd.n253 4.5
R47666 vdd.n262 vdd.n261 4.5
R47667 vdd.n271 vdd.n270 4.5
R47668 vdd.n170 vdd.n169 4.5
R47669 vdd.n183 vdd.n182 4.5
R47670 vdd.n195 vdd.n194 4.5
R47671 vdd.n4 vdd.n3 4.5
R47672 vdd.n13 vdd.n12 4.5
R47673 vdd.n24 vdd.n23 4.5
R47674 vdd.n36 vdd.n35 4.5
R47675 vdd.n47 vdd.n46 4.5
R47676 vdd.n450 vdd.n449 4.5
R47677 vdd.n465 vdd.n464 4.5
R47678 vdd.n483 vdd.n482 4.5
R47679 vdd.n581 vdd.n580 4.5
R47680 vdd.n570 vdd.n569 4.5
R47681 vdd.n518 vdd.n517 4.5
R47682 vdd.n5894 vdd.n5893 4.5
R47683 vdd.n5908 vdd.n5907 4.5
R47684 vdd.n5920 vdd.n5919 4.5
R47685 vdd.n5857 vdd.n5856 4.5
R47686 vdd.n5783 vdd.n5782 4.5
R47687 vdd.n5790 vdd.n5789 4.5
R47688 vdd.n5802 vdd.n5801 4.5
R47689 vdd.n5814 vdd.n5813 4.5
R47690 vdd.n5989 vdd.n5988 4.5
R47691 vdd.n5947 vdd.n5946 4.5
R47692 vdd.n5937 vdd.n5936 4.5
R47693 vdd.n6038 vdd.n6037 4.5
R47694 vdd.n6056 vdd.n6055 4.5
R47695 vdd.n6069 vdd.n6068 4.5
R47696 vdd.n6090 vdd.n6089 4.5
R47697 vdd.n6101 vdd.n6100 4.5
R47698 vdd.n6184 vdd.n6183 4.5
R47699 vdd.n6172 vdd.n6171 4.5
R47700 vdd.n6240 vdd.n6239 4.5
R47701 vdd.n6158 vdd.n6157 4.5
R47702 vdd.n6144 vdd.n6143 4.5
R47703 vdd.n6345 vdd.n6344 4.5
R47704 vdd.n6267 vdd.n6266 4.5
R47705 vdd.n6279 vdd.n6278 4.5
R47706 vdd.n5466 vdd.n5465 4.5
R47707 vdd.n5454 vdd.n5453 4.5
R47708 vdd.n5502 vdd.n5501 4.5
R47709 vdd.n5514 vdd.n5513 4.5
R47710 vdd.n5400 vdd.n5399 4.5
R47711 vdd.n5409 vdd.n5408 4.5
R47712 vdd.n5421 vdd.n5420 4.5
R47713 vdd.n5704 vdd.n5703 4.5
R47714 vdd.n5723 vdd.n5722 4.5
R47715 vdd.n5651 vdd.n5650 4.5
R47716 vdd.n5641 vdd.n5640 4.5
R47717 vdd.n5762 vdd.n5761 4.5
R47718 vdd.n5525 vdd.n5524 4.5
R47719 vdd.n5536 vdd.n5535 4.5
R47720 vdd.n5549 vdd.n5548 4.5
R47721 vdd.n5558 vdd.n5557 4.5
R47722 vdd.n5239 vdd.n5238 4.5
R47723 vdd.n5252 vdd.n5251 4.5
R47724 vdd.n5205 vdd.n5204 4.5
R47725 vdd.n5269 vdd.n5268 4.5
R47726 vdd.n5281 vdd.n5280 4.5
R47727 vdd.n5381 vdd.n5380 4.5
R47728 vdd.n5304 vdd.n5303 4.5
R47729 vdd.n5315 vdd.n5314 4.5
R47730 vdd.n4898 vdd.n4897 4.5
R47731 vdd.n4888 vdd.n4887 4.5
R47732 vdd.n4933 vdd.n4932 4.5
R47733 vdd.n4945 vdd.n4944 4.5
R47734 vdd.n4805 vdd.n4804 4.5
R47735 vdd.n4814 vdd.n4813 4.5
R47736 vdd.n4825 vdd.n4824 4.5
R47737 vdd.n4833 vdd.n4832 4.5
R47738 vdd.n4843 vdd.n4842 4.5
R47739 vdd.n5081 vdd.n5080 4.5
R47740 vdd.n5148 vdd.n5147 4.5
R47741 vdd.n5161 vdd.n5160 4.5
R47742 vdd.n5175 vdd.n5174 4.5
R47743 vdd.n4956 vdd.n4955 4.5
R47744 vdd.n4967 vdd.n4966 4.5
R47745 vdd.n5046 vdd.n5045 4.5
R47746 vdd.n4980 vdd.n4979 4.5
R47747 vdd.n4989 vdd.n4988 4.5
R47748 vdd.n4752 vdd.n4751 4.5
R47749 vdd.n4765 vdd.n4764 4.5
R47750 vdd.n4782 vdd.n4781 4.5
R47751 vdd.n4794 vdd.n4793 4.5
R47752 vdd.n4702 vdd.n4701 4.5
R47753 vdd.n4628 vdd.n4627 4.5
R47754 vdd.n4635 vdd.n4634 4.5
R47755 vdd.n4293 vdd.n4292 4.5
R47756 vdd.n4281 vdd.n4280 4.5
R47757 vdd.n4329 vdd.n4328 4.5
R47758 vdd.n4341 vdd.n4340 4.5
R47759 vdd.n4230 vdd.n4229 4.5
R47760 vdd.n4239 vdd.n4238 4.5
R47761 vdd.n4251 vdd.n4250 4.5
R47762 vdd.n4531 vdd.n4530 4.5
R47763 vdd.n4553 vdd.n4552 4.5
R47764 vdd.n4478 vdd.n4477 4.5
R47765 vdd.n4468 vdd.n4467 4.5
R47766 vdd.n4592 vdd.n4591 4.5
R47767 vdd.n4352 vdd.n4351 4.5
R47768 vdd.n4363 vdd.n4362 4.5
R47769 vdd.n4376 vdd.n4375 4.5
R47770 vdd.n4384 vdd.n4383 4.5
R47771 vdd.n4069 vdd.n4068 4.5
R47772 vdd.n4082 vdd.n4081 4.5
R47773 vdd.n4035 vdd.n4034 4.5
R47774 vdd.n4099 vdd.n4098 4.5
R47775 vdd.n4111 vdd.n4110 4.5
R47776 vdd.n4211 vdd.n4210 4.5
R47777 vdd.n4134 vdd.n4133 4.5
R47778 vdd.n4146 vdd.n4145 4.5
R47779 vdd.n1880 vdd.n1879 4.5
R47780 vdd.n1180 vdd.n1179 4.5
R47781 vdd.n1911 vdd.n1910 4.5
R47782 vdd.n1204 vdd.n1203 4.5
R47783 vdd.n1934 vdd.n1933 4.5
R47784 vdd.n1187 vdd.n1186 4.5
R47785 vdd.n2068 vdd.n2067 4.5
R47786 vdd.n2673 vdd.n2672 4.5
R47787 vdd.n2004 vdd.n2003 4.5
R47788 vdd.n2576 vdd.n2575 4.5
R47789 vdd.n2533 vdd.n2532 4.5
R47790 vdd.n2424 vdd.n2423 4.5
R47791 vdd.n2407 vdd.n2406 4.5
R47792 vdd.n2386 vdd.n2385 4.5
R47793 vdd.n2045 vdd.n2044 4.5
R47794 vdd.n2031 vdd.n2030 4.5
R47795 vdd.n2116 vdd.n2115 4.5
R47796 vdd.n2141 vdd.n2140 4.5
R47797 vdd.n2024 vdd.n2023 4.5
R47798 vdd.n2126 vdd.n2125 4.5
R47799 vdd.n2162 vdd.n2161 4.5
R47800 vdd.n2145 vdd.n2144 4.5
R47801 vdd.n2184 vdd.n2183 4.5
R47802 vdd.n2201 vdd.n2200 4.5
R47803 vdd.n2019 vdd.n2018 4.5
R47804 vdd.n3760 vdd.n3759 4.5
R47805 vdd.n3745 vdd.n3744 4.5
R47806 vdd.n2683 vdd.n2682 4.5
R47807 vdd.n2691 vdd.n2690 4.5
R47808 vdd.n2678 vdd.n2677 4.5
R47809 vdd.n3729 vdd.n3728 4.5
R47810 vdd.n2704 vdd.n2703 4.5
R47811 vdd.n2727 vdd.n2726 4.5
R47812 vdd.n2060 vdd.n2059 4.5
R47813 vdd.n31288 vdd.n31280 4.5
R47814 vdd.n31042 vdd.n31041 4.5
R47815 vdd.n32452 vdd.n32451 4.5
R47816 vdd.n31518 vdd.n31517 4.5
R47817 vdd.n32274 vdd.n32273 4.5
R47818 vdd.n31553 vdd.n31552 4.5
R47819 vdd.n32183 vdd.n32182 4.5
R47820 vdd.n32132 vdd.n32131 4.5
R47821 vdd.n31587 vdd.n31586 4.5
R47822 vdd.n32074 vdd.n32073 4.5
R47823 vdd.n32103 vdd.n32102 4.5
R47824 vdd.n32161 vdd.n32160 4.5
R47825 vdd.n31561 vdd.n31560 4.5
R47826 vdd.n32240 vdd.n32239 4.5
R47827 vdd.n31543 vdd.n31542 4.5
R47828 vdd.n31537 vdd.n31536 4.5
R47829 vdd.n32293 vdd.n32292 4.5
R47830 vdd.n31528 vdd.n31527 4.5
R47831 vdd.n31069 vdd.n31068 4.5
R47832 vdd.n31032 vdd.n31031 4.5
R47833 vdd.n31022 vdd.n31021 4.5
R47834 vdd.n31025 vdd.n31024 4.5
R47835 vdd.n31286 vdd.n31285 4.5
R47836 vdd.n31924 vdd.n31923 4.5
R47837 vdd.n31690 vdd.n31689 4.5
R47838 vdd.n31705 vdd.n31704 4.5
R47839 vdd.n31727 vdd.n31726 4.5
R47840 vdd.n27214 vdd.n27213 4.5
R47841 vdd.n26154 vdd.n26153 4.5
R47842 vdd.n26396 vdd.n26395 4.5
R47843 vdd.n31739 vdd.n31738 4.5
R47844 vdd.n31780 vdd.n31779 4.5
R47845 vdd.n31716 vdd.n31715 4.5
R47846 vdd.n31684 vdd.n31683 4.5
R47847 vdd.n31929 vdd.n31928 4.5
R47848 vdd.n31948 vdd.n31947 4.5
R47849 vdd.n9260 vdd.n9253 4.5
R47850 vdd.n11622 vdd.n11621 4.5
R47851 vdd.n11606 vdd.n11605 4.5
R47852 vdd.n11609 vdd.n11580 4.5
R47853 vdd.n11619 vdd.n11618 4.5
R47854 vdd.n11618 vdd.n11617 4.5
R47855 vdd.n11612 vdd.n11610 4.5
R47856 vdd.n13140 vdd.n13139 4.5
R47857 vdd.n13141 vdd.n13140 4.5
R47858 vdd.n11593 vdd.n11592 4.5
R47859 vdd.n11595 vdd.n11594 4.5
R47860 vdd.n11604 vdd.n11603 4.5
R47861 vdd.n11591 vdd.n11588 4.5
R47862 vdd.n11939 vdd.n11557 4.5
R47863 vdd.n11939 vdd.n11938 4.5
R47864 vdd.n11951 vdd.n11950 4.5
R47865 vdd.n11556 vdd.n11555 4.5
R47866 vdd.n11538 vdd.n11452 4.5
R47867 vdd.n11538 vdd.n11537 4.5
R47868 vdd.n11541 vdd.n11450 4.5
R47869 vdd.n11953 vdd.n11952 4.5
R47870 vdd.n11954 vdd.n11953 4.5
R47871 vdd.n11515 vdd.n11514 4.5
R47872 vdd.n11516 vdd.n11515 4.5
R47873 vdd.n11513 vdd.n11462 4.5
R47874 vdd.n11532 vdd.n11456 4.5
R47875 vdd.n11532 vdd.n11531 4.5
R47876 vdd.n11508 vdd.n11502 4.5
R47877 vdd.n11511 vdd.n11460 4.5
R47878 vdd.n11460 vdd.n11458 4.5
R47879 vdd.n11498 vdd.n11463 4.5
R47880 vdd.n11501 vdd.n11435 4.5
R47881 vdd.n11497 vdd.n11496 4.5
R47882 vdd.n11492 vdd.n11491 4.5
R47883 vdd.n11495 vdd.n11494 4.5
R47884 vdd.n11470 vdd.n11468 4.5
R47885 vdd.n11490 vdd.n11467 4.5
R47886 vdd.n10197 vdd.n10196 4.5
R47887 vdd.n10203 vdd.n10202 4.5
R47888 vdd.n10210 vdd.n10209 4.5
R47889 vdd.n10215 vdd.n10214 4.5
R47890 vdd.n10220 vdd.n10219 4.5
R47891 vdd.n10250 vdd.n10128 4.5
R47892 vdd.n12580 vdd.n12579 4.5
R47893 vdd.n12573 vdd.n10258 4.5
R47894 vdd.n12572 vdd.n12571 4.5
R47895 vdd.n12572 vdd.n10260 4.5
R47896 vdd.n12574 vdd.n10267 4.5
R47897 vdd.n10267 vdd.n10258 4.5
R47898 vdd.n10254 vdd.n10127 4.5
R47899 vdd.n10252 vdd.n10251 4.5
R47900 vdd.n10216 vdd.n10070 4.5
R47901 vdd.n10211 vdd.n10076 4.5
R47902 vdd.n12579 vdd.n10253 4.5
R47903 vdd.n10129 vdd.n10128 4.5
R47904 vdd.n10222 vdd.n10221 4.5
R47905 vdd.n10220 vdd.n10217 4.5
R47906 vdd.n10215 vdd.n10212 4.5
R47907 vdd.n10210 vdd.n10207 4.5
R47908 vdd.n10203 vdd.n10200 4.5
R47909 vdd.n10204 vdd.n10079 4.5
R47910 vdd.n10079 vdd.n10065 4.5
R47911 vdd.n10197 vdd.n10136 4.5
R47912 vdd.n10194 vdd.n10087 4.5
R47913 vdd.n10197 vdd.n10085 4.5
R47914 vdd.n10203 vdd.n10089 4.5
R47915 vdd.n10210 vdd.n10077 4.5
R47916 vdd.n10215 vdd.n10095 4.5
R47917 vdd.n10220 vdd.n10071 4.5
R47918 vdd.n10221 vdd.n10134 4.5
R47919 vdd.n10131 vdd.n10128 4.5
R47920 vdd.n12579 vdd.n12578 4.5
R47921 vdd.n12575 vdd.n10258 4.5
R47922 vdd.n12575 vdd.n12574 4.5
R47923 vdd.n12574 vdd.n12573 4.5
R47924 vdd.n10178 vdd.n10083 4.5
R47925 vdd.n10178 vdd.n10084 4.5
R47926 vdd.n10181 vdd.n10180 4.5
R47927 vdd.n10184 vdd.n10082 4.5
R47928 vdd.n10180 vdd.n10143 4.5
R47929 vdd.n10177 vdd.n10053 4.5
R47930 vdd.n12618 vdd.n10053 4.5
R47931 vdd.n10173 vdd.n10144 4.5
R47932 vdd.n10173 vdd.n10050 4.5
R47933 vdd.n10176 vdd.n10052 4.5
R47934 vdd.n10166 vdd.n10165 4.5
R47935 vdd.n10169 vdd.n10168 4.5
R47936 vdd.n11762 vdd.n11678 4.5
R47937 vdd.n11759 vdd.n11680 4.5
R47938 vdd.n11695 vdd.n11683 4.5
R47939 vdd.n11755 vdd.n11685 4.5
R47940 vdd.n11756 vdd.n11755 4.5
R47941 vdd.n11748 vdd.n11720 4.5
R47942 vdd.n11750 vdd.n11719 4.5
R47943 vdd.n11747 vdd.n11721 4.5
R47944 vdd.n11724 vdd.n11721 4.5
R47945 vdd.n11775 vdd.n11774 4.5
R47946 vdd.n11677 vdd.n11676 4.5
R47947 vdd.n11769 vdd.n11768 4.5
R47948 vdd.n11768 vdd.n11670 4.5
R47949 vdd.n11686 vdd.n11683 4.5
R47950 vdd.n11873 vdd.n11805 4.5
R47951 vdd.n11892 vdd.n11796 4.5
R47952 vdd.n11894 vdd.n11893 4.5
R47953 vdd.n11802 vdd.n11801 4.5
R47954 vdd.n11879 vdd.n11878 4.5
R47955 vdd.n11887 vdd.n11886 4.5
R47956 vdd.n11886 vdd.n11885 4.5
R47957 vdd.n11889 vdd.n11888 4.5
R47958 vdd.n11812 vdd.n11811 4.5
R47959 vdd.n11812 vdd.n11807 4.5
R47960 vdd.n11820 vdd.n11819 4.5
R47961 vdd.n11867 vdd.n11809 4.5
R47962 vdd.n11868 vdd.n11867 4.5
R47963 vdd.n11897 vdd.n11794 4.5
R47964 vdd.n11903 vdd.n11902 4.5
R47965 vdd.n11915 vdd.n11787 4.5
R47966 vdd.n11907 vdd.n11663 4.5
R47967 vdd.n11909 vdd.n11787 4.5
R47968 vdd.n11911 vdd.n11663 4.5
R47969 vdd.n22466 vdd.n22465 4.5
R47970 vdd.n22451 vdd.n22450 4.5
R47971 vdd.n22436 vdd.n22435 4.5
R47972 vdd.n22421 vdd.n22420 4.5
R47973 vdd.n22406 vdd.n22405 4.5
R47974 vdd.n22382 vdd.n22381 4.5
R47975 vdd.n22349 vdd.n22348 4.5
R47976 vdd.n22213 vdd.n22212 4.5
R47977 vdd.n22229 vdd.n22228 4.5
R47978 vdd.n22255 vdd.n22254 4.5
R47979 vdd.n22322 vdd.n22321 4.5
R47980 vdd.n22307 vdd.n22306 4.5
R47981 vdd.n22292 vdd.n22291 4.5
R47982 vdd.n24366 vdd.n24365 4.5
R47983 vdd.n24351 vdd.n24350 4.5
R47984 vdd.n24327 vdd.n24326 4.5
R47985 vdd.n22065 vdd.n22064 4.5
R47986 vdd.n22077 vdd.n22076 4.5
R47987 vdd.n22105 vdd.n22104 4.5
R47988 vdd.n22131 vdd.n22130 4.5
R47989 vdd.n24294 vdd.n24293 4.5
R47990 vdd.n24279 vdd.n24278 4.5
R47991 vdd.n24264 vdd.n24263 4.5
R47992 vdd.n24249 vdd.n24248 4.5
R47993 vdd.n24234 vdd.n24233 4.5
R47994 vdd.n24210 vdd.n24209 4.5
R47995 vdd.n21628 vdd.n21627 4.5
R47996 vdd.n21651 vdd.n21650 4.5
R47997 vdd.n21682 vdd.n21681 4.5
R47998 vdd.n18403 vdd.n18402 4.5
R47999 vdd.n18376 vdd.n18375 4.5
R48000 vdd.n18382 vdd.n18381 4.5
R48001 vdd.n18356 vdd.n18355 4.5
R48002 vdd.n18369 vdd.n18368 4.5
R48003 vdd.n18348 vdd.n18347 4.5
R48004 vdd.n15122 vdd.n15121 4.5
R48005 vdd.n16702 vdd.n16701 4.5
R48006 vdd.n16730 vdd.n16729 4.5
R48007 vdd.n16717 vdd.n16716 4.5
R48008 vdd.n16752 vdd.n16751 4.5
R48009 vdd.n16762 vdd.n16761 4.5
R48010 vdd.n16582 vdd.n16581 4.5
R48011 vdd.n16768 vdd.n16767 4.5
R48012 vdd.n21769 vdd.n21768 4.5
R48013 vdd.n21853 vdd.n21848 4.5
R48014 vdd.n21964 vdd.n21896 4.5
R48015 vdd.n21983 vdd.n21887 4.5
R48016 vdd.n21985 vdd.n21984 4.5
R48017 vdd.n21893 vdd.n21892 4.5
R48018 vdd.n21970 vdd.n21969 4.5
R48019 vdd.n21978 vdd.n21977 4.5
R48020 vdd.n21977 vdd.n21976 4.5
R48021 vdd.n21980 vdd.n21979 4.5
R48022 vdd.n21903 vdd.n21902 4.5
R48023 vdd.n21903 vdd.n21898 4.5
R48024 vdd.n21911 vdd.n21910 4.5
R48025 vdd.n21958 vdd.n21900 4.5
R48026 vdd.n21959 vdd.n21958 4.5
R48027 vdd.n21988 vdd.n21885 4.5
R48028 vdd.n21994 vdd.n21993 4.5
R48029 vdd.n21755 vdd.n21754 4.5
R48030 vdd.n10357 vdd.n10344 4.493
R48031 vdd.n9442 vdd.n9435 4.493
R48032 vdd.n12985 vdd.n12984 4.493
R48033 vdd.n12974 vdd.n9454 4.493
R48034 vdd.n9608 vdd.n9571 4.493
R48035 vdd.n9630 vdd.n9615 4.493
R48036 vdd.n9648 vdd.n9647 4.493
R48037 vdd.t355 vdd.n12841 4.493
R48038 vdd.n9801 vdd.n9794 4.493
R48039 vdd.n12777 vdd.n12776 4.493
R48040 vdd.n12766 vdd.n9814 4.493
R48041 vdd.n9968 vdd.n9930 4.493
R48042 vdd.n9990 vdd.n9975 4.493
R48043 vdd.n10008 vdd.n10007 4.493
R48044 vdd.n10244 vdd.n10239 4.493
R48045 vdd.n10494 vdd.n10493 4.493
R48046 vdd.n12527 vdd.n10518 4.493
R48047 vdd.n12442 vdd.n12441 4.493
R48048 vdd.n12425 vdd.n10671 4.493
R48049 vdd.t310 vdd.n10774 4.493
R48050 vdd.n12341 vdd.n10817 4.493
R48051 vdd.n12324 vdd.n12323 4.493
R48052 vdd.n12242 vdd.n11003 4.493
R48053 vdd.n12224 vdd.n12223 4.493
R48054 vdd.n12144 vdd.n11146 4.493
R48055 vdd.n11210 vdd.n11209 4.493
R48056 vdd.n11273 vdd.t302 4.493
R48057 vdd.n12035 vdd.n11326 4.493
R48058 vdd.n12018 vdd.n12017 4.493
R48059 vdd.n11933 vdd.n11560 4.493
R48060 vdd.t370 vdd.n11560 4.493
R48061 vdd.n15426 vdd.n15425 4.493
R48062 vdd.n15659 vdd.n15658 4.493
R48063 vdd.n15679 vdd.n15678 4.493
R48064 vdd.n15695 vdd.n15694 4.493
R48065 vdd.n15915 vdd.n15914 4.493
R48066 vdd.n15935 vdd.n15934 4.493
R48067 vdd.n15951 vdd.n15950 4.493
R48068 vdd.t18 vdd.n16023 4.493
R48069 vdd.n16171 vdd.n16170 4.493
R48070 vdd.n16191 vdd.n16190 4.493
R48071 vdd.n16207 vdd.n16206 4.493
R48072 vdd.n16427 vdd.n16426 4.493
R48073 vdd.n16447 vdd.n16446 4.493
R48074 vdd.n16463 vdd.n16462 4.493
R48075 vdd.n16642 vdd.n16641 4.493
R48076 vdd.n15084 vdd.n15083 4.493
R48077 vdd.n16869 vdd.n16868 4.493
R48078 vdd.n17087 vdd.n17086 4.493
R48079 vdd.n17139 vdd.n17138 4.493
R48080 vdd.n17311 vdd.t270 4.493
R48081 vdd.n17359 vdd.n17358 4.493
R48082 vdd.n17411 vdd.n17410 4.493
R48083 vdd.n17617 vdd.n17616 4.493
R48084 vdd.n17669 vdd.n17668 4.493
R48085 vdd.n17888 vdd.n17887 4.493
R48086 vdd.n17940 vdd.n17939 4.493
R48087 vdd.n18063 vdd.t264 4.493
R48088 vdd.n18160 vdd.n18159 4.493
R48089 vdd.n18212 vdd.n18211 4.493
R48090 vdd.n15015 vdd.n15011 4.493
R48091 vdd.t27 vdd.n15015 4.493
R48092 vdd.n12600 vdd.n10072 4.479
R48093 vdd.n16743 vdd.n16597 4.479
R48094 vdd.n13133 vdd.n9263 4.478
R48095 vdd.n13205 vdd.n13204 4.478
R48096 vdd.n38184 vdd.n37596 4.47
R48097 vdd.n37432 vdd.n37431 4.47
R48098 vdd.n33106 vdd.n33102 4.47
R48099 vdd.n37048 vdd.n37045 4.47
R48100 vdd.n37030 vdd.n35676 4.47
R48101 vdd.n33099 vdd.n33090 4.47
R48102 vdd.n37411 vdd.n37391 4.47
R48103 vdd.n38184 vdd.n37595 4.47
R48104 vdd.n37432 vdd.n37426 4.47
R48105 vdd.n37411 vdd.n37400 4.47
R48106 vdd.n33099 vdd.n33094 4.47
R48107 vdd.n33106 vdd.n33101 4.47
R48108 vdd.n37048 vdd.n37043 4.47
R48109 vdd.n37030 vdd.n35675 4.47
R48110 vdd.n33150 vdd.n33149 4.47
R48111 vdd.n35644 vdd.n35643 4.47
R48112 vdd.n37328 vdd.n37325 4.47
R48113 vdd.n37364 vdd.n37355 4.47
R48114 vdd.n35673 vdd.n35670 4.47
R48115 vdd.n32835 vdd.n32832 4.47
R48116 vdd.n28833 vdd.n28820 4.47
R48117 vdd.n28029 vdd.n27781 4.47
R48118 vdd.n28022 vdd.n28021 4.47
R48119 vdd.n29783 vdd.n29699 4.47
R48120 vdd.n29773 vdd.n29772 4.47
R48121 vdd.n29773 vdd.n29700 4.47
R48122 vdd.n29783 vdd.n29698 4.47
R48123 vdd.n28022 vdd.n27825 4.47
R48124 vdd.n28029 vdd.n27780 4.47
R48125 vdd.n28833 vdd.n28819 4.47
R48126 vdd.n30536 vdd.n30320 4.47
R48127 vdd.n30510 vdd.n30322 4.47
R48128 vdd.n30536 vdd.n30319 4.47
R48129 vdd.n25535 vdd.n25534 4.47
R48130 vdd.n25584 vdd.n25583 4.47
R48131 vdd.n3684 vdd.n2708 4.47
R48132 vdd.n2248 vdd.n2204 4.47
R48133 vdd.n2261 vdd.n2166 4.47
R48134 vdd.n2631 vdd.n2586 4.47
R48135 vdd.n2661 vdd.n2571 4.47
R48136 vdd.n3684 vdd.n2706 4.47
R48137 vdd.n2248 vdd.n2203 4.47
R48138 vdd.n2261 vdd.n2164 4.47
R48139 vdd.n2631 vdd.n2585 4.47
R48140 vdd.n2661 vdd.n2569 4.47
R48141 vdd.n26155 vdd.n26150 4.47
R48142 vdd.n31916 vdd.n31677 4.47
R48143 vdd.n32288 vdd.n31531 4.47
R48144 vdd.n31959 vdd.n31662 4.47
R48145 vdd.n32315 vdd.n31502 4.47
R48146 vdd.n26155 vdd.n26148 4.47
R48147 vdd.n31916 vdd.n31676 4.47
R48148 vdd.n31959 vdd.n31957 4.47
R48149 vdd.n32288 vdd.n31530 4.47
R48150 vdd.n32315 vdd.n32313 4.47
R48151 vdd.n13371 vdd.n9065 4.47
R48152 vdd.n13400 vdd.n9050 4.47
R48153 vdd.n13663 vdd.n8845 4.47
R48154 vdd.n13693 vdd.n8829 4.47
R48155 vdd.n8667 vdd.n8662 4.47
R48156 vdd.n8609 vdd.n8608 4.47
R48157 vdd.n8444 vdd.n8441 4.47
R48158 vdd.n8387 vdd.n8386 4.47
R48159 vdd.n14708 vdd.n8115 4.47
R48160 vdd.n8117 vdd.n8116 4.47
R48161 vdd.n14854 vdd.n8027 4.47
R48162 vdd.n14881 vdd.n8026 4.47
R48163 vdd.n20149 vdd.n20015 4.47
R48164 vdd.n20156 vdd.n20014 4.47
R48165 vdd.n20385 vdd.n19989 4.47
R48166 vdd.n20392 vdd.n19988 4.47
R48167 vdd.n20729 vdd.n19936 4.47
R48168 vdd.n20736 vdd.n19924 4.47
R48169 vdd.n20918 vdd.n19868 4.47
R48170 vdd.n20925 vdd.n19856 4.47
R48171 vdd.n19728 vdd.n19202 4.47
R48172 vdd.n19721 vdd.n19214 4.47
R48173 vdd.n19527 vdd.n19258 4.47
R48174 vdd.n19520 vdd.n19270 4.47
R48175 vdd.n25161 vdd.n24986 4.47
R48176 vdd.n25166 vdd.n24985 4.47
R48177 vdd.n24750 vdd.n24516 4.47
R48178 vdd.n24745 vdd.n24517 4.47
R48179 vdd.n2529 vdd.n2528 4.447
R48180 vdd.n1846 vdd.n1242 4.447
R48181 vdd.n3866 vdd.n3821 4.447
R48182 vdd.n31157 vdd.n31156 4.444
R48183 vdd.n32044 vdd.n31600 4.398
R48184 vdd.n26317 vdd.n26313 4.398
R48185 vdd.n32368 vdd.n31463 4.398
R48186 vdd.n259 vdd.n258 4.384
R48187 vdd.n37537 vdd.n37536 4.384
R48188 vdd.n33003 vdd.n33002 4.384
R48189 vdd.n37293 vdd.n37287 4.384
R48190 vdd.n37153 vdd.n37141 4.384
R48191 vdd.n33188 vdd.n33187 4.384
R48192 vdd.n32878 vdd.n32860 4.384
R48193 vdd.n37537 vdd.n37530 4.384
R48194 vdd.n32878 vdd.n32875 4.384
R48195 vdd.n33003 vdd.n32996 4.384
R48196 vdd.n37293 vdd.n37286 4.384
R48197 vdd.n37153 vdd.n37133 4.384
R48198 vdd.n33188 vdd.n33186 4.384
R48199 vdd.n37472 vdd.n37461 4.384
R48200 vdd.n32931 vdd.n32920 4.384
R48201 vdd.n37099 vdd.n37077 4.384
R48202 vdd.n33258 vdd.n33257 4.384
R48203 vdd.n37230 vdd.n37222 4.384
R48204 vdd.n33064 vdd.n33042 4.384
R48205 vdd.n30550 vdd.n30316 4.384
R48206 vdd.n25552 vdd.n25551 4.384
R48207 vdd.n25568 vdd.n25563 4.384
R48208 vdd.n13503 vdd.n8984 4.384
R48209 vdd.n13542 vdd.n13541 4.384
R48210 vdd.n13783 vdd.n8769 4.384
R48211 vdd.n13827 vdd.n13826 4.384
R48212 vdd.n8555 vdd.n8517 4.384
R48213 vdd.n8520 vdd.n8519 4.384
R48214 vdd.n20817 vdd.n19898 4.384
R48215 vdd.n20847 vdd.n19893 4.384
R48216 vdd.n19831 vdd.n19161 4.384
R48217 vdd.n19811 vdd.n19177 4.384
R48218 vdd.n19639 vdd.n19228 4.384
R48219 vdd.n19609 vdd.n19233 4.384
R48220 ldomc_0.otaldom_0.pcsm_0.vdd vdd.n13784 4.332
R48221 bandgapmd_0.otam_1.pcsm_0.vdd vdd.n19828 4.332
R48222 vdd.n9100 vdd.n9099 4.332
R48223 vdd.n13418 vdd.n13417 4.332
R48224 vdd.n13565 vdd.n8940 4.332
R48225 vdd.n13690 vdd.n8831 4.332
R48226 vdd.n8670 vdd.n8661 4.332
R48227 vdd.n14044 vdd.n14043 4.332
R48228 vdd.n14182 vdd.n8464 4.332
R48229 vdd.n8353 vdd.n8352 4.332
R48230 vdd.n19500 vdd.n19283 4.332
R48231 vdd.n19562 vdd.n19234 4.332
R48232 vdd.n19667 vdd.n19227 4.332
R48233 vdd.n19731 vdd.n19190 4.332
R48234 vdd.n20928 vdd.n19844 4.332
R48235 vdd.n20864 vdd.n19881 4.332
R48236 vdd.n20770 vdd.n19899 4.332
R48237 vdd.n20709 vdd.n19949 4.332
R48238 vdd.n10 vdd.n9 4.328
R48239 vdd.n33494 vdd.n33493 4.326
R48240 vdd.n984 vdd.n983 4.326
R48241 vdd.n25542 vdd.n25541 4.326
R48242 vdd.n30311 vdd.n30310 4.326
R48243 vdd.n2130 vdd.n2129 4.326
R48244 vdd.n38198 vdd.n37592 4.302
R48245 vdd.n32936 vdd.n32935 4.302
R48246 vdd.n32952 vdd.n32948 4.302
R48247 vdd.n37238 vdd.n37237 4.302
R48248 vdd.n37193 vdd.n37192 4.302
R48249 vdd.n37015 vdd.n35680 4.302
R48250 vdd.n33272 vdd.n33256 4.302
R48251 vdd.n38198 vdd.n37590 4.302
R48252 vdd.n32936 vdd.n32933 4.302
R48253 vdd.n32952 vdd.n32946 4.302
R48254 vdd.n37238 vdd.n37232 4.302
R48255 vdd.n37193 vdd.n37190 4.302
R48256 vdd.n37015 vdd.n35678 4.302
R48257 vdd.n33272 vdd.n33254 4.302
R48258 vdd.n36987 vdd.n35687 4.302
R48259 vdd.n37152 vdd.n37151 4.302
R48260 vdd.n37188 vdd.n37179 4.302
R48261 vdd.n32995 vdd.n32992 4.302
R48262 vdd.n32981 vdd.n32978 4.302
R48263 vdd.n37529 vdd.n37526 4.302
R48264 vdd.n37573 vdd.n37572 4.302
R48265 vdd.n29725 vdd.n29724 4.302
R48266 vdd.n30557 vdd.n30556 4.302
R48267 vdd.n30557 vdd.n30314 4.302
R48268 vdd.n25513 vdd.n25509 4.302
R48269 vdd.n25615 vdd.n25424 4.302
R48270 vdd.n9098 vdd.n9066 4.302
R48271 vdd.n13397 vdd.n13394 4.302
R48272 vdd.n8878 vdd.n8846 4.302
R48273 vdd.n13689 vdd.n13686 4.302
R48274 vdd.n13912 vdd.n8671 4.302
R48275 vdd.n13983 vdd.n8607 4.302
R48276 vdd.n14202 vdd.n8447 4.302
R48277 vdd.n14273 vdd.n8385 4.302
R48278 vdd.n20726 vdd.n19948 4.302
R48279 vdd.n20739 vdd.n19912 4.302
R48280 vdd.n20915 vdd.n19880 4.302
R48281 vdd.n20929 vdd.n19843 4.302
R48282 vdd.n19732 vdd.n19189 4.302
R48283 vdd.n19718 vdd.n19226 4.302
R48284 vdd.n19530 vdd.n19246 4.302
R48285 vdd.n19517 vdd.n19282 4.302
R48286 vdd.t120 vdd.n13365 4.282
R48287 vdd.n13428 vdd.n13427 4.282
R48288 vdd.n13499 vdd.n13498 4.282
R48289 vdd.n13720 vdd.n13719 4.282
R48290 vdd.n14012 vdd.n14011 4.282
R48291 vdd.n14078 vdd.n8552 4.282
R48292 vdd.n14302 vdd.n14301 4.282
R48293 vdd.n14548 vdd.n14547 4.282
R48294 vdd.n32395 vdd.n32394 4.266
R48295 vdd.n29822 vdd.n29821 4.261
R48296 vdd.n25466 vdd.n25465 4.223
R48297 vdd.n25422 vdd.n25416 4.223
R48298 vdd.n21560 vdd.n21559 4.222
R48299 vdd.n21478 vdd.n21477 4.222
R48300 vdd.n21301 vdd.n21300 4.222
R48301 vdd.n21219 vdd.n21218 4.222
R48302 vdd.n21042 vdd.n21041 4.222
R48303 vdd.t347 vdd.n19124 4.222
R48304 vdd.n19112 vdd.n19111 4.222
R48305 vdd.n18935 vdd.n18934 4.222
R48306 vdd.n18853 vdd.n18852 4.222
R48307 vdd.n18676 vdd.n18675 4.222
R48308 vdd.n18594 vdd.n18593 4.222
R48309 vdd.n10465 vdd.n10279 4.194
R48310 vdd.n10431 vdd.n10430 4.194
R48311 vdd.n15287 vdd.n15286 4.194
R48312 vdd.n15338 vdd.n15337 4.194
R48313 vdd.n13050 vdd.n9317 4.172
R48314 vdd.n13030 vdd.n9355 4.172
R48315 vdd.n9368 vdd.n9355 4.172
R48316 vdd.n12949 vdd.n9475 4.172
R48317 vdd.n12929 vdd.n12928 4.172
R48318 vdd.n12928 vdd.n9525 4.172
R48319 vdd.n12842 vdd.n9679 4.172
R48320 vdd.n12822 vdd.n9715 4.172
R48321 vdd.n9728 vdd.n9715 4.172
R48322 vdd.n12741 vdd.n9835 4.172
R48323 vdd.n12721 vdd.n12720 4.172
R48324 vdd.n12720 vdd.n9886 4.172
R48325 vdd.n12634 vdd.n10039 4.172
R48326 vdd.n12613 vdd.n10057 4.172
R48327 vdd.n10139 vdd.n10057 4.172
R48328 vdd.n10577 vdd.n10573 4.172
R48329 vdd.n12472 vdd.n12471 4.172
R48330 vdd.n12394 vdd.n10720 4.172
R48331 vdd.n12371 vdd.n12370 4.172
R48332 vdd.n12292 vdd.n10906 4.172
R48333 vdd.n12277 vdd.n10922 4.172
R48334 vdd.n12192 vdd.n12191 4.172
R48335 vdd.n12173 vdd.n11105 4.172
R48336 vdd.n11260 vdd.n11259 4.172
R48337 vdd.n12065 vdd.n12064 4.172
R48338 vdd.n11986 vdd.n11414 4.172
R48339 vdd.n11971 vdd.n11431 4.172
R48340 vdd.n15512 vdd.n15508 4.172
R48341 vdd.n15575 vdd.n15572 4.172
R48342 vdd.n15575 vdd.n15574 4.172
R48343 vdd.n15768 vdd.n15764 4.172
R48344 vdd.n15831 vdd.n15828 4.172
R48345 vdd.n15831 vdd.n15830 4.172
R48346 vdd.n16024 vdd.n16020 4.172
R48347 vdd.n16087 vdd.n16084 4.172
R48348 vdd.n16087 vdd.n16086 4.172
R48349 vdd.n16280 vdd.n16276 4.172
R48350 vdd.n16343 vdd.n16340 4.172
R48351 vdd.n16343 vdd.n16342 4.172
R48352 vdd.n16536 vdd.n16532 4.172
R48353 vdd.n16554 vdd.n16552 4.172
R48354 vdd.n16552 vdd.n16550 4.172
R48355 vdd.n16946 vdd.n16943 4.172
R48356 vdd.n17006 vdd.n17003 4.172
R48357 vdd.n17218 vdd.n17215 4.172
R48358 vdd.n17278 vdd.n17275 4.172
R48359 vdd.n17490 vdd.n17487 4.172
R48360 vdd.n17550 vdd.n17547 4.172
R48361 vdd.n17748 vdd.n17745 4.172
R48362 vdd.n17808 vdd.n17805 4.172
R48363 vdd.n18019 vdd.n18016 4.172
R48364 vdd.n18079 vdd.n18076 4.172
R48365 vdd.n18286 vdd.n18284 4.172
R48366 vdd.n18326 vdd.n18324 4.172
R48367 vdd.n15353 vdd.n15350 4.163
R48368 vdd.n12 vdd.n10 4.162
R48369 vdd.n33500 vdd.n33498 4.154
R48370 vdd.n34362 vdd.n34360 4.154
R48371 vdd.n35378 vdd.n35376 4.154
R48372 vdd.n34788 vdd.n34786 4.154
R48373 vdd.n990 vdd.n988 4.154
R48374 vdd.n6068 vdd.n6066 4.154
R48375 vdd.n5535 vdd.n5533 4.154
R48376 vdd.n4781 vdd.n4780 4.154
R48377 vdd.n4362 vdd.n4360 4.154
R48378 vdd.n27474 vdd.n27472 4.154
R48379 vdd.n11884 vdd.n11883 4.145
R48380 vdd.n21975 vdd.n21974 4.145
R48381 vdd.n31536 vdd.n31535 4.141
R48382 vdd.n31536 vdd.n31533 4.141
R48383 vdd.n31552 vdd.n31551 4.141
R48384 vdd.n31560 vdd.n31558 4.141
R48385 vdd.n31558 vdd.n31557 4.141
R48386 vdd.n31931 vdd.n31930 4.141
R48387 vdd.n31038 vdd.n31037 4.141
R48388 vdd.n31143 vdd.n31142 4.141
R48389 vdd.n30344 vdd.n30343 4.141
R48390 vdd.n35708 vdd.n35707 4.141
R48391 vdd.n35997 vdd.n35996 4.141
R48392 vdd.n36067 vdd.n36066 4.141
R48393 vdd.n36228 vdd.n36227 4.141
R48394 vdd.n36298 vdd.n36297 4.141
R48395 vdd.n36459 vdd.n36458 4.141
R48396 vdd.n36529 vdd.n36528 4.141
R48397 vdd.n36690 vdd.n36689 4.141
R48398 vdd.n36760 vdd.n36759 4.141
R48399 vdd.n36921 vdd.n36920 4.141
R48400 vdd.n37002 vdd.n37001 4.141
R48401 vdd.n33168 vdd.n33167 4.141
R48402 vdd.n33130 vdd.n33129 4.141
R48403 vdd.n37309 vdd.n37308 4.141
R48404 vdd.n37381 vdd.n37380 4.141
R48405 vdd.n32842 vdd.n32841 4.141
R48406 vdd.n38206 vdd.n38205 4.141
R48407 vdd.n38046 vdd.n38045 4.141
R48408 vdd.n37976 vdd.n37975 4.141
R48409 vdd.n37815 vdd.n37814 4.141
R48410 vdd.n37745 vdd.n37744 4.141
R48411 vdd.n28187 vdd.n28186 4.141
R48412 vdd.n28257 vdd.n28256 4.141
R48413 vdd.n28418 vdd.n28417 4.141
R48414 vdd.n28488 vdd.n28487 4.141
R48415 vdd.n28649 vdd.n28648 4.141
R48416 vdd.n28719 vdd.n28718 4.141
R48417 vdd.n27832 vdd.n27831 4.141
R48418 vdd.n27907 vdd.n27906 4.141
R48419 vdd.n30193 vdd.n30184 4.141
R48420 vdd.n25457 vdd.n25455 4.141
R48421 vdd.n25412 vdd.n25411 4.141
R48422 vdd.n1677 vdd.n1676 4.141
R48423 vdd.n1623 vdd.n1622 4.141
R48424 vdd.n1496 vdd.n1495 4.141
R48425 vdd.n1442 vdd.n1441 4.141
R48426 vdd.n1315 vdd.n1314 4.141
R48427 vdd.n26781 vdd.n26780 4.141
R48428 vdd.n26908 vdd.n26907 4.141
R48429 vdd.n26962 vdd.n26961 4.141
R48430 vdd.n27089 vdd.n27088 4.141
R48431 vdd.n27143 vdd.n27142 4.141
R48432 vdd.n1185 vdd.n1184 4.141
R48433 vdd.n1186 vdd.n1185 4.141
R48434 vdd.n2667 vdd.n2666 4.141
R48435 vdd.n2396 vdd.n2395 4.141
R48436 vdd.n2114 vdd.n2113 4.141
R48437 vdd.n2159 vdd.n2151 4.141
R48438 vdd.n3743 vdd.n3742 4.141
R48439 vdd.n2700 vdd.n2699 4.141
R48440 vdd.n2737 vdd.n2736 4.141
R48441 vdd.n2861 vdd.n2860 4.141
R48442 vdd.n2915 vdd.n2914 4.141
R48443 vdd.n3042 vdd.n3041 4.141
R48444 vdd.n3096 vdd.n3095 4.141
R48445 vdd.n3223 vdd.n3222 4.141
R48446 vdd.n3277 vdd.n3276 4.141
R48447 vdd.n3404 vdd.n3403 4.141
R48448 vdd.n3458 vdd.n3457 4.141
R48449 vdd.n3585 vdd.n3584 4.141
R48450 vdd.n3648 vdd.n3647 4.141
R48451 vdd.n31738 vdd.n31737 4.141
R48452 vdd.n31702 vdd.n31701 4.141
R48453 vdd.n31704 vdd.n31702 4.141
R48454 vdd.n13120 vdd.n9271 4.141
R48455 vdd.n13122 vdd.n9267 4.141
R48456 vdd.n13340 vdd.n13339 4.141
R48457 vdd.n13346 vdd.n13345 4.141
R48458 vdd.n13412 vdd.n9040 4.141
R48459 vdd.n13414 vdd.n9036 4.141
R48460 vdd.n13632 vdd.n13631 4.141
R48461 vdd.n13638 vdd.n13637 4.141
R48462 vdd.n13706 vdd.n8819 4.141
R48463 vdd.n13708 vdd.n8815 4.141
R48464 vdd.n8689 vdd.n8674 4.141
R48465 vdd.n8675 vdd.n8672 4.141
R48466 vdd.n13990 vdd.n13989 4.141
R48467 vdd.n8606 vdd.n8605 4.141
R48468 vdd.n8466 vdd.n8450 4.141
R48469 vdd.n8451 vdd.n8448 4.141
R48470 vdd.n14281 vdd.n14280 4.141
R48471 vdd.n8384 vdd.n8383 4.141
R48472 vdd.n14491 vdd.n8218 4.141
R48473 vdd.n14498 vdd.n14497 4.141
R48474 vdd.n14676 vdd.n8131 4.141
R48475 vdd.n14677 vdd.n14676 4.141
R48476 vdd.n14733 vdd.n8109 4.141
R48477 vdd.n14733 vdd.n14722 4.141
R48478 vdd.n14848 vdd.n8041 4.141
R48479 vdd.n14849 vdd.n14848 4.141
R48480 vdd.n14890 vdd.n14887 4.141
R48481 vdd.n14887 vdd.n8014 4.141
R48482 vdd.n13174 vdd.n9228 4.141
R48483 vdd.n13227 vdd.n13226 4.141
R48484 vdd.n13314 vdd.n9134 4.141
R48485 vdd.n9135 vdd.n9108 4.141
R48486 vdd.n13467 vdd.n13466 4.141
R48487 vdd.n13519 vdd.n13518 4.141
R48488 vdd.n13606 vdd.n8912 4.141
R48489 vdd.n8913 vdd.n8887 4.141
R48490 vdd.n13799 vdd.n8758 4.141
R48491 vdd.n8763 vdd.n8762 4.141
R48492 vdd.n13881 vdd.n8697 4.141
R48493 vdd.n8699 vdd.n8698 4.141
R48494 vdd.n14086 vdd.n8545 4.141
R48495 vdd.n8550 vdd.n8549 4.141
R48496 vdd.n14170 vdd.n8474 4.141
R48497 vdd.n8476 vdd.n8475 4.141
R48498 vdd.n8330 vdd.n8329 4.141
R48499 vdd.n14384 vdd.n14383 4.141
R48500 vdd.n14470 vdd.n8230 4.141
R48501 vdd.n14472 vdd.n8227 4.141
R48502 vdd.n24231 vdd.n24224 4.141
R48503 vdd.n24233 vdd.n24231 4.141
R48504 vdd.n24131 vdd.n24124 4.141
R48505 vdd.n24049 vdd.n24042 4.141
R48506 vdd.n23899 vdd.n23892 4.141
R48507 vdd.n23817 vdd.n23810 4.141
R48508 vdd.n23667 vdd.n23660 4.141
R48509 vdd.n23129 vdd.n23122 4.141
R48510 vdd.n23211 vdd.n23204 4.141
R48511 vdd.n23361 vdd.n23354 4.141
R48512 vdd.n23443 vdd.n23436 4.141
R48513 vdd.n23593 vdd.n23586 4.141
R48514 vdd.n22550 vdd.n22543 4.141
R48515 vdd.n22632 vdd.n22625 4.141
R48516 vdd.n22782 vdd.n22775 4.141
R48517 vdd.n22864 vdd.n22857 4.141
R48518 vdd.n23014 vdd.n23007 4.141
R48519 vdd.n22403 vdd.n22396 4.141
R48520 vdd.n22405 vdd.n22403 4.141
R48521 vdd.n24348 vdd.n24341 4.141
R48522 vdd.n24350 vdd.n24348 4.141
R48523 vdd.n19301 vdd.n19300 4.141
R48524 vdd.n19504 vdd.n19503 4.141
R48525 vdd.n19534 vdd.n19533 4.141
R48526 vdd.n19705 vdd.n19704 4.141
R48527 vdd.n19736 vdd.n19735 4.141
R48528 vdd.n20933 vdd.n20932 4.141
R48529 vdd.n20902 vdd.n20901 4.141
R48530 vdd.n20743 vdd.n20742 4.141
R48531 vdd.n20713 vdd.n20712 4.141
R48532 vdd.n19971 vdd.n19970 4.141
R48533 vdd.n21553 vdd.n21552 4.141
R48534 vdd.n21471 vdd.n21470 4.141
R48535 vdd.n21294 vdd.n21293 4.141
R48536 vdd.n21212 vdd.n21211 4.141
R48537 vdd.n21035 vdd.n21034 4.141
R48538 vdd.n19105 vdd.n19104 4.141
R48539 vdd.n18928 vdd.n18927 4.141
R48540 vdd.n18846 vdd.n18845 4.141
R48541 vdd.n18669 vdd.n18668 4.141
R48542 vdd.n18587 vdd.n18586 4.141
R48543 vdd.n20438 vdd.n20429 4.141
R48544 vdd.n20348 vdd.n20339 4.141
R48545 vdd.n20202 vdd.n20193 4.141
R48546 vdd.n20112 vdd.n20103 4.141
R48547 vdd.n24716 vdd.n24711 4.141
R48548 vdd.n24781 vdd.n24776 4.141
R48549 vdd.n25199 vdd.n25194 4.141
R48550 vdd.n25134 vdd.n25129 4.141
R48551 vdd.n27933 vdd.n27929 4.14
R48552 vdd.n11780 vdd.n11778 4.139
R48553 vdd.n21871 vdd.n21870 4.139
R48554 vdd.n32510 vdd.n32508 4.106
R48555 vdd.n19366 vdd.n19363 4.104
R48556 vdd.n19480 vdd.t152 4.104
R48557 vdd.n19479 vdd.n19476 4.104
R48558 vdd.n19572 vdd.n19569 4.104
R48559 vdd.n19679 vdd.n19676 4.104
R48560 vdd.n19774 vdd.n19771 4.104
R48561 vdd.t168 vdd.n19806 4.104
R48562 vdd.n19807 vdd.t168 4.104
R48563 vdd.n20999 vdd.t160 4.104
R48564 vdd.t160 vdd.n19156 4.104
R48565 vdd.n20971 vdd.n20968 4.104
R48566 vdd.n20876 vdd.n20873 4.104
R48567 vdd.n20780 vdd.n20777 4.104
R48568 vdd.n20688 vdd.n20685 4.104
R48569 vdd.n20689 vdd.t156 4.104
R48570 vdd.n20575 vdd.n20572 4.104
R48571 vdd.n19977 vdd.n19976 4.104
R48572 vdd.n20314 vdd.n20313 4.104
R48573 vdd.n20232 vdd.n20231 4.104
R48574 vdd.n20078 vdd.n20077 4.104
R48575 vdd.n14759 vdd.n14758 4.094
R48576 vdd.n14817 vdd.n14816 4.094
R48577 vdd.n14932 vdd.n14931 4.094
R48578 vdd.n10600 vdd.n10591 4.029
R48579 vdd.n10686 vdd.n10680 4.029
R48580 vdd.n10759 vdd.n10751 4.029
R48581 vdd.n12332 vdd.n10829 4.029
R48582 vdd.n12283 vdd.n10919 4.029
R48583 vdd.n11031 vdd.n11015 4.029
R48584 vdd.n12181 vdd.n11092 4.029
R48585 vdd.n12125 vdd.n12124 4.029
R48586 vdd.n12076 vdd.n11268 4.029
R48587 vdd.n12026 vdd.n11338 4.029
R48588 vdd.n11977 vdd.n11428 4.029
R48589 vdd.n11602 vdd.n11598 4.029
R48590 vdd.n16978 vdd.n16971 4.029
R48591 vdd.n17126 vdd.n17125 4.029
R48592 vdd.n17250 vdd.n17243 4.029
R48593 vdd.n17398 vdd.n17397 4.029
R48594 vdd.n17522 vdd.n17515 4.029
R48595 vdd.n17656 vdd.n17655 4.029
R48596 vdd.n17780 vdd.n17773 4.029
R48597 vdd.n17927 vdd.n17926 4.029
R48598 vdd.n18051 vdd.n18044 4.029
R48599 vdd.n18199 vdd.n18198 4.029
R48600 vdd.n16817 vdd.n16811 4.029
R48601 vdd.n21702 vdd.n15018 4.029
R48602 vdd.n3900 vdd.n3899 4.015
R48603 vdd.n11603 vdd.n11602 4
R48604 vdd.n21702 vdd.n21701 4
R48605 vdd.n11674 vdd.n11673 3.983
R48606 vdd.n21850 vdd.n21849 3.983
R48607 vdd.n38155 vdd.n38154 3.98
R48608 vdd.n13366 vdd.n9070 3.976
R48609 vdd.n13578 vdd.n8930 3.976
R48610 vdd.n13658 vdd.n8850 3.976
R48611 vdd.n8664 vdd.n8663 3.976
R48612 vdd.n14160 vdd.n14159 3.976
R48613 vdd.n8438 vdd.n8420 3.976
R48614 vdd.n14277 vdd.t287 3.976
R48615 vdd.n14440 vdd.n14439 3.976
R48616 vdd.n33487 vdd.n33486 3.951
R48617 vdd.n974 vdd.n973 3.951
R48618 vdd.n4821 vdd.n4820 3.95
R48619 vdd.n25491 vdd.n25490 3.95
R48620 vdd.n36031 vdd.n36027 3.931
R48621 vdd.n36045 vdd.n36041 3.931
R48622 vdd.n36262 vdd.n36258 3.931
R48623 vdd.n36276 vdd.n36272 3.931
R48624 vdd.n36493 vdd.n36489 3.931
R48625 vdd.n36507 vdd.n36503 3.931
R48626 vdd.n36724 vdd.n36720 3.931
R48627 vdd.n36738 vdd.n36734 3.931
R48628 vdd.n36955 vdd.n36951 3.931
R48629 vdd.n36969 vdd.n36965 3.931
R48630 vdd.n33147 vdd.n33143 3.931
R48631 vdd.n35641 vdd.n35637 3.931
R48632 vdd.n37323 vdd.n37319 3.931
R48633 vdd.n37353 vdd.n37349 3.931
R48634 vdd.n35668 vdd.n35664 3.931
R48635 vdd.n32830 vdd.n32826 3.931
R48636 vdd.n38024 vdd.n38020 3.931
R48637 vdd.n38010 vdd.n38006 3.931
R48638 vdd.n37793 vdd.n37789 3.931
R48639 vdd.n37779 vdd.n37775 3.931
R48640 vdd.n28221 vdd.n28217 3.931
R48641 vdd.n28235 vdd.n28231 3.931
R48642 vdd.n28452 vdd.n28448 3.931
R48643 vdd.n28466 vdd.n28462 3.931
R48644 vdd.n28683 vdd.n28679 3.931
R48645 vdd.n28697 vdd.n28693 3.931
R48646 vdd.n26700 vdd.n26699 3.931
R48647 vdd.n26309 vdd.n26308 3.931
R48648 vdd.n27985 vdd.n27981 3.931
R48649 vdd.n27882 vdd.n27878 3.931
R48650 vdd.n31459 vdd.n31458 3.931
R48651 vdd.n32402 vdd.n32401 3.931
R48652 vdd.n2886 vdd.n2885 3.931
R48653 vdd.n2896 vdd.n2895 3.931
R48654 vdd.n3067 vdd.n3066 3.931
R48655 vdd.n3077 vdd.n3076 3.931
R48656 vdd.n3248 vdd.n3247 3.931
R48657 vdd.n3258 vdd.n3257 3.931
R48658 vdd.n3429 vdd.n3428 3.931
R48659 vdd.n3439 vdd.n3438 3.931
R48660 vdd.n3610 vdd.n3609 3.931
R48661 vdd.n3620 vdd.n3619 3.931
R48662 vdd.n3897 vdd.n3896 3.931
R48663 vdd.n3814 vdd.n3813 3.931
R48664 vdd.n2525 vdd.n2524 3.931
R48665 vdd.n2495 vdd.n2494 3.931
R48666 vdd.n1240 vdd.n1239 3.931
R48667 vdd.n1816 vdd.n1815 3.931
R48668 vdd.n1658 vdd.n1657 3.931
R48669 vdd.n1648 vdd.n1647 3.931
R48670 vdd.n1477 vdd.n1476 3.931
R48671 vdd.n1467 vdd.n1466 3.931
R48672 vdd.n1296 vdd.n1295 3.931
R48673 vdd.n26762 vdd.n26761 3.931
R48674 vdd.n26933 vdd.n26932 3.931
R48675 vdd.n26943 vdd.n26942 3.931
R48676 vdd.n27114 vdd.n27113 3.931
R48677 vdd.n27124 vdd.n27123 3.931
R48678 vdd.n26702 vdd.n26695 3.931
R48679 vdd.n26311 vdd.n26304 3.931
R48680 vdd.n31614 vdd.n31613 3.931
R48681 vdd.n31598 vdd.n31597 3.931
R48682 vdd.n31461 vdd.n31454 3.931
R48683 vdd.n32404 vdd.n32397 3.931
R48684 vdd.n13358 vdd.n9069 3.931
R48685 vdd.n13403 vdd.n9048 3.931
R48686 vdd.n13650 vdd.n8849 3.931
R48687 vdd.n13696 vdd.n8827 3.931
R48688 vdd.n13966 vdd.n8622 3.931
R48689 vdd.n13977 vdd.n8612 3.931
R48690 vdd.n14256 vdd.n8400 3.931
R48691 vdd.n14267 vdd.n8390 3.931
R48692 vdd.n14686 vdd.n14683 3.931
R48693 vdd.n14715 vdd.n8112 3.931
R48694 vdd.n14860 vdd.n14857 3.931
R48695 vdd.n14905 vdd.n8023 3.931
R48696 vdd.n13239 vdd.n9180 3.931
R48697 vdd.n13277 vdd.n9152 3.931
R48698 vdd.n13531 vdd.n8959 3.931
R48699 vdd.n13569 vdd.n8931 3.931
R48700 vdd.n13819 vdd.n8740 3.931
R48701 vdd.n13857 vdd.n8706 3.931
R48702 vdd.n14106 vdd.n8527 3.931
R48703 vdd.n14146 vdd.n8483 3.931
R48704 vdd.n14410 vdd.n8296 3.931
R48705 vdd.n8268 vdd.n8240 3.931
R48706 vdd.n19268 vdd.n19262 3.931
R48707 vdd.n19256 vdd.n19250 3.931
R48708 vdd.n19212 vdd.n19206 3.931
R48709 vdd.n19200 vdd.n19194 3.931
R48710 vdd.n19854 vdd.n19848 3.931
R48711 vdd.n19866 vdd.n19860 3.931
R48712 vdd.n19922 vdd.n19916 3.931
R48713 vdd.n19934 vdd.n19928 3.931
R48714 vdd.n21529 vdd.n21523 3.931
R48715 vdd.n21511 vdd.n21505 3.931
R48716 vdd.n21270 vdd.n21264 3.931
R48717 vdd.n21252 vdd.n21246 3.931
R48718 vdd.n19146 vdd.n19145 3.931
R48719 vdd.n19138 vdd.n19137 3.931
R48720 vdd.n18904 vdd.n18898 3.931
R48721 vdd.n18886 vdd.n18880 3.931
R48722 vdd.n18645 vdd.n18639 3.931
R48723 vdd.n18627 vdd.n18621 3.931
R48724 vdd.n20396 vdd.n20395 3.931
R48725 vdd.n20373 vdd.n20372 3.931
R48726 vdd.n20160 vdd.n20159 3.931
R48727 vdd.n20137 vdd.n20136 3.931
R48728 vdd.n24754 vdd.n24753 3.931
R48729 vdd.n25156 vdd.n25155 3.931
R48730 vdd.n10392 vdd.n10326 3.872
R48731 vdd.n10393 vdd.n9297 3.872
R48732 vdd.n10347 vdd.n10346 3.87
R48733 vdd.n10376 vdd.n10375 3.87
R48734 vdd.n9445 vdd.n9425 3.87
R48735 vdd.n9449 vdd.n9419 3.87
R48736 vdd.n12893 vdd.n12892 3.87
R48737 vdd.n9638 vdd.n9635 3.87
R48738 vdd.n9804 vdd.n9785 3.87
R48739 vdd.n9808 vdd.n9780 3.87
R48740 vdd.n12685 vdd.n12684 3.87
R48741 vdd.n9998 vdd.n9995 3.87
R48742 vdd.n15256 vdd.n15255 3.87
R48743 vdd.n15245 vdd.n15244 3.87
R48744 vdd.n15234 vdd.n15233 3.87
R48745 vdd.n15220 vdd.n15219 3.87
R48746 vdd.n15206 vdd.n15205 3.87
R48747 vdd.n15180 vdd.n15179 3.87
R48748 vdd.n15178 vdd.n15177 3.87
R48749 vdd.n15164 vdd.n15163 3.87
R48750 vdd.n15150 vdd.n15149 3.87
R48751 vdd.n15136 vdd.n15135 3.87
R48752 vdd.n10369 vdd.n10368 3.851
R48753 vdd.n13001 vdd.n9407 3.851
R48754 vdd.n9439 vdd.t360 3.851
R48755 vdd.n12986 vdd.n12985 3.851
R48756 vdd.n12974 vdd.n12973 3.851
R48757 vdd.t366 vdd.n9555 3.851
R48758 vdd.n9596 vdd.n9570 3.851
R48759 vdd.n12879 vdd.n9615 3.851
R48760 vdd.n9649 vdd.n9648 3.851
R48761 vdd.n12793 vdd.n9767 3.851
R48762 vdd.n12778 vdd.n12777 3.851
R48763 vdd.n12766 vdd.n12765 3.851
R48764 vdd.n9956 vdd.n9929 3.851
R48765 vdd.n12671 vdd.n9975 3.851
R48766 vdd.n10009 vdd.n10008 3.851
R48767 vdd.n12595 vdd.t83 3.851
R48768 vdd.n10486 vdd.n10485 3.851
R48769 vdd.t80 vdd.n10486 3.851
R48770 vdd.n10493 vdd.n10479 3.851
R48771 vdd.n12520 vdd.n12519 3.851
R48772 vdd.n12453 vdd.n10623 3.851
R48773 vdd.n12415 vdd.n12414 3.851
R48774 vdd.n12343 vdd.n10816 3.851
R48775 vdd.n10885 vdd.n10884 3.851
R48776 vdd.n12252 vdd.n12251 3.851
R48777 vdd.n11050 vdd.n11047 3.851
R48778 vdd.t298 vdd.n11169 3.851
R48779 vdd.n12115 vdd.n11191 3.851
R48780 vdd.n12037 vdd.n11325 3.851
R48781 vdd.n11394 vdd.n11393 3.851
R48782 vdd.t186 vdd.n11926 3.851
R48783 vdd.n15440 vdd.n15439 3.851
R48784 vdd.n15642 vdd.n15641 3.851
R48785 vdd.n15229 vdd.t28 3.851
R48786 vdd.n15678 vdd.n15677 3.851
R48787 vdd.n15696 vdd.n15695 3.851
R48788 vdd.t34 vdd.n15845 3.851
R48789 vdd.n15898 vdd.n15897 3.851
R48790 vdd.n15934 vdd.n15933 3.851
R48791 vdd.n15952 vdd.n15951 3.851
R48792 vdd.n16154 vdd.n16153 3.851
R48793 vdd.n16190 vdd.n16189 3.851
R48794 vdd.n16208 vdd.n16207 3.851
R48795 vdd.n16410 vdd.n16409 3.851
R48796 vdd.n16446 vdd.n16445 3.851
R48797 vdd.n16464 vdd.n16463 3.851
R48798 vdd.t337 vdd.n16633 3.851
R48799 vdd.n15074 vdd.n15073 3.851
R48800 vdd.t336 vdd.n15074 3.851
R48801 vdd.n15085 vdd.n15084 3.851
R48802 vdd.n16883 vdd.n16882 3.851
R48803 vdd.n17071 vdd.n17070 3.851
R48804 vdd.n17155 vdd.n17154 3.851
R48805 vdd.n17343 vdd.n17342 3.851
R48806 vdd.n17427 vdd.n17426 3.851
R48807 vdd.n17601 vdd.n17600 3.851
R48808 vdd.n17685 vdd.n17684 3.851
R48809 vdd.t258 vdd.n17872 3.851
R48810 vdd.n17956 vdd.n17955 3.851
R48811 vdd.n18144 vdd.n18143 3.851
R48812 vdd.n18227 vdd.n18226 3.851
R48813 vdd.n21706 vdd.t177 3.851
R48814 vdd.n24727 vdd.n24726 3.85
R48815 vdd.n25185 vdd.n25184 3.85
R48816 vdd.n25184 vdd.n25183 3.85
R48817 vdd.n24726 vdd.n24725 3.85
R48818 vdd.n11486 vdd.n11469 3.85
R48819 vdd.n11466 vdd.n11433 3.85
R48820 vdd.n16818 vdd.n16810 3.85
R48821 vdd.n15038 vdd.n15037 3.85
R48822 vdd.n33527 vdd.n33526 3.843
R48823 vdd.n1010 vdd.n1009 3.843
R48824 vdd.n15394 vdd.n15393 3.843
R48825 vdd.n15409 vdd.n15408 3.843
R48826 vdd.n13153 vdd.n13152 3.838
R48827 vdd.n13187 vdd.n13186 3.838
R48828 vdd.n5078 vdd.n5077 3.836
R48829 vdd.n34119 vdd.n34118 3.829
R48830 vdd.n35506 vdd.n35505 3.829
R48831 vdd.n34973 vdd.n34972 3.829
R48832 vdd.n5986 vdd.n5985 3.829
R48833 vdd.n5720 vdd.n5719 3.829
R48834 vdd.n4550 vdd.n4549 3.829
R48835 vdd.n27395 vdd.n27394 3.829
R48836 vdd.n25841 vdd.n25840 3.829
R48837 vdd.n268 vdd.n267 3.821
R48838 vdd.n33580 vdd.n33579 3.814
R48839 vdd.n923 vdd.n922 3.814
R48840 vdd.n22212 vdd.n22211 3.808
R48841 vdd.n22076 vdd.n22075 3.808
R48842 vdd.n32092 vdd.n32091 3.8
R48843 vdd.n32408 vdd.n32407 3.799
R48844 vdd.n10385 vdd.n10384 3.792
R48845 vdd.n10383 vdd.n10342 3.792
R48846 vdd.n9437 vdd.n9418 3.792
R48847 vdd.n12991 vdd.n12990 3.792
R48848 vdd.n12885 vdd.n9605 3.792
R48849 vdd.n12884 vdd.n12883 3.792
R48850 vdd.n9796 vdd.n9779 3.792
R48851 vdd.n12783 vdd.n12782 3.792
R48852 vdd.n12677 vdd.n9965 3.792
R48853 vdd.n12676 vdd.n12675 3.792
R48854 vdd.n10185 vdd.n10184 3.792
R48855 vdd.n10593 vdd.n10590 3.792
R48856 vdd.n12475 vdd.n10588 3.792
R48857 vdd.n12434 vdd.n10661 3.792
R48858 vdd.n10686 vdd.n10678 3.792
R48859 vdd.n12379 vdd.n12378 3.792
R48860 vdd.n10786 vdd.n10754 3.792
R48861 vdd.n10848 vdd.n10847 3.792
R48862 vdd.n10858 vdd.n10829 3.792
R48863 vdd.n10943 vdd.n10942 3.792
R48864 vdd.n10947 vdd.n10924 3.792
R48865 vdd.n11026 vdd.n11019 3.792
R48866 vdd.n12232 vdd.n11015 3.792
R48867 vdd.n12183 vdd.n12182 3.792
R48868 vdd.n11123 vdd.n11122 3.792
R48869 vdd.n12130 vdd.n11176 3.792
R48870 vdd.n12124 vdd.n11182 3.792
R48871 vdd.n12080 vdd.n11245 3.792
R48872 vdd.n11295 vdd.n11271 3.792
R48873 vdd.n11357 vdd.n11356 3.792
R48874 vdd.n11367 vdd.n11338 3.792
R48875 vdd.n15247 vdd.n15246 3.792
R48876 vdd.n15236 vdd.n15235 3.792
R48877 vdd.n15222 vdd.n15221 3.792
R48878 vdd.n15208 vdd.n15207 3.792
R48879 vdd.n15182 vdd.n15181 3.792
R48880 vdd.n15191 vdd.n15190 3.792
R48881 vdd.n15166 vdd.n15165 3.792
R48882 vdd.n15152 vdd.n15151 3.792
R48883 vdd.n15138 vdd.n15137 3.792
R48884 vdd.n15124 vdd.n15123 3.792
R48885 vdd.n16716 vdd.n16715 3.792
R48886 vdd.n16979 vdd.n16970 3.792
R48887 vdd.n16995 vdd.n16994 3.792
R48888 vdd.n17105 vdd.n17096 3.792
R48889 vdd.n17125 vdd.n17112 3.792
R48890 vdd.n17251 vdd.n17242 3.792
R48891 vdd.n17267 vdd.n17266 3.792
R48892 vdd.n17377 vdd.n17368 3.792
R48893 vdd.n17397 vdd.n17384 3.792
R48894 vdd.n17523 vdd.n17514 3.792
R48895 vdd.n17539 vdd.n17538 3.792
R48896 vdd.n17635 vdd.n17626 3.792
R48897 vdd.n17655 vdd.n17642 3.792
R48898 vdd.n17781 vdd.n17772 3.792
R48899 vdd.n17797 vdd.n17796 3.792
R48900 vdd.n17906 vdd.n17897 3.792
R48901 vdd.n17926 vdd.n17913 3.792
R48902 vdd.n18052 vdd.n18043 3.792
R48903 vdd.n18068 vdd.n18067 3.792
R48904 vdd.n18178 vdd.n18169 3.792
R48905 vdd.n18198 vdd.n18185 3.792
R48906 vdd.n33581 vdd.n33580 3.764
R48907 vdd.n34374 vdd.n34373 3.764
R48908 vdd.n35397 vdd.n35396 3.764
R48909 vdd.n34800 vdd.n34799 3.764
R48910 vdd.n924 vdd.n923 3.764
R48911 vdd.n6088 vdd.n6087 3.764
R48912 vdd.n5547 vdd.n5546 3.764
R48913 vdd.n4763 vdd.n4762 3.764
R48914 vdd.n4841 vdd.n4840 3.764
R48915 vdd.n4374 vdd.n4373 3.764
R48916 vdd.n31277 vdd.n31270 3.764
R48917 vdd.n30516 vdd.n30512 3.764
R48918 vdd.n35871 vdd.n35864 3.764
R48919 vdd.n35976 vdd.n35969 3.764
R48920 vdd.n36102 vdd.n36095 3.764
R48921 vdd.n36207 vdd.n36200 3.764
R48922 vdd.n36333 vdd.n36326 3.764
R48923 vdd.n36438 vdd.n36431 3.764
R48924 vdd.n36564 vdd.n36557 3.764
R48925 vdd.n36669 vdd.n36662 3.764
R48926 vdd.n36795 vdd.n36788 3.764
R48927 vdd.n36900 vdd.n36893 3.764
R48928 vdd.n37040 vdd.n37036 3.764
R48929 vdd.n37113 vdd.n37109 3.764
R48930 vdd.n33114 vdd.n33110 3.764
R48931 vdd.n33035 vdd.n33031 3.764
R48932 vdd.n37409 vdd.n37402 3.764
R48933 vdd.n32868 vdd.n32864 3.764
R48934 vdd.n38182 vdd.n38178 3.764
R48935 vdd.n38081 vdd.n38074 3.764
R48936 vdd.n37955 vdd.n37948 3.764
R48937 vdd.n37850 vdd.n37843 3.764
R48938 vdd.n37724 vdd.n37717 3.764
R48939 vdd.n37619 vdd.n37612 3.764
R48940 vdd.n28292 vdd.n28285 3.764
R48941 vdd.n28397 vdd.n28390 3.764
R48942 vdd.n28523 vdd.n28516 3.764
R48943 vdd.n28628 vdd.n28621 3.764
R48944 vdd.n28754 vdd.n28747 3.764
R48945 vdd.n30206 vdd.n30205 3.764
R48946 vdd.n27268 vdd.n27267 3.764
R48947 vdd.n25923 vdd.n25922 3.764
R48948 vdd.n1284 vdd.n1277 3.764
R48949 vdd.n1703 vdd.n1699 3.764
R48950 vdd.n1605 vdd.n1601 3.764
R48951 vdd.n1522 vdd.n1518 3.764
R48952 vdd.n1424 vdd.n1420 3.764
R48953 vdd.n1341 vdd.n1337 3.764
R48954 vdd.n26807 vdd.n26803 3.764
R48955 vdd.n26890 vdd.n26886 3.764
R48956 vdd.n26988 vdd.n26984 3.764
R48957 vdd.n27071 vdd.n27067 3.764
R48958 vdd.n27169 vdd.n27165 3.764
R48959 vdd.n2115 vdd.n2114 3.764
R48960 vdd.n2125 vdd.n2124 3.764
R48961 vdd.n2161 vdd.n2160 3.764
R48962 vdd.n2144 vdd.n2143 3.764
R48963 vdd.n3795 vdd.n3794 3.764
R48964 vdd.n2760 vdd.n2756 3.764
R48965 vdd.n2843 vdd.n2839 3.764
R48966 vdd.n2941 vdd.n2937 3.764
R48967 vdd.n3024 vdd.n3020 3.764
R48968 vdd.n3122 vdd.n3118 3.764
R48969 vdd.n3205 vdd.n3201 3.764
R48970 vdd.n3303 vdd.n3299 3.764
R48971 vdd.n3386 vdd.n3382 3.764
R48972 vdd.n3484 vdd.n3480 3.764
R48973 vdd.n3567 vdd.n3563 3.764
R48974 vdd.n13196 vdd.n13195 3.764
R48975 vdd.n13195 vdd.n9217 3.764
R48976 vdd.n13291 vdd.n9145 3.764
R48977 vdd.n13301 vdd.n9145 3.764
R48978 vdd.n13490 vdd.n13489 3.764
R48979 vdd.n13489 vdd.n8997 3.764
R48980 vdd.n13583 vdd.n8924 3.764
R48981 vdd.n13593 vdd.n8924 3.764
R48982 vdd.n13770 vdd.n13769 3.764
R48983 vdd.n13769 vdd.n8780 3.764
R48984 vdd.n13850 vdd.n8685 3.764
R48985 vdd.n13897 vdd.n8685 3.764
R48986 vdd.n14048 vdd.n8572 3.764
R48987 vdd.n14048 vdd.n14047 3.764
R48988 vdd.n14139 vdd.n8461 3.764
R48989 vdd.n14186 vdd.n8461 3.764
R48990 vdd.n14323 vdd.n8355 3.764
R48991 vdd.n14323 vdd.n14322 3.764
R48992 vdd.n14455 vdd.n14454 3.764
R48993 vdd.n14454 vdd.n8249 3.764
R48994 vdd.n14648 vdd.n8153 3.764
R48995 vdd.n8157 vdd.n8155 3.764
R48996 vdd.n14752 vdd.n8096 3.764
R48997 vdd.n14762 vdd.n8092 3.764
R48998 vdd.n14820 vdd.n14809 3.764
R48999 vdd.n14813 vdd.n14811 3.764
R49000 vdd.n14922 vdd.n8005 3.764
R49001 vdd.n14928 vdd.n8006 3.764
R49002 vdd.n13164 vdd.n9232 3.764
R49003 vdd.n13164 vdd.n9233 3.764
R49004 vdd.n9120 vdd.n9119 3.764
R49005 vdd.n9119 vdd.n9113 3.764
R49006 vdd.n9012 vdd.n9009 3.764
R49007 vdd.n13458 vdd.n9009 3.764
R49008 vdd.n8899 vdd.n8898 3.764
R49009 vdd.n8898 vdd.n8892 3.764
R49010 vdd.n13748 vdd.n8790 3.764
R49011 vdd.n13748 vdd.n8787 3.764
R49012 vdd.n8654 vdd.n8653 3.764
R49013 vdd.n8653 vdd.n8639 3.764
R49014 vdd.n14036 vdd.n8578 3.764
R49015 vdd.n14036 vdd.n8579 3.764
R49016 vdd.n8434 vdd.n8433 3.764
R49017 vdd.n8433 vdd.n8417 3.764
R49018 vdd.n8360 vdd.n8321 3.764
R49019 vdd.n14370 vdd.n8321 3.764
R49020 vdd.n14533 vdd.n8194 3.764
R49021 vdd.n14534 vdd.n14533 3.764
R49022 vdd.n24254 vdd.n24253 3.764
R49023 vdd.n24263 vdd.n24262 3.764
R49024 vdd.n24152 vdd.n24151 3.764
R49025 vdd.n24014 vdd.n24013 3.764
R49026 vdd.n23920 vdd.n23919 3.764
R49027 vdd.n23782 vdd.n23781 3.764
R49028 vdd.n23688 vdd.n23687 3.764
R49029 vdd.n23094 vdd.n23093 3.764
R49030 vdd.n23232 vdd.n23231 3.764
R49031 vdd.n23326 vdd.n23325 3.764
R49032 vdd.n23464 vdd.n23463 3.764
R49033 vdd.n23558 vdd.n23557 3.764
R49034 vdd.n22515 vdd.n22514 3.764
R49035 vdd.n22653 vdd.n22652 3.764
R49036 vdd.n22747 vdd.n22746 3.764
R49037 vdd.n22885 vdd.n22884 3.764
R49038 vdd.n22979 vdd.n22978 3.764
R49039 vdd.n22426 vdd.n22425 3.764
R49040 vdd.n22435 vdd.n22434 3.764
R49041 vdd.n22282 vdd.n22281 3.764
R49042 vdd.n22291 vdd.n22290 3.764
R49043 vdd.n19369 vdd.n19360 3.764
R49044 vdd.n19482 vdd.n19473 3.764
R49045 vdd.n19575 vdd.n19566 3.764
R49046 vdd.n19682 vdd.n19673 3.764
R49047 vdd.n19777 vdd.n19768 3.764
R49048 vdd.n20974 vdd.n20965 3.764
R49049 vdd.n20879 vdd.n20870 3.764
R49050 vdd.n20783 vdd.n20774 3.764
R49051 vdd.n20691 vdd.n20682 3.764
R49052 vdd.n20578 vdd.n20569 3.764
R49053 vdd.n21594 vdd.n21585 3.764
R49054 vdd.n21448 vdd.n21439 3.764
R49055 vdd.n21335 vdd.n21326 3.764
R49056 vdd.n21189 vdd.n21180 3.764
R49057 vdd.n21076 vdd.n21067 3.764
R49058 vdd.n19082 vdd.n19073 3.764
R49059 vdd.n18969 vdd.n18960 3.764
R49060 vdd.n18823 vdd.n18814 3.764
R49061 vdd.n18710 vdd.n18701 3.764
R49062 vdd.n18564 vdd.n18555 3.764
R49063 vdd.n20307 vdd.n20306 3.764
R49064 vdd.n20225 vdd.n20224 3.764
R49065 vdd.n20071 vdd.n20070 3.764
R49066 vdd.n24687 vdd.n24686 3.764
R49067 vdd.n24800 vdd.n24799 3.764
R49068 vdd.n25218 vdd.n25217 3.764
R49069 vdd.n25105 vdd.n25104 3.764
R49070 vdd.n31527 vdd.n31524 3.739
R49071 vdd.n2159 vdd.n2158 3.699
R49072 vdd.n13237 vdd.n9178 3.67
R49073 vdd.n13266 vdd.n9165 3.67
R49074 vdd.n13375 vdd.n9062 3.67
R49075 vdd.n13404 vdd.n9045 3.67
R49076 vdd.n13390 vdd.n13389 3.67
R49077 vdd.n13446 vdd.n13445 3.67
R49078 vdd.n13548 vdd.n8949 3.67
R49079 vdd.n13558 vdd.n8944 3.67
R49080 vdd.n13620 vdd.t328 3.67
R49081 vdd.n13667 vdd.n8842 3.67
R49082 vdd.n13697 vdd.n8824 3.67
R49083 vdd.n13682 vdd.n13681 3.67
R49084 vdd.n13737 vdd.n13736 3.67
R49085 vdd.n13761 vdd.n13760 3.67
R49086 vdd.n13821 vdd.n13820 3.67
R49087 vdd.n13961 vdd.n8629 3.67
R49088 vdd.n13974 vdd.n8614 3.67
R49089 vdd.n14004 vdd.n8594 3.67
R49090 vdd.n14021 vdd.n8574 3.67
R49091 vdd.n14096 vdd.n8536 3.67
R49092 vdd.n14153 vdd.n8490 3.67
R49093 vdd.n14251 vdd.n8407 3.67
R49094 vdd.n14264 vdd.n8392 3.67
R49095 vdd.n14295 vdd.n8372 3.67
R49096 vdd.n14310 vdd.n8357 3.67
R49097 vdd.n14345 vdd.n8327 3.67
R49098 vdd.n14406 vdd.n8297 3.67
R49099 vdd.n14430 vdd.n8273 3.67
R49100 vdd.n14559 vdd.n8188 3.67
R49101 vdd.n14602 vdd.n14567 3.67
R49102 vdd.n12522 vdd.n10519 3.638
R49103 vdd.n12444 vdd.n10655 3.638
R49104 vdd.n12424 vdd.n10674 3.638
R49105 vdd.n10818 vdd.n10815 3.638
R49106 vdd.n10875 vdd.n10857 3.638
R49107 vdd.n11001 vdd.n10995 3.638
R49108 vdd.n12221 vdd.n11036 3.638
R49109 vdd.n12143 vdd.n11147 3.638
R49110 vdd.n11212 vdd.n11199 3.638
R49111 vdd.n11327 vdd.n11324 3.638
R49112 vdd.n11384 vdd.n11366 3.638
R49113 vdd.n11934 vdd.n11550 3.638
R49114 vdd.n10395 vdd.n10391 3.638
R49115 vdd.n10371 vdd.n10355 3.638
R49116 vdd.n9432 vdd.n9408 3.638
R49117 vdd.n12983 vdd.n9422 3.638
R49118 vdd.n12897 vdd.n9573 3.638
R49119 vdd.n9645 vdd.n9631 3.638
R49120 vdd.n9792 vdd.n9768 3.638
R49121 vdd.n12775 vdd.n9782 3.638
R49122 vdd.n12689 vdd.n9932 3.638
R49123 vdd.n10005 vdd.n9991 3.638
R49124 vdd.n10489 vdd.n10488 3.638
R49125 vdd.n16837 vdd.n16836 3.638
R49126 vdd.n17082 vdd.n17081 3.638
R49127 vdd.n17134 vdd.n17133 3.638
R49128 vdd.n17354 vdd.n17353 3.638
R49129 vdd.n17406 vdd.n17405 3.638
R49130 vdd.n17612 vdd.n17611 3.638
R49131 vdd.n17664 vdd.n17663 3.638
R49132 vdd.n17883 vdd.n17882 3.638
R49133 vdd.n17935 vdd.n17934 3.638
R49134 vdd.n18155 vdd.n18154 3.638
R49135 vdd.n18207 vdd.n18206 3.638
R49136 vdd.n15013 vdd.n15012 3.638
R49137 vdd.n15411 vdd.n15406 3.638
R49138 vdd.n15428 vdd.n15424 3.638
R49139 vdd.n15661 vdd.n15654 3.638
R49140 vdd.n15681 vdd.n15674 3.638
R49141 vdd.n15917 vdd.n15910 3.638
R49142 vdd.n15937 vdd.n15930 3.638
R49143 vdd.n16173 vdd.n16166 3.638
R49144 vdd.n16193 vdd.n16186 3.638
R49145 vdd.n16429 vdd.n16422 3.638
R49146 vdd.n16449 vdd.n16442 3.638
R49147 vdd.n15078 vdd.n15077 3.638
R49148 vdd.n28133 vdd.n28132 3.635
R49149 vdd.n35911 vdd.n35910 3.576
R49150 vdd.n35932 vdd.n35931 3.576
R49151 vdd.n36142 vdd.n36141 3.576
R49152 vdd.n36163 vdd.n36162 3.576
R49153 vdd.n36373 vdd.n36372 3.576
R49154 vdd.n36394 vdd.n36393 3.576
R49155 vdd.n36604 vdd.n36603 3.576
R49156 vdd.n36625 vdd.n36624 3.576
R49157 vdd.n36835 vdd.n36834 3.576
R49158 vdd.n36856 vdd.n36855 3.576
R49159 vdd.n33266 vdd.n33265 3.576
R49160 vdd.n33248 vdd.n33247 3.576
R49161 vdd.n33072 vdd.n33071 3.576
R49162 vdd.n37258 vdd.n37257 3.576
R49163 vdd.n37444 vdd.n37442 3.576
R49164 vdd.n32912 vdd.n32911 3.576
R49165 vdd.n38123 vdd.n38122 3.576
R49166 vdd.n38134 vdd.n38133 3.576
R49167 vdd.n37911 vdd.n37909 3.576
R49168 vdd.n37890 vdd.n37889 3.576
R49169 vdd.n37680 vdd.n37678 3.576
R49170 vdd.n37659 vdd.n37658 3.576
R49171 vdd.n28332 vdd.n28331 3.576
R49172 vdd.n28353 vdd.n28352 3.576
R49173 vdd.n28563 vdd.n28562 3.576
R49174 vdd.n28584 vdd.n28583 3.576
R49175 vdd.n28794 vdd.n28793 3.576
R49176 vdd.n28151 vdd.n28150 3.576
R49177 vdd.n27766 vdd.n27764 3.576
R49178 vdd.n31891 vdd.n31887 3.576
R49179 vdd.n32229 vdd.n32225 3.576
R49180 vdd.n29692 vdd.n29691 3.576
R49181 vdd.n30298 vdd.n30296 3.576
R49182 vdd.n30566 vdd.n30565 3.576
R49183 vdd.n34094 vdd.n34093 3.573
R49184 vdd.n35255 vdd.n35254 3.573
R49185 vdd.n34671 vdd.n34670 3.573
R49186 vdd.n5799 vdd.n5798 3.573
R49187 vdd.n5418 vdd.n5417 3.573
R49188 vdd.n4248 vdd.n4247 3.573
R49189 vdd.n27369 vdd.n27368 3.573
R49190 vdd.n25737 vdd.n25736 3.573
R49191 vdd.n28143 vdd.n28142 3.573
R49192 vdd.n250 vdd.n249 3.572
R49193 vdd.n25578 vdd.n25575 3.572
R49194 vdd.n10451 vdd.n10288 3.555
R49195 vdd.n10451 vdd.n10450 3.555
R49196 vdd.n10301 vdd.n10299 3.555
R49197 vdd.n10439 vdd.n10299 3.555
R49198 vdd.n9345 vdd.n9335 3.555
R49199 vdd.n9346 vdd.n9345 3.555
R49200 vdd.n13035 vdd.n9333 3.555
R49201 vdd.n13035 vdd.n13034 3.555
R49202 vdd.n12944 vdd.n12943 3.555
R49203 vdd.n12943 vdd.n9511 3.555
R49204 vdd.n9536 vdd.n9535 3.555
R49205 vdd.n9543 vdd.n9536 3.555
R49206 vdd.n9705 vdd.n9695 3.555
R49207 vdd.n9706 vdd.n9705 3.555
R49208 vdd.n12827 vdd.n9693 3.555
R49209 vdd.n12827 vdd.n12826 3.555
R49210 vdd.n12736 vdd.n12735 3.555
R49211 vdd.n12735 vdd.n9871 3.555
R49212 vdd.n9897 vdd.n9896 3.555
R49213 vdd.n9903 vdd.n9897 3.555
R49214 vdd.n10159 vdd.n10152 3.555
R49215 vdd.n10594 vdd.n10569 3.555
R49216 vdd.n12480 vdd.n10587 3.555
R49217 vdd.n12434 vdd.n10662 3.555
R49218 vdd.n10694 vdd.n10675 3.555
R49219 vdd.n12380 vdd.n10747 3.555
R49220 vdd.n10760 vdd.n10753 3.555
R49221 vdd.n10849 vdd.n10848 3.555
R49222 vdd.n12327 vdd.n12326 3.555
R49223 vdd.n10941 vdd.n10927 3.555
R49224 vdd.n12282 vdd.n12281 3.555
R49225 vdd.n11026 vdd.n11020 3.555
R49226 vdd.n12226 vdd.n11016 3.555
R49227 vdd.n11097 vdd.n11090 3.555
R49228 vdd.n11115 vdd.n11112 3.555
R49229 vdd.n12130 vdd.n12129 3.555
R49230 vdd.n11207 vdd.n11201 3.555
R49231 vdd.n12082 vdd.n12081 3.555
R49232 vdd.n12070 vdd.n12069 3.555
R49233 vdd.n11358 vdd.n11357 3.555
R49234 vdd.n12021 vdd.n12020 3.555
R49235 vdd.n11485 vdd.n11471 3.555
R49236 vdd.n11976 vdd.n11975 3.555
R49237 vdd.n15305 vdd.n15296 3.555
R49238 vdd.n15307 vdd.n15305 3.555
R49239 vdd.n15327 vdd.n15326 3.555
R49240 vdd.n15326 vdd.n15317 3.555
R49241 vdd.n15533 vdd.n15521 3.555
R49242 vdd.n15535 vdd.n15533 3.555
R49243 vdd.n15561 vdd.n15560 3.555
R49244 vdd.n15560 vdd.n15545 3.555
R49245 vdd.n15789 vdd.n15777 3.555
R49246 vdd.n15791 vdd.n15789 3.555
R49247 vdd.n15817 vdd.n15816 3.555
R49248 vdd.n15816 vdd.n15801 3.555
R49249 vdd.n16045 vdd.n16033 3.555
R49250 vdd.n16047 vdd.n16045 3.555
R49251 vdd.n16073 vdd.n16072 3.555
R49252 vdd.n16072 vdd.n16057 3.555
R49253 vdd.n16301 vdd.n16289 3.555
R49254 vdd.n16303 vdd.n16301 3.555
R49255 vdd.n16329 vdd.n16328 3.555
R49256 vdd.n16328 vdd.n16313 3.555
R49257 vdd.n16573 vdd.n16544 3.555
R49258 vdd.n16956 vdd.n16955 3.555
R49259 vdd.n16984 vdd.n16983 3.555
R49260 vdd.n17107 vdd.n17105 3.555
R49261 vdd.n17142 vdd.n17141 3.555
R49262 vdd.n17228 vdd.n17227 3.555
R49263 vdd.n17256 vdd.n17255 3.555
R49264 vdd.n17379 vdd.n17377 3.555
R49265 vdd.n17414 vdd.n17413 3.555
R49266 vdd.n17500 vdd.n17499 3.555
R49267 vdd.n17528 vdd.n17527 3.555
R49268 vdd.n17637 vdd.n17635 3.555
R49269 vdd.n17672 vdd.n17671 3.555
R49270 vdd.n17758 vdd.n17757 3.555
R49271 vdd.n17786 vdd.n17785 3.555
R49272 vdd.n17908 vdd.n17906 3.555
R49273 vdd.n17943 vdd.n17942 3.555
R49274 vdd.n18029 vdd.n18028 3.555
R49275 vdd.n18057 vdd.n18056 3.555
R49276 vdd.n18180 vdd.n18178 3.555
R49277 vdd.n18215 vdd.n18214 3.555
R49278 vdd.n18296 vdd.n18295 3.555
R49279 vdd.n15028 vdd.n15027 3.555
R49280 vdd.n10467 vdd.n10277 3.549
R49281 vdd.n10318 vdd.n10307 3.549
R49282 vdd.n15273 vdd.n15272 3.549
R49283 vdd.t138 vdd.t100 3.538
R49284 vdd.n24846 vdd.n24843 3.538
R49285 vdd.n13074 vdd.t296 3.53
R49286 vdd.n13060 vdd.n13059 3.53
R49287 vdd.n9354 vdd.n9329 3.53
R49288 vdd.n9386 vdd.n9385 3.53
R49289 vdd.n9499 vdd.n9474 3.53
R49290 vdd.n9539 vdd.n9538 3.53
R49291 vdd.n12919 vdd.n12918 3.53
R49292 vdd.n9714 vdd.n9689 3.53
R49293 vdd.n9746 vdd.n9745 3.53
R49294 vdd.n9859 vdd.n9834 3.53
R49295 vdd.n9900 vdd.n9899 3.53
R49296 vdd.n12711 vdd.n12710 3.53
R49297 vdd.n12644 vdd.n12643 3.53
R49298 vdd.n10056 vdd.n10047 3.53
R49299 vdd.n10191 vdd.n10190 3.53
R49300 vdd.n10614 vdd.n10605 3.53
R49301 vdd.n10739 vdd.n10738 3.53
R49302 vdd.n10797 vdd.n10796 3.53
R49303 vdd.n10909 vdd.n10905 3.53
R49304 vdd.n12270 vdd.n12269 3.53
R49305 vdd.n12203 vdd.n11057 3.53
R49306 vdd.n12163 vdd.n12162 3.53
R49307 vdd.n12090 vdd.n11231 3.53
R49308 vdd.n11306 vdd.n11305 3.53
R49309 vdd.n11418 vdd.n11415 3.53
R49310 vdd.n11964 vdd.n11963 3.53
R49311 vdd.n15461 vdd.t249 3.53
R49312 vdd.n15495 vdd.n15491 3.53
R49313 vdd.n15558 vdd.n15555 3.53
R49314 vdd.n15592 vdd.n15591 3.53
R49315 vdd.n15751 vdd.n15747 3.53
R49316 vdd.n15814 vdd.n15811 3.53
R49317 vdd.n15848 vdd.n15847 3.53
R49318 vdd.n16070 vdd.n16067 3.53
R49319 vdd.n16104 vdd.n16103 3.53
R49320 vdd.n16263 vdd.n16259 3.53
R49321 vdd.n16326 vdd.n16323 3.53
R49322 vdd.n16360 vdd.n16359 3.53
R49323 vdd.n16519 vdd.n16515 3.53
R49324 vdd.n16560 vdd.n16558 3.53
R49325 vdd.n16611 vdd.n16610 3.53
R49326 vdd.n17022 vdd.n17019 3.53
R49327 vdd.n17202 vdd.n17199 3.53
R49328 vdd.n17294 vdd.n17291 3.53
R49329 vdd.n17474 vdd.n17471 3.53
R49330 vdd.n17566 vdd.n17563 3.53
R49331 vdd.n17732 vdd.n17729 3.53
R49332 vdd.n17824 vdd.n17821 3.53
R49333 vdd.n18003 vdd.n18000 3.53
R49334 vdd.n18095 vdd.n18092 3.53
R49335 vdd.n18271 vdd.n18269 3.53
R49336 vdd.n18343 vdd.n18341 3.53
R49337 vdd.n24200 vdd.n24196 3.529
R49338 vdd.n23978 vdd.n23974 3.529
R49339 vdd.n23968 vdd.n23964 3.529
R49340 vdd.n23746 vdd.n23742 3.529
R49341 vdd.n23736 vdd.n23732 3.529
R49342 vdd.n23058 vdd.n23054 3.529
R49343 vdd.n23280 vdd.n23276 3.529
R49344 vdd.n23290 vdd.n23286 3.529
R49345 vdd.n23512 vdd.n23508 3.529
R49346 vdd.n23522 vdd.n23518 3.529
R49347 vdd.n22479 vdd.n22475 3.529
R49348 vdd.n22701 vdd.n22697 3.529
R49349 vdd.n22711 vdd.n22707 3.529
R49350 vdd.n22933 vdd.n22929 3.529
R49351 vdd.n22943 vdd.n22939 3.529
R49352 vdd.n22183 vdd.n22179 3.529
R49353 vdd.n22266 vdd.n22261 3.529
R49354 vdd.n22277 vdd.n22273 3.529
R49355 vdd.n22151 vdd.n22146 3.529
R49356 vdd.n22162 vdd.n22158 3.529
R49357 vdd.n15353 vdd.n15352 3.523
R49358 vdd.n13118 vdd.n9245 3.518
R49359 vdd.n13229 vdd.n9191 3.518
R49360 vdd.n21615 vdd.n21611 3.518
R49361 vdd.n21429 vdd.n21426 3.518
R49362 vdd.n21348 vdd.n21345 3.518
R49363 vdd.n21250 vdd.t276 3.518
R49364 vdd.n21170 vdd.n21167 3.518
R49365 vdd.n21085 vdd.n21082 3.518
R49366 vdd.n19063 vdd.n19060 3.518
R49367 vdd.n18982 vdd.n18979 3.518
R49368 vdd.n18902 vdd.t344 3.518
R49369 vdd.n18804 vdd.n18801 3.518
R49370 vdd.n18723 vdd.n18720 3.518
R49371 vdd.n18545 vdd.n18542 3.518
R49372 vdd.n19335 vdd.n19334 3.518
R49373 vdd.n19511 vdd.n19510 3.518
R49374 vdd.n19541 vdd.n19540 3.518
R49375 vdd.n19712 vdd.n19711 3.518
R49376 vdd.n19743 vdd.n19742 3.518
R49377 vdd.n20940 vdd.n20939 3.518
R49378 vdd.n20909 vdd.n20908 3.518
R49379 vdd.n20750 vdd.n20749 3.518
R49380 vdd.n20720 vdd.n20719 3.518
R49381 vdd.n20544 vdd.n20543 3.518
R49382 vdd.n20451 vdd.t262 3.518
R49383 vdd.n20435 vdd.n20432 3.518
R49384 vdd.n20345 vdd.n20344 3.518
R49385 vdd.n20199 vdd.n20196 3.518
R49386 vdd.n20109 vdd.n20108 3.518
R49387 vdd.n20094 vdd.t256 3.518
R49388 vdd.n14673 vdd.n14672 3.509
R49389 vdd.n14730 vdd.n14729 3.509
R49390 vdd.n14845 vdd.n14844 3.509
R49391 vdd.n14914 vdd.n14913 3.509
R49392 vdd.t300 vdd.n8009 3.509
R49393 vdd.n51 vdd.n50 3.475
R49394 vdd.n28016 vdd.n28015 3.469
R49395 vdd.n33489 vdd.n33487 3.416
R49396 vdd.n34096 vdd.n34094 3.416
R49397 vdd.n35257 vdd.n35255 3.416
R49398 vdd.n34673 vdd.n34671 3.416
R49399 vdd.n976 vdd.n974 3.416
R49400 vdd.n5801 vdd.n5799 3.416
R49401 vdd.n5420 vdd.n5418 3.416
R49402 vdd.n4250 vdd.n4248 3.416
R49403 vdd.n27371 vdd.n27369 3.416
R49404 vdd.n25739 vdd.n25737 3.416
R49405 vdd.n3894 vdd.n3893 3.413
R49406 vdd.n10237 vdd.n10230 3.401
R49407 vdd.n16645 vdd.n16607 3.401
R49408 vdd.n1179 vdd.n1178 3.388
R49409 vdd.n30228 vdd.n30227 3.388
R49410 vdd.n32273 vdd.n32272 3.388
R49411 vdd.n32126 vdd.n32125 3.388
R49412 vdd.n32490 vdd.n32488 3.388
R49413 vdd.n31152 vdd.n31151 3.388
R49414 vdd.n30334 vdd.n30333 3.388
R49415 vdd.n35850 vdd.n35849 3.388
R49416 vdd.n35983 vdd.n35982 3.388
R49417 vdd.n36081 vdd.n36080 3.388
R49418 vdd.n36214 vdd.n36213 3.388
R49419 vdd.n36312 vdd.n36311 3.388
R49420 vdd.n36445 vdd.n36444 3.388
R49421 vdd.n36543 vdd.n36542 3.388
R49422 vdd.n36676 vdd.n36675 3.388
R49423 vdd.n36774 vdd.n36773 3.388
R49424 vdd.n36907 vdd.n36906 3.388
R49425 vdd.n37017 vdd.n37016 3.388
R49426 vdd.n33190 vdd.n33189 3.388
R49427 vdd.n37199 vdd.n37198 3.388
R49428 vdd.n33009 vdd.n33008 3.388
R49429 vdd.n32954 vdd.n32953 3.388
R49430 vdd.n37505 vdd.n37504 3.388
R49431 vdd.n38192 vdd.n38191 3.388
R49432 vdd.n38060 vdd.n38059 3.388
R49433 vdd.n37962 vdd.n37961 3.388
R49434 vdd.n37829 vdd.n37828 3.388
R49435 vdd.n37731 vdd.n37730 3.388
R49436 vdd.n37598 vdd.n37597 3.388
R49437 vdd.n28271 vdd.n28270 3.388
R49438 vdd.n28404 vdd.n28403 3.388
R49439 vdd.n28502 vdd.n28501 3.388
R49440 vdd.n28635 vdd.n28634 3.388
R49441 vdd.n28733 vdd.n28732 3.388
R49442 vdd.n28815 vdd.n28814 3.388
R49443 vdd.n28057 vdd.n28056 3.388
R49444 vdd.n29890 vdd.n29889 3.388
R49445 vdd.n29819 vdd.n29812 3.388
R49446 vdd.n29758 vdd.n29757 3.388
R49447 vdd.n25540 vdd.n25539 3.388
R49448 vdd.n25577 vdd.n25576 3.388
R49449 vdd.n1266 vdd.n1265 3.388
R49450 vdd.n1688 vdd.n1687 3.388
R49451 vdd.n1612 vdd.n1611 3.388
R49452 vdd.n1507 vdd.n1506 3.388
R49453 vdd.n1431 vdd.n1430 3.388
R49454 vdd.n1326 vdd.n1325 3.388
R49455 vdd.n26792 vdd.n26791 3.388
R49456 vdd.n26897 vdd.n26896 3.388
R49457 vdd.n26973 vdd.n26972 3.388
R49458 vdd.n27078 vdd.n27077 3.388
R49459 vdd.n27154 vdd.n27153 3.388
R49460 vdd.n1900 vdd.n1899 3.388
R49461 vdd.n2382 vdd.n2381 3.388
R49462 vdd.n2745 vdd.n2744 3.388
R49463 vdd.n2850 vdd.n2849 3.388
R49464 vdd.n2926 vdd.n2925 3.388
R49465 vdd.n3031 vdd.n3030 3.388
R49466 vdd.n3107 vdd.n3106 3.388
R49467 vdd.n3212 vdd.n3211 3.388
R49468 vdd.n3288 vdd.n3287 3.388
R49469 vdd.n3393 vdd.n3392 3.388
R49470 vdd.n3469 vdd.n3468 3.388
R49471 vdd.n3574 vdd.n3573 3.388
R49472 vdd.n3628 vdd.n3627 3.388
R49473 vdd.n13130 vdd.n13129 3.388
R49474 vdd.n9269 vdd.n9268 3.388
R49475 vdd.n13299 vdd.n9146 3.388
R49476 vdd.n13338 vdd.n9101 3.388
R49477 vdd.n13424 vdd.n13423 3.388
R49478 vdd.n9038 vdd.n9037 3.388
R49479 vdd.n13591 vdd.n8925 3.388
R49480 vdd.n13630 vdd.n8880 3.388
R49481 vdd.n13716 vdd.n13715 3.388
R49482 vdd.n8817 vdd.n8816 3.388
R49483 vdd.n13895 vdd.n8686 3.388
R49484 vdd.n8691 vdd.n8690 3.388
R49485 vdd.n14060 vdd.n8568 3.388
R49486 vdd.n14055 vdd.n8569 3.388
R49487 vdd.n14184 vdd.n8462 3.388
R49488 vdd.n8468 vdd.n8467 3.388
R49489 vdd.n14335 vdd.n8350 3.388
R49490 vdd.n14330 vdd.n8351 3.388
R49491 vdd.n8258 vdd.n8255 3.388
R49492 vdd.n14490 vdd.n8220 3.388
R49493 vdd.n14665 vdd.n14664 3.388
R49494 vdd.n14665 vdd.n8136 3.388
R49495 vdd.n14725 vdd.n8098 3.388
R49496 vdd.n14750 vdd.n8098 3.388
R49497 vdd.n14837 vdd.n14836 3.388
R49498 vdd.n14837 vdd.n8046 3.388
R49499 vdd.n14918 vdd.n8012 3.388
R49500 vdd.n14924 vdd.n8012 3.388
R49501 vdd.n13168 vdd.n13167 3.388
R49502 vdd.n13175 vdd.n9227 3.388
R49503 vdd.n13333 vdd.n13332 3.388
R49504 vdd.n9112 vdd.n9109 3.388
R49505 vdd.n13460 vdd.n9006 3.388
R49506 vdd.n13465 vdd.n9007 3.388
R49507 vdd.n13625 vdd.n13624 3.388
R49508 vdd.n8891 vdd.n8888 3.388
R49509 vdd.n13752 vdd.n8788 3.388
R49510 vdd.n13801 vdd.n13800 3.388
R49511 vdd.n13925 vdd.n8649 3.388
R49512 vdd.n13920 vdd.n8650 3.388
R49513 vdd.n14033 vdd.n14032 3.388
R49514 vdd.n14088 vdd.n14087 3.388
R49515 vdd.n14215 vdd.n8429 3.388
R49516 vdd.n14210 vdd.n8430 3.388
R49517 vdd.n14368 vdd.n8322 3.388
R49518 vdd.n8331 vdd.n8325 3.388
R49519 vdd.n14485 vdd.n14484 3.388
R49520 vdd.n14478 vdd.n8228 3.388
R49521 vdd.n24246 vdd.n24239 3.388
R49522 vdd.n24248 vdd.n24246 3.388
R49523 vdd.n24145 vdd.n24138 3.388
R49524 vdd.n24035 vdd.n24028 3.388
R49525 vdd.n23913 vdd.n23906 3.388
R49526 vdd.n23803 vdd.n23796 3.388
R49527 vdd.n23681 vdd.n23674 3.388
R49528 vdd.n23115 vdd.n23108 3.388
R49529 vdd.n23225 vdd.n23218 3.388
R49530 vdd.n23347 vdd.n23340 3.388
R49531 vdd.n23457 vdd.n23450 3.388
R49532 vdd.n23579 vdd.n23572 3.388
R49533 vdd.n22536 vdd.n22529 3.388
R49534 vdd.n22646 vdd.n22639 3.388
R49535 vdd.n22768 vdd.n22761 3.388
R49536 vdd.n22878 vdd.n22871 3.388
R49537 vdd.n23000 vdd.n22993 3.388
R49538 vdd.n22418 vdd.n22411 3.388
R49539 vdd.n22420 vdd.n22418 3.388
R49540 vdd.n22228 vdd.n22227 3.388
R49541 vdd.n22227 vdd.n22219 3.388
R49542 vdd.n24363 vdd.n24356 3.388
R49543 vdd.n24365 vdd.n24363 3.388
R49544 vdd.n22104 vdd.n22103 3.388
R49545 vdd.n22103 vdd.n22095 3.388
R49546 vdd.n19344 vdd.n19343 3.388
R49547 vdd.n19489 vdd.n19488 3.388
R49548 vdd.n19550 vdd.n19549 3.388
R49549 vdd.n19689 vdd.n19688 3.388
R49550 vdd.n19752 vdd.n19751 3.388
R49551 vdd.n20949 vdd.n20948 3.388
R49552 vdd.n20886 vdd.n20885 3.388
R49553 vdd.n20759 vdd.n20758 3.388
R49554 vdd.n20698 vdd.n20697 3.388
R49555 vdd.n20553 vdd.n20552 3.388
R49556 vdd.n21569 vdd.n21568 3.388
R49557 vdd.n21455 vdd.n21454 3.388
R49558 vdd.n21310 vdd.n21309 3.388
R49559 vdd.n21196 vdd.n21195 3.388
R49560 vdd.n21051 vdd.n21050 3.388
R49561 vdd.n19089 vdd.n19088 3.388
R49562 vdd.n18944 vdd.n18943 3.388
R49563 vdd.n18830 vdd.n18829 3.388
R49564 vdd.n18685 vdd.n18684 3.388
R49565 vdd.n18571 vdd.n18570 3.388
R49566 vdd.n20453 vdd.n20445 3.388
R49567 vdd.n20332 vdd.n20323 3.388
R49568 vdd.n20218 vdd.n20209 3.388
R49569 vdd.n20096 vdd.n20087 3.388
R49570 vdd.n24704 vdd.n24699 3.388
R49571 vdd.n24793 vdd.n24788 3.388
R49572 vdd.n25211 vdd.n25206 3.388
R49573 vdd.n25122 vdd.n25117 3.388
R49574 vdd.n13316 vdd.n9130 3.364
R49575 vdd.n13348 vdd.n9094 3.364
R49576 vdd.n13410 vdd.n9021 3.364
R49577 vdd.n13640 vdd.n8874 3.364
R49578 vdd.n13704 vdd.n8801 3.364
R49579 vdd.n13792 vdd.n13791 3.364
R49580 vdd.n13879 vdd.n8693 3.364
R49581 vdd.n13905 vdd.n8656 3.364
R49582 vdd.n13992 vdd.n8600 3.364
R49583 vdd.t124 vdd.n8565 3.364
R49584 vdd.n14079 vdd.n8512 3.364
R49585 vdd.n8535 vdd.t122 3.364
R49586 vdd.n14195 vdd.n14194 3.364
R49587 vdd.n14283 vdd.n8378 3.364
R49588 vdd.n14381 vdd.n8303 3.364
R49589 vdd.n14468 vdd.n8232 3.364
R49590 vdd.n14500 vdd.n8216 3.364
R49591 vdd.n36029 vdd.n36028 3.352
R49592 vdd.n36043 vdd.n36042 3.352
R49593 vdd.n36260 vdd.n36259 3.352
R49594 vdd.n36274 vdd.n36273 3.352
R49595 vdd.n36491 vdd.n36490 3.352
R49596 vdd.n36505 vdd.n36504 3.352
R49597 vdd.n36722 vdd.n36721 3.352
R49598 vdd.n36736 vdd.n36735 3.352
R49599 vdd.n36953 vdd.n36952 3.352
R49600 vdd.n36967 vdd.n36966 3.352
R49601 vdd.n33145 vdd.n33144 3.352
R49602 vdd.n35639 vdd.n35638 3.352
R49603 vdd.n37321 vdd.n37320 3.352
R49604 vdd.n37351 vdd.n37350 3.352
R49605 vdd.n35666 vdd.n35665 3.352
R49606 vdd.n32828 vdd.n32827 3.352
R49607 vdd.n38022 vdd.n38021 3.352
R49608 vdd.n38008 vdd.n38007 3.352
R49609 vdd.n37791 vdd.n37790 3.352
R49610 vdd.n37777 vdd.n37776 3.352
R49611 vdd.n28219 vdd.n28218 3.352
R49612 vdd.n28233 vdd.n28232 3.352
R49613 vdd.n28450 vdd.n28449 3.352
R49614 vdd.n28464 vdd.n28463 3.352
R49615 vdd.n28681 vdd.n28680 3.352
R49616 vdd.n28695 vdd.n28694 3.352
R49617 vdd.n26697 vdd.n26696 3.352
R49618 vdd.n26306 vdd.n26305 3.352
R49619 vdd.n27983 vdd.n27982 3.352
R49620 vdd.n27880 vdd.n27879 3.352
R49621 vdd.n31456 vdd.n31455 3.352
R49622 vdd.n32399 vdd.n32398 3.352
R49623 vdd.n10398 vdd.n10397 3.318
R49624 vdd.n10338 vdd.n10334 3.318
R49625 vdd.n10353 vdd.n10351 3.318
R49626 vdd.n10360 vdd.n10354 3.318
R49627 vdd.n9429 vdd.n9427 3.318
R49628 vdd.n9444 vdd.n9431 3.318
R49629 vdd.n12982 vdd.n9423 3.318
R49630 vdd.n12977 vdd.n9424 3.318
R49631 vdd.n9600 vdd.n9574 3.318
R49632 vdd.n9604 vdd.n9575 3.318
R49633 vdd.n9637 vdd.n9632 3.318
R49634 vdd.n9640 vdd.n9633 3.318
R49635 vdd.n9789 vdd.n9787 3.318
R49636 vdd.n9803 vdd.n9791 3.318
R49637 vdd.n12774 vdd.n9783 3.318
R49638 vdd.n12769 vdd.n9784 3.318
R49639 vdd.n9960 vdd.n9933 3.318
R49640 vdd.n9964 vdd.n9934 3.318
R49641 vdd.n9997 vdd.n9992 3.318
R49642 vdd.n10000 vdd.n9993 3.318
R49643 vdd.n12525 vdd.n12524 3.318
R49644 vdd.n12493 vdd.n12492 3.318
R49645 vdd.n12467 vdd.n10607 3.318
R49646 vdd.n12439 vdd.n10654 3.318
R49647 vdd.n12423 vdd.n10675 3.318
R49648 vdd.n12390 vdd.n10724 3.318
R49649 vdd.n10793 vdd.n10784 3.318
R49650 vdd.n10841 vdd.n10832 3.318
R49651 vdd.n12326 vdd.n10854 3.318
R49652 vdd.n10931 vdd.n10929 3.318
R49653 vdd.n10973 vdd.n10925 3.318
R49654 vdd.n12244 vdd.n10999 3.318
R49655 vdd.n12226 vdd.n11035 3.318
R49656 vdd.n12188 vdd.n12187 3.318
R49657 vdd.n12166 vdd.n11110 3.318
R49658 vdd.n12142 vdd.n12141 3.318
R49659 vdd.n11207 vdd.n11198 3.318
R49660 vdd.n11264 vdd.n11263 3.318
R49661 vdd.n11302 vdd.n11292 3.318
R49662 vdd.n11350 vdd.n11341 3.318
R49663 vdd.n12020 vdd.n11363 3.318
R49664 vdd.n11475 vdd.n11473 3.318
R49665 vdd.n11506 vdd.n11434 3.318
R49666 vdd.n11935 vdd.n11558 3.318
R49667 vdd.n15413 vdd.n15402 3.318
R49668 vdd.n15404 vdd.n15403 3.318
R49669 vdd.n15422 vdd.n15421 3.318
R49670 vdd.n15431 vdd.n15430 3.318
R49671 vdd.n15663 vdd.n15650 3.318
R49672 vdd.n15652 vdd.n15651 3.318
R49673 vdd.n15672 vdd.n15671 3.318
R49674 vdd.n15684 vdd.n15683 3.318
R49675 vdd.n15919 vdd.n15906 3.318
R49676 vdd.n15908 vdd.n15907 3.318
R49677 vdd.n15928 vdd.n15927 3.318
R49678 vdd.n15940 vdd.n15939 3.318
R49679 vdd.n16175 vdd.n16162 3.318
R49680 vdd.n16164 vdd.n16163 3.318
R49681 vdd.n16184 vdd.n16183 3.318
R49682 vdd.n16196 vdd.n16195 3.318
R49683 vdd.n16431 vdd.n16418 3.318
R49684 vdd.n16420 vdd.n16419 3.318
R49685 vdd.n16440 vdd.n16439 3.318
R49686 vdd.n16452 vdd.n16451 3.318
R49687 vdd.n16871 vdd.n16834 3.318
R49688 vdd.n16966 vdd.n16954 3.318
R49689 vdd.n17011 vdd.n17010 3.318
R49690 vdd.n17089 vdd.n17080 3.318
R49691 vdd.n17141 vdd.n17132 3.318
R49692 vdd.n17238 vdd.n17226 3.318
R49693 vdd.n17283 vdd.n17282 3.318
R49694 vdd.n17361 vdd.n17352 3.318
R49695 vdd.n17413 vdd.n17404 3.318
R49696 vdd.n17510 vdd.n17498 3.318
R49697 vdd.n17555 vdd.n17554 3.318
R49698 vdd.n17619 vdd.n17610 3.318
R49699 vdd.n17671 vdd.n17662 3.318
R49700 vdd.n17768 vdd.n17756 3.318
R49701 vdd.n17813 vdd.n17812 3.318
R49702 vdd.n17890 vdd.n17881 3.318
R49703 vdd.n17942 vdd.n17933 3.318
R49704 vdd.n18039 vdd.n18027 3.318
R49705 vdd.n18084 vdd.n18083 3.318
R49706 vdd.n18162 vdd.n18153 3.318
R49707 vdd.n18214 vdd.n18205 3.318
R49708 vdd.n18305 vdd.n18294 3.318
R49709 vdd.n18411 vdd.n18410 3.318
R49710 vdd.n25174 vdd.n25173 3.246
R49711 vdd.n24742 vdd.n24741 3.246
R49712 vdd.n10405 vdd.n10404 3.226
R49713 vdd.n13080 vdd.n9290 3.209
R49714 vdd.n13013 vdd.n13012 3.209
R49715 vdd.n12994 vdd.n12993 3.209
R49716 vdd.n9465 vdd.n9464 3.209
R49717 vdd.n9593 vdd.n9579 3.209
R49718 vdd.n12872 vdd.n9622 3.209
R49719 vdd.n12805 vdd.n12804 3.209
R49720 vdd.n9825 vdd.n9824 3.209
R49721 vdd.n9953 vdd.n9939 3.209
R49722 vdd.n9974 vdd.n9970 3.209
R49723 vdd.n12664 vdd.n9982 3.209
R49724 vdd.n10111 vdd.n10104 3.209
R49725 vdd.n12588 vdd.n12587 3.209
R49726 vdd.n10553 vdd.n10552 3.209
R49727 vdd.n10647 vdd.n10646 3.209
R49728 vdd.n10713 vdd.n10710 3.209
R49729 vdd.n12353 vdd.n12352 3.209
R49730 vdd.n12317 vdd.n10866 3.209
R49731 vdd.n12263 vdd.n10960 3.209
R49732 vdd.n12210 vdd.n12209 3.209
R49733 vdd.n12150 vdd.n11138 3.209
R49734 vdd.n12105 vdd.n12104 3.209
R49735 vdd.n12047 vdd.n12046 3.209
R49736 vdd.n12011 vdd.n11375 3.209
R49737 vdd.n11957 vdd.n11445 3.209
R49738 vdd.t190 vdd.n11944 3.209
R49739 vdd.n11660 vdd.n11565 3.209
R49740 vdd.n15457 vdd.n15456 3.209
R49741 vdd.n15625 vdd.n15624 3.209
R49742 vdd.n15214 vdd.n15213 3.209
R49743 vdd.n15713 vdd.n15712 3.209
R49744 vdd.n15881 vdd.n15880 3.209
R49745 vdd.n15969 vdd.n15968 3.209
R49746 vdd.n16137 vdd.n16136 3.209
R49747 vdd.n16225 vdd.n16224 3.209
R49748 vdd.n16393 vdd.n16392 3.209
R49749 vdd.n15130 vdd.n15129 3.209
R49750 vdd.n16481 vdd.n16480 3.209
R49751 vdd.n16626 vdd.n16625 3.209
R49752 vdd.n16661 vdd.n16658 3.209
R49753 vdd.n16899 vdd.n16898 3.209
R49754 vdd.n17055 vdd.n17054 3.209
R49755 vdd.n17171 vdd.n17170 3.209
R49756 vdd.n17327 vdd.n17326 3.209
R49757 vdd.n17443 vdd.n17442 3.209
R49758 vdd.n17596 vdd.n16827 3.209
R49759 vdd.n17701 vdd.n17700 3.209
R49760 vdd.n17857 vdd.n17856 3.209
R49761 vdd.n17972 vdd.n17971 3.209
R49762 vdd.n18128 vdd.n18127 3.209
R49763 vdd.n18242 vdd.n18241 3.209
R49764 vdd.n15023 vdd.n15022 3.209
R49765 vdd.n15009 vdd.t220 3.209
R49766 vdd.n21709 vdd.n21708 3.209
R49767 vdd.n15380 vdd.n15379 3.202
R49768 vdd.n32099 vdd.n32098 3.2
R49769 vdd.n13198 vdd.n9213 3.198
R49770 vdd.n13162 vdd.n9222 3.198
R49771 vdd.n240 vdd.n239 3.197
R49772 vdd.n33732 vdd.n33731 3.195
R49773 vdd.n933 vdd.n932 3.195
R49774 vdd.n25620 vdd.n25619 3.195
R49775 vdd.n30316 vdd.n30315 3.168
R49776 vdd.n31769 vdd.n31768 3.142
R49777 vdd.n35897 vdd.n35896 3.129
R49778 vdd.n35946 vdd.n35945 3.129
R49779 vdd.n36128 vdd.n36127 3.129
R49780 vdd.n36177 vdd.n36176 3.129
R49781 vdd.n36359 vdd.n36358 3.129
R49782 vdd.n36408 vdd.n36407 3.129
R49783 vdd.n36590 vdd.n36589 3.129
R49784 vdd.n36639 vdd.n36638 3.129
R49785 vdd.n36821 vdd.n36820 3.129
R49786 vdd.n36870 vdd.n36869 3.129
R49787 vdd.n37056 vdd.n37055 3.129
R49788 vdd.n37095 vdd.n37094 3.129
R49789 vdd.n2156 vdd.n2155 3.129
R49790 vdd.n33057 vdd.n33056 3.129
R49791 vdd.n32927 vdd.n32926 3.129
R49792 vdd.n37468 vdd.n37467 3.129
R49793 vdd.n38150 vdd.n38149 3.129
R49794 vdd.n38107 vdd.n38106 3.129
R49795 vdd.n37925 vdd.n37924 3.129
R49796 vdd.n37876 vdd.n37875 3.129
R49797 vdd.n37694 vdd.n37693 3.129
R49798 vdd.n37645 vdd.n37644 3.129
R49799 vdd.n28318 vdd.n28317 3.129
R49800 vdd.n28367 vdd.n28366 3.129
R49801 vdd.n28549 vdd.n28548 3.129
R49802 vdd.n28598 vdd.n28597 3.129
R49803 vdd.n28780 vdd.n28779 3.129
R49804 vdd.n28163 vdd.n28162 3.129
R49805 vdd.n31846 vdd.n31842 3.129
R49806 vdd.n29028 vdd.n29027 3.129
R49807 vdd.n29870 vdd.n29869 3.129
R49808 vdd.n29836 vdd.n29835 3.129
R49809 vdd.n31094 vdd.n31090 3.129
R49810 vdd.n30545 vdd.n30544 3.129
R49811 vdd.n10475 vdd.n10271 3.105
R49812 vdd.n15259 vdd.n15258 3.105
R49813 vdd.n33632 vdd.n33631 3.105
R49814 vdd.n33319 vdd.n33318 3.105
R49815 vdd.n33409 vdd.n33408 3.105
R49816 vdd.n34283 vdd.n34282 3.105
R49817 vdd.n33916 vdd.n33915 3.105
R49818 vdd.n34395 vdd.n34394 3.105
R49819 vdd.n34002 vdd.n34001 3.105
R49820 vdd.n35164 vdd.n35163 3.105
R49821 vdd.n35062 vdd.n35061 3.105
R49822 vdd.n35411 vdd.n35410 3.105
R49823 vdd.n35549 vdd.n35548 3.105
R49824 vdd.n34919 vdd.n34918 3.105
R49825 vdd.n34475 vdd.n34474 3.105
R49826 vdd.n34815 vdd.n34814 3.105
R49827 vdd.n34584 vdd.n34583 3.105
R49828 vdd.n1089 vdd.n1088 3.105
R49829 vdd.n629 vdd.n628 3.105
R49830 vdd.n733 vdd.n732 3.105
R49831 vdd.n131 vdd.n130 3.105
R49832 vdd.n424 vdd.n423 3.105
R49833 vdd.n529 vdd.n528 3.105
R49834 vdd.n6295 vdd.n6294 3.105
R49835 vdd.n6190 vdd.n6189 3.105
R49836 vdd.n6108 vdd.n6107 3.105
R49837 vdd.n5962 vdd.n5961 3.105
R49838 vdd.n5666 vdd.n5665 3.105
R49839 vdd.n5222 vdd.n5221 3.105
R49840 vdd.n5562 vdd.n5561 3.105
R49841 vdd.n5331 vdd.n5330 3.105
R49842 vdd.n4646 vdd.n4645 3.105
R49843 vdd.n4738 vdd.n4737 3.105
R49844 vdd.n4993 vdd.n4992 3.105
R49845 vdd.n5122 vdd.n5121 3.105
R49846 vdd.n4493 vdd.n4492 3.105
R49847 vdd.n4052 vdd.n4051 3.105
R49848 vdd.n4388 vdd.n4387 3.105
R49849 vdd.n4162 vdd.n4161 3.105
R49850 vdd.n27424 vdd.n27423 3.105
R49851 vdd.n27507 vdd.n27506 3.105
R49852 vdd.n27530 vdd.n27529 3.105
R49853 vdd.n27635 vdd.n27634 3.105
R49854 vdd.n25870 vdd.n25869 3.105
R49855 vdd.n25944 vdd.n25943 3.105
R49856 vdd.n25967 vdd.n25966 3.105
R49857 vdd.n26056 vdd.n26055 3.105
R49858 vdd.n10684 vdd.n10680 3.1
R49859 vdd.n12332 vdd.n12331 3.1
R49860 vdd.n11032 vdd.n11031 3.1
R49861 vdd.n12126 vdd.n12125 3.1
R49862 vdd.n12026 vdd.n12025 3.1
R49863 vdd.n17127 vdd.n17126 3.1
R49864 vdd.n17399 vdd.n17398 3.1
R49865 vdd.n17657 vdd.n17656 3.1
R49866 vdd.n17928 vdd.n17927 3.1
R49867 vdd.n18200 vdd.n18199 3.1
R49868 vdd.n24626 vdd.n24625 3.096
R49869 vdd.n33600 vdd.n33599 3.09
R49870 vdd.n1111 vdd.n1110 3.09
R49871 vdd.n24990 vdd.n24989 3.089
R49872 vdd.n25256 vdd.n25255 3.086
R49873 vdd.n10463 vdd.n10462 3.081
R49874 vdd.n10462 vdd.n10282 3.081
R49875 vdd.n10433 vdd.n10300 3.081
R49876 vdd.n10433 vdd.n10305 3.081
R49877 vdd.n13052 vdd.n9313 3.081
R49878 vdd.n13052 vdd.n9314 3.081
R49879 vdd.n9376 vdd.n9374 3.081
R49880 vdd.n9376 vdd.n9370 3.081
R49881 vdd.n12952 vdd.n12951 3.081
R49882 vdd.n12951 vdd.n9479 3.081
R49883 vdd.n12926 vdd.n9528 3.081
R49884 vdd.n12926 vdd.n9529 3.081
R49885 vdd.n12844 vdd.n9674 3.081
R49886 vdd.n12844 vdd.n9675 3.081
R49887 vdd.n9736 vdd.n9734 3.081
R49888 vdd.n9736 vdd.n9730 3.081
R49889 vdd.n12744 vdd.n12743 3.081
R49890 vdd.n12743 vdd.n9839 3.081
R49891 vdd.n12718 vdd.n9889 3.081
R49892 vdd.n12718 vdd.n9890 3.081
R49893 vdd.n12636 vdd.n10034 3.081
R49894 vdd.n12636 vdd.n10035 3.081
R49895 vdd.n10543 vdd.n10542 3.081
R49896 vdd.n10575 vdd.n10568 3.081
R49897 vdd.n12474 vdd.n10603 3.081
R49898 vdd.n12439 vdd.n12438 3.081
R49899 vdd.n12417 vdd.n10676 3.081
R49900 vdd.n12392 vdd.n12391 3.081
R49901 vdd.n10788 vdd.n10787 3.081
R49902 vdd.n10841 vdd.n10833 3.081
R49903 vdd.n10882 vdd.n10876 3.081
R49904 vdd.n10930 vdd.n10901 3.081
R49905 vdd.n12275 vdd.n12274 3.081
R49906 vdd.n12244 vdd.n11000 3.081
R49907 vdd.n12218 vdd.n11038 3.081
R49908 vdd.n12189 vdd.n11084 3.081
R49909 vdd.n12171 vdd.n11109 3.081
R49910 vdd.n12141 vdd.n11150 3.081
R49911 vdd.n11215 vdd.n11195 3.081
R49912 vdd.n11262 vdd.n11247 3.081
R49913 vdd.n11297 vdd.n11296 3.081
R49914 vdd.n11350 vdd.n11342 3.081
R49915 vdd.n11391 vdd.n11385 3.081
R49916 vdd.n11474 vdd.n11410 3.081
R49917 vdd.n11969 vdd.n11968 3.081
R49918 vdd.n11586 vdd.n11558 3.081
R49919 vdd.n15289 vdd.n15282 3.081
R49920 vdd.n15291 vdd.n15289 3.081
R49921 vdd.n15341 vdd.n15340 3.081
R49922 vdd.n15340 vdd.n15333 3.081
R49923 vdd.n15514 vdd.n15504 3.081
R49924 vdd.n15516 vdd.n15514 3.081
R49925 vdd.n15578 vdd.n15577 3.081
R49926 vdd.n15577 vdd.n15567 3.081
R49927 vdd.n15770 vdd.n15760 3.081
R49928 vdd.n15772 vdd.n15770 3.081
R49929 vdd.n15834 vdd.n15833 3.081
R49930 vdd.n15833 vdd.n15823 3.081
R49931 vdd.n16026 vdd.n16016 3.081
R49932 vdd.n16028 vdd.n16026 3.081
R49933 vdd.n16090 vdd.n16089 3.081
R49934 vdd.n16089 vdd.n16079 3.081
R49935 vdd.n16282 vdd.n16272 3.081
R49936 vdd.n16284 vdd.n16282 3.081
R49937 vdd.n16346 vdd.n16345 3.081
R49938 vdd.n16345 vdd.n16335 3.081
R49939 vdd.n16538 vdd.n16528 3.081
R49940 vdd.n16540 vdd.n16538 3.081
R49941 vdd.n16886 vdd.n16885 3.081
R49942 vdd.n16940 vdd.n16939 3.081
R49943 vdd.n17000 vdd.n16999 3.081
R49944 vdd.n17091 vdd.n17089 3.081
R49945 vdd.n17158 vdd.n17157 3.081
R49946 vdd.n17212 vdd.n17211 3.081
R49947 vdd.n17272 vdd.n17271 3.081
R49948 vdd.n17363 vdd.n17361 3.081
R49949 vdd.n17430 vdd.n17429 3.081
R49950 vdd.n17484 vdd.n17483 3.081
R49951 vdd.n17544 vdd.n17543 3.081
R49952 vdd.n17621 vdd.n17619 3.081
R49953 vdd.n17688 vdd.n17687 3.081
R49954 vdd.n17742 vdd.n17741 3.081
R49955 vdd.n17802 vdd.n17801 3.081
R49956 vdd.n17892 vdd.n17890 3.081
R49957 vdd.n17959 vdd.n17958 3.081
R49958 vdd.n18013 vdd.n18012 3.081
R49959 vdd.n18073 vdd.n18072 3.081
R49960 vdd.n18164 vdd.n18162 3.081
R49961 vdd.n18230 vdd.n18229 3.081
R49962 vdd.n18281 vdd.n18280 3.081
R49963 vdd.n18320 vdd.n18319 3.081
R49964 vdd.n18413 vdd.n18411 3.081
R49965 vdd.n9158 vdd.n9150 3.058
R49966 vdd.n9089 vdd.n9071 3.058
R49967 vdd.n13492 vdd.n8993 3.058
R49968 vdd.n13455 vdd.n9002 3.058
R49969 vdd.n13556 vdd.t283 3.058
R49970 vdd.n8936 vdd.n8929 3.058
R49971 vdd.n8869 vdd.n8851 3.058
R49972 vdd.n13746 vdd.n8785 3.058
R49973 vdd.n8721 vdd.n8719 3.058
R49974 vdd.n13934 vdd.n8619 3.058
R49975 vdd.n14051 vdd.n14050 3.058
R49976 vdd.n14038 vdd.n8576 3.058
R49977 vdd.n14224 vdd.n8397 3.058
R49978 vdd.n14326 vdd.n14325 3.058
R49979 vdd.n14372 vdd.n8317 3.058
R49980 vdd.n14437 vdd.n8241 3.058
R49981 vdd.n14531 vdd.n8197 3.058
R49982 vdd.n14646 vdd.n14645 3.058
R49983 vdd.n9995 vdd.n9994 3.049
R49984 vdd.n12684 vdd.n9963 3.049
R49985 vdd.n9807 vdd.n9780 3.049
R49986 vdd.n9806 vdd.n9785 3.049
R49987 vdd.n9635 vdd.n9634 3.049
R49988 vdd.n12892 vdd.n9603 3.049
R49989 vdd.n9448 vdd.n9419 3.049
R49990 vdd.n9447 vdd.n9425 3.049
R49991 vdd.n10376 vdd.n10350 3.049
R49992 vdd.n10349 vdd.n10346 3.049
R49993 vdd.n16436 vdd.n15136 3.049
R49994 vdd.n16435 vdd.n15150 3.049
R49995 vdd.n16180 vdd.n15164 3.049
R49996 vdd.n16179 vdd.n15178 3.049
R49997 vdd.n15924 vdd.n15180 3.049
R49998 vdd.n15923 vdd.n15206 3.049
R49999 vdd.n15668 vdd.n15220 3.049
R50000 vdd.n15667 vdd.n15234 3.049
R50001 vdd.n15418 vdd.n15245 3.049
R50002 vdd.n15417 vdd.n15256 3.049
R50003 vdd.n2619 vdd.n2618 3.041
R50004 vdd.n2236 vdd.n2235 3.041
R50005 vdd.n3949 vdd.n3948 3.041
R50006 vdd.n253 vdd.n251 3.033
R50007 vdd.n4824 vdd.n4822 3.033
R50008 vdd.n27290 vdd.n27289 3.033
R50009 vdd.n27272 vdd.n27271 3.033
R50010 vdd.n27594 vdd.n27593 3.033
R50011 vdd.n25833 vdd.n25832 3.033
R50012 vdd.n25709 vdd.n25708 3.033
R50013 vdd.n26010 vdd.n26009 3.033
R50014 vdd.n25458 vdd.n25457 3.033
R50015 vdd.n25612 vdd.n25611 3.033
R50016 vdd.n25603 vdd.n25602 3.033
R50017 vdd.n25668 vdd.n25667 3.033
R50018 vdd.n30207 vdd.n30206 3.033
R50019 vdd.n29891 vdd.n29890 3.033
R50020 vdd.n27988 vdd.n27987 3.033
R50021 vdd.n28981 vdd.n28980 3.033
R50022 vdd.n33582 vdd.n33581 3.033
R50023 vdd.n33511 vdd.n33510 3.033
R50024 vdd.n33459 vdd.n33458 3.033
R50025 vdd.n34116 vdd.n34115 3.033
R50026 vdd.n34431 vdd.n34430 3.033
R50027 vdd.n34068 vdd.n34067 3.033
R50028 vdd.n35472 vdd.n35471 3.033
R50029 vdd.n35389 vdd.n35388 3.033
R50030 vdd.n35229 vdd.n35228 3.033
R50031 vdd.n34950 vdd.n34949 3.033
R50032 vdd.n34861 vdd.n34860 3.033
R50033 vdd.n34642 vdd.n34641 3.033
R50034 vdd.n925 vdd.n924 3.033
R50035 vdd.n1035 vdd.n1034 3.033
R50036 vdd.n778 vdd.n777 3.033
R50037 vdd.n204 vdd.n203 3.033
R50038 vdd.n473 vdd.n472 3.033
R50039 vdd.n5824 vdd.n5823 3.033
R50040 vdd.n6082 vdd.n6081 3.033
R50041 vdd.n6352 vdd.n6351 3.033
R50042 vdd.n5697 vdd.n5696 3.033
R50043 vdd.n5608 vdd.n5607 3.033
R50044 vdd.n5389 vdd.n5388 3.033
R50045 vdd.n5183 vdd.n5182 3.033
R50046 vdd.n4723 vdd.n4722 3.033
R50047 vdd.n4524 vdd.n4523 3.033
R50048 vdd.n4435 vdd.n4434 3.033
R50049 vdd.n4219 vdd.n4218 3.033
R50050 vdd.n27884 vdd.n27883 3.033
R50051 vdd.n11595 vdd.n11586 3.033
R50052 vdd.n11950 vdd.n11949 3.033
R50053 vdd.n11967 vdd.n11435 3.033
R50054 vdd.n11864 vdd.n11812 3.033
R50055 vdd.n22374 vdd.n22373 3.033
R50056 vdd.n24319 vdd.n24318 3.033
R50057 vdd.n18414 vdd.n18413 3.033
R50058 vdd.n18388 vdd.n18387 3.033
R50059 vdd.n18330 vdd.n18329 3.033
R50060 vdd.n21955 vdd.n21903 3.033
R50061 vdd.n11744 vdd.n11724 3.027
R50062 vdd.n21826 vdd.n21806 3.027
R50063 vdd.n11885 vdd.n11800 3.027
R50064 vdd.n21976 vdd.n21891 3.027
R50065 vdd.n31496 vdd.n31495 3.024
R50066 vdd.n31649 vdd.n31648 3.024
R50067 vdd.n32427 vdd.n32426 3.024
R50068 vdd.n26172 vdd.n26171 3.024
R50069 vdd.n33521 vdd.n33520 3.011
R50070 vdd.n33980 vdd.n33979 3.011
R50071 vdd.n33896 vdd.n33895 3.011
R50072 vdd.n35142 vdd.n35141 3.011
R50073 vdd.n35090 vdd.n35089 3.011
R50074 vdd.n34555 vdd.n34554 3.011
R50075 vdd.n34503 vdd.n34502 3.011
R50076 vdd.n1002 vdd.n1001 3.011
R50077 vdd.n364 vdd.n363 3.011
R50078 vdd.n269 vdd.n268 3.011
R50079 vdd.n6265 vdd.n6264 3.011
R50080 vdd.n6170 vdd.n6169 3.011
R50081 vdd.n5302 vdd.n5301 3.011
R50082 vdd.n5250 vdd.n5249 3.011
R50083 vdd.n4978 vdd.n4977 3.011
R50084 vdd.n5159 vdd.n5158 3.011
R50085 vdd.n4132 vdd.n4131 3.011
R50086 vdd.n4080 vdd.n4079 3.011
R50087 vdd.n31586 vdd.n31585 3.011
R50088 vdd.n31156 vdd.n31152 3.011
R50089 vdd.n30341 vdd.n30334 3.011
R50090 vdd.n35857 vdd.n35850 3.011
R50091 vdd.n35990 vdd.n35983 3.011
R50092 vdd.n36088 vdd.n36081 3.011
R50093 vdd.n36221 vdd.n36214 3.011
R50094 vdd.n36319 vdd.n36312 3.011
R50095 vdd.n36452 vdd.n36445 3.011
R50096 vdd.n36550 vdd.n36543 3.011
R50097 vdd.n36683 vdd.n36676 3.011
R50098 vdd.n36781 vdd.n36774 3.011
R50099 vdd.n36914 vdd.n36907 3.011
R50100 vdd.n37021 vdd.n37017 3.011
R50101 vdd.n33197 vdd.n33190 3.011
R50102 vdd.n37206 vdd.n37199 3.011
R50103 vdd.n33013 vdd.n33009 3.011
R50104 vdd.n32961 vdd.n32954 3.011
R50105 vdd.n37509 vdd.n37505 3.011
R50106 vdd.n38196 vdd.n38192 3.011
R50107 vdd.n38067 vdd.n38060 3.011
R50108 vdd.n37969 vdd.n37962 3.011
R50109 vdd.n37836 vdd.n37829 3.011
R50110 vdd.n37738 vdd.n37731 3.011
R50111 vdd.n37605 vdd.n37598 3.011
R50112 vdd.n28278 vdd.n28271 3.011
R50113 vdd.n28411 vdd.n28404 3.011
R50114 vdd.n28509 vdd.n28502 3.011
R50115 vdd.n28642 vdd.n28635 3.011
R50116 vdd.n28740 vdd.n28733 3.011
R50117 vdd.n28065 vdd.n28058 3.011
R50118 vdd.n27938 vdd.n27937 3.011
R50119 vdd.n29876 vdd.n29875 3.011
R50120 vdd.n29857 vdd.n29856 3.011
R50121 vdd.n29858 vdd.n29857 3.011
R50122 vdd.n29765 vdd.n29758 3.011
R50123 vdd.n27553 vdd.n27552 3.011
R50124 vdd.n27258 vdd.n27257 3.011
R50125 vdd.n25990 vdd.n25989 3.011
R50126 vdd.n26026 vdd.n26025 3.011
R50127 vdd.n26754 vdd.n26750 3.011
R50128 vdd.n1273 vdd.n1266 3.011
R50129 vdd.n1692 vdd.n1688 3.011
R50130 vdd.n1616 vdd.n1612 3.011
R50131 vdd.n1511 vdd.n1507 3.011
R50132 vdd.n1435 vdd.n1431 3.011
R50133 vdd.n1330 vdd.n1326 3.011
R50134 vdd.n26796 vdd.n26792 3.011
R50135 vdd.n26901 vdd.n26897 3.011
R50136 vdd.n26977 vdd.n26973 3.011
R50137 vdd.n27082 vdd.n27078 3.011
R50138 vdd.n27158 vdd.n27154 3.011
R50139 vdd.n1878 vdd.n1877 3.011
R50140 vdd.n2575 vdd.n2573 3.011
R50141 vdd.n3787 vdd.n3786 3.011
R50142 vdd.n2749 vdd.n2745 3.011
R50143 vdd.n2854 vdd.n2850 3.011
R50144 vdd.n2930 vdd.n2926 3.011
R50145 vdd.n3035 vdd.n3031 3.011
R50146 vdd.n3111 vdd.n3107 3.011
R50147 vdd.n3216 vdd.n3212 3.011
R50148 vdd.n3292 vdd.n3288 3.011
R50149 vdd.n3397 vdd.n3393 3.011
R50150 vdd.n3473 vdd.n3469 3.011
R50151 vdd.n3578 vdd.n3574 3.011
R50152 vdd.n3635 vdd.n3628 3.011
R50153 vdd.n13129 vdd.n13128 3.011
R50154 vdd.n13128 vdd.n9269 3.011
R50155 vdd.n13295 vdd.n9146 3.011
R50156 vdd.n13295 vdd.n9101 3.011
R50157 vdd.n13423 vdd.n13422 3.011
R50158 vdd.n13422 vdd.n9038 3.011
R50159 vdd.n13587 vdd.n8925 3.011
R50160 vdd.n13587 vdd.n8880 3.011
R50161 vdd.n13715 vdd.n13714 3.011
R50162 vdd.n13714 vdd.n8817 3.011
R50163 vdd.n13891 vdd.n8686 3.011
R50164 vdd.n13891 vdd.n8691 3.011
R50165 vdd.n14060 vdd.n14059 3.011
R50166 vdd.n14059 vdd.n8569 3.011
R50167 vdd.n14180 vdd.n8462 3.011
R50168 vdd.n14180 vdd.n8468 3.011
R50169 vdd.n14335 vdd.n14334 3.011
R50170 vdd.n14334 vdd.n8351 3.011
R50171 vdd.n8255 vdd.n8254 3.011
R50172 vdd.n8254 vdd.n8220 3.011
R50173 vdd.n14664 vdd.n8138 3.011
R50174 vdd.n14669 vdd.n8136 3.011
R50175 vdd.n14726 vdd.n14725 3.011
R50176 vdd.n14751 vdd.n14750 3.011
R50177 vdd.n14836 vdd.n8048 3.011
R50178 vdd.n14841 vdd.n8046 3.011
R50179 vdd.n14918 vdd.n14917 3.011
R50180 vdd.n14924 vdd.n14923 3.011
R50181 vdd.n9260 vdd.n9259 3.011
R50182 vdd.n13155 vdd.n9237 3.011
R50183 vdd.n13170 vdd.n13168 3.011
R50184 vdd.n13170 vdd.n9227 3.011
R50185 vdd.n13332 vdd.n13331 3.011
R50186 vdd.n13331 vdd.n9109 3.011
R50187 vdd.n13470 vdd.n9006 3.011
R50188 vdd.n13470 vdd.n9007 3.011
R50189 vdd.n13624 vdd.n13623 3.011
R50190 vdd.n13623 vdd.n8888 3.011
R50191 vdd.n8788 vdd.n8757 3.011
R50192 vdd.n13801 vdd.n8757 3.011
R50193 vdd.n13925 vdd.n13924 3.011
R50194 vdd.n13924 vdd.n8650 3.011
R50195 vdd.n14032 vdd.n8544 3.011
R50196 vdd.n14088 vdd.n8544 3.011
R50197 vdd.n14215 vdd.n14214 3.011
R50198 vdd.n14214 vdd.n8430 3.011
R50199 vdd.n14364 vdd.n8322 3.011
R50200 vdd.n14364 vdd.n8325 3.011
R50201 vdd.n14484 vdd.n14483 3.011
R50202 vdd.n14483 vdd.n8228 3.011
R50203 vdd.n24239 vdd.n24238 3.011
R50204 vdd.n24248 vdd.n24247 3.011
R50205 vdd.n24138 vdd.n24137 3.011
R50206 vdd.n24028 vdd.n24027 3.011
R50207 vdd.n23906 vdd.n23905 3.011
R50208 vdd.n23796 vdd.n23795 3.011
R50209 vdd.n23674 vdd.n23673 3.011
R50210 vdd.n23108 vdd.n23107 3.011
R50211 vdd.n23218 vdd.n23217 3.011
R50212 vdd.n23340 vdd.n23339 3.011
R50213 vdd.n23450 vdd.n23449 3.011
R50214 vdd.n23572 vdd.n23571 3.011
R50215 vdd.n22529 vdd.n22528 3.011
R50216 vdd.n22639 vdd.n22638 3.011
R50217 vdd.n22761 vdd.n22760 3.011
R50218 vdd.n22871 vdd.n22870 3.011
R50219 vdd.n22993 vdd.n22992 3.011
R50220 vdd.n22411 vdd.n22410 3.011
R50221 vdd.n22420 vdd.n22419 3.011
R50222 vdd.n22228 vdd.n22217 3.011
R50223 vdd.n22219 vdd.n22218 3.011
R50224 vdd.n24356 vdd.n24355 3.011
R50225 vdd.n24365 vdd.n24364 3.011
R50226 vdd.n22104 vdd.n22093 3.011
R50227 vdd.n22095 vdd.n22094 3.011
R50228 vdd.n19353 vdd.n19344 3.011
R50229 vdd.n19498 vdd.n19489 3.011
R50230 vdd.n19559 vdd.n19550 3.011
R50231 vdd.n19698 vdd.n19689 3.011
R50232 vdd.n19761 vdd.n19752 3.011
R50233 vdd.n20958 vdd.n20949 3.011
R50234 vdd.n20895 vdd.n20886 3.011
R50235 vdd.n20768 vdd.n20759 3.011
R50236 vdd.n20707 vdd.n20698 3.011
R50237 vdd.n20562 vdd.n20553 3.011
R50238 vdd.n21627 vdd.n21626 3.011
R50239 vdd.n21578 vdd.n21569 3.011
R50240 vdd.n21464 vdd.n21455 3.011
R50241 vdd.n21319 vdd.n21310 3.011
R50242 vdd.n21205 vdd.n21196 3.011
R50243 vdd.n21060 vdd.n21051 3.011
R50244 vdd.n19098 vdd.n19089 3.011
R50245 vdd.n18953 vdd.n18944 3.011
R50246 vdd.n18839 vdd.n18830 3.011
R50247 vdd.n18694 vdd.n18685 3.011
R50248 vdd.n18580 vdd.n18571 3.011
R50249 vdd.n20445 vdd.n20444 3.011
R50250 vdd.n20323 vdd.n20322 3.011
R50251 vdd.n20209 vdd.n20208 3.011
R50252 vdd.n20087 vdd.n20086 3.011
R50253 vdd.n24699 vdd.n24698 3.011
R50254 vdd.n24788 vdd.n24787 3.011
R50255 vdd.n25206 vdd.n25205 3.011
R50256 vdd.n25117 vdd.n25116 3.011
R50257 vdd.n33699 vdd.n33574 2.953
R50258 vdd.n33572 vdd.n33476 2.953
R50259 vdd.n33364 vdd.n33289 2.953
R50260 vdd.n34158 vdd.n34075 2.953
R50261 vdd.n34341 vdd.n34239 2.953
R50262 vdd.n34345 vdd.n34235 2.953
R50263 vdd.n34345 vdd.n34238 2.953
R50264 vdd.n34071 vdd.n33967 2.953
R50265 vdd.n34071 vdd.n33970 2.953
R50266 vdd.n35233 vdd.n35132 2.953
R50267 vdd.n35233 vdd.n35134 2.953
R50268 vdd.n35608 vdd.n35466 2.953
R50269 vdd.n35355 vdd.n35278 2.953
R50270 vdd.n34771 vdd.n34694 2.953
R50271 vdd.n35020 vdd.n34881 2.953
R50272 vdd.n35024 vdd.n34877 2.953
R50273 vdd.n35024 vdd.n34880 2.953
R50274 vdd.n34646 vdd.n34542 2.953
R50275 vdd.n34646 vdd.n34547 2.953
R50276 vdd.n1166 vdd.n1050 2.953
R50277 vdd.n1170 vdd.n1048 2.953
R50278 vdd.n683 vdd.n599 2.953
R50279 vdd.n208 vdd.n88 2.953
R50280 vdd.n574 vdd.n507 2.953
R50281 vdd.n6356 vdd.n6252 2.953
R50282 vdd.n6356 vdd.n6255 2.953
R50283 vdd.n6043 vdd.n5924 2.953
R50284 vdd.n5846 vdd.n5844 2.953
R50285 vdd.n5518 vdd.n5441 2.953
R50286 vdd.n5767 vdd.n5628 2.953
R50287 vdd.n5771 vdd.n5624 2.953
R50288 vdd.n5771 vdd.n5627 2.953
R50289 vdd.n5393 vdd.n5288 2.953
R50290 vdd.n5393 vdd.n5294 2.953
R50291 vdd.n4707 vdd.n4617 2.953
R50292 vdd.n5067 vdd.n5063 2.953
R50293 vdd.n5067 vdd.n5065 2.953
R50294 vdd.n4949 vdd.n4874 2.953
R50295 vdd.n4345 vdd.n4268 2.953
R50296 vdd.n4597 vdd.n4455 2.953
R50297 vdd.n4601 vdd.n4451 2.953
R50298 vdd.n4601 vdd.n4454 2.953
R50299 vdd.n4223 vdd.n4119 2.953
R50300 vdd.n4223 vdd.n4124 2.953
R50301 vdd.n28806 vdd.n28133 2.953
R50302 vdd.n29038 vdd.n29021 2.953
R50303 vdd.n27785 vdd.n27783 2.953
R50304 vdd.n29035 vdd.n29023 2.953
R50305 vdd.n29849 vdd.n29684 2.953
R50306 vdd.n29952 vdd.n29853 2.953
R50307 vdd.n27358 vdd.n27305 2.953
R50308 vdd.n27465 vdd.n27285 2.953
R50309 vdd.n27466 vdd.n27284 2.953
R50310 vdd.n27466 vdd.n27281 2.953
R50311 vdd.n27592 vdd.n27265 2.953
R50312 vdd.n27592 vdd.n27262 2.953
R50313 vdd.n25810 vdd.n25757 2.953
R50314 vdd.n25911 vdd.n25731 2.953
R50315 vdd.n25912 vdd.n25730 2.953
R50316 vdd.n25912 vdd.n25727 2.953
R50317 vdd.n26008 vdd.n25682 2.953
R50318 vdd.n26008 vdd.n25680 2.953
R50319 vdd.n25558 vdd.n25430 2.953
R50320 vdd.n25559 vdd.n25429 2.953
R50321 vdd.n25568 vdd.n25567 2.953
R50322 vdd.n29823 vdd.n29822 2.953
R50323 vdd.n28005 vdd.n27841 2.953
R50324 vdd.n28120 vdd.n28118 2.953
R50325 vdd.n33391 vdd.n33386 2.953
R50326 vdd.n33391 vdd.n33384 2.953
R50327 vdd.n35465 vdd.n35363 2.953
R50328 vdd.n35465 vdd.n35360 2.953
R50329 vdd.n705 vdd.n699 2.953
R50330 vdd.n705 vdd.n696 2.953
R50331 vdd.n503 vdd.n498 2.953
R50332 vdd.n503 vdd.n495 2.953
R50333 vdd.n6136 vdd.n6051 2.953
R50334 vdd.n6136 vdd.n6049 2.953
R50335 vdd.n4711 vdd.n4613 2.953
R50336 vdd.n4711 vdd.n4610 2.953
R50337 vdd.n22326 vdd.n22279 2.953
R50338 vdd.n22328 vdd.n22268 2.953
R50339 vdd.n24298 vdd.n22164 2.953
R50340 vdd.n24300 vdd.n22153 2.953
R50341 vdd.n22470 vdd.n22185 2.953
R50342 vdd.n19382 vdd.n19379 2.932
R50343 vdd.n19463 vdd.n19460 2.932
R50344 vdd.n19588 vdd.n19585 2.932
R50345 vdd.t154 vdd.n19634 2.932
R50346 vdd.n19663 vdd.n19660 2.932
R50347 vdd.n19790 vdd.n19787 2.932
R50348 vdd.n20987 vdd.n20984 2.932
R50349 vdd.n19889 vdd.n19886 2.932
R50350 vdd.t172 vdd.n20839 2.932
R50351 vdd.n20796 vdd.n20793 2.932
R50352 vdd.n20672 vdd.n20669 2.932
R50353 vdd.n20591 vdd.n20588 2.932
R50354 vdd.n20471 vdd.n20470 2.932
R50355 vdd.n20298 vdd.n20297 2.932
R50356 vdd.n20248 vdd.n20247 2.932
R50357 vdd.n20062 vdd.n20061 2.932
R50358 vdd.n14773 vdd.n8082 2.924
R50359 vdd.n14828 vdd.n8055 2.924
R50360 vdd.n14942 vdd.n8001 2.924
R50361 vdd.n11914 vdd.n11910 2.919
R50362 vdd.n22000 vdd.n21999 2.919
R50363 vdd.n36015 vdd.n36014 2.905
R50364 vdd.n36057 vdd.n36056 2.905
R50365 vdd.n36246 vdd.n36245 2.905
R50366 vdd.n36288 vdd.n36287 2.905
R50367 vdd.n36477 vdd.n36476 2.905
R50368 vdd.n36519 vdd.n36518 2.905
R50369 vdd.n36708 vdd.n36707 2.905
R50370 vdd.n36750 vdd.n36749 2.905
R50371 vdd.n36805 vdd.t39 2.905
R50372 vdd.n36939 vdd.n36938 2.905
R50373 vdd.n3642 vdd.n3641 2.905
R50374 vdd.n37147 vdd.n37146 2.905
R50375 vdd.n37175 vdd.n37174 2.905
R50376 vdd.n32988 vdd.n32987 2.905
R50377 vdd.n32974 vdd.n32973 2.905
R50378 vdd.n37522 vdd.n37521 2.905
R50379 vdd.n37568 vdd.n37567 2.905
R50380 vdd.n38036 vdd.n38035 2.905
R50381 vdd.n37994 vdd.n37993 2.905
R50382 vdd.n37805 vdd.n37804 2.905
R50383 vdd.n37763 vdd.n37762 2.905
R50384 vdd.n28205 vdd.n28204 2.905
R50385 vdd.n28247 vdd.n28246 2.905
R50386 vdd.n28436 vdd.n28435 2.905
R50387 vdd.n28478 vdd.n28477 2.905
R50388 vdd.n28610 vdd.t36 2.905
R50389 vdd.n28667 vdd.n28666 2.905
R50390 vdd.n28709 vdd.n28708 2.905
R50391 vdd.n28112 vdd.n28111 2.905
R50392 vdd.n28086 vdd.n28085 2.905
R50393 vdd.n31625 vdd.n31624 2.905
R50394 vdd.n32063 vdd.n32062 2.905
R50395 vdd.n29720 vdd.n29719 2.905
R50396 vdd.n30188 vdd.n30187 2.905
R50397 vdd.n10476 vdd.n10272 2.904
R50398 vdd.n10417 vdd.n10416 2.904
R50399 vdd.n15262 vdd.n15261 2.904
R50400 vdd.n13071 vdd.n9298 2.888
R50401 vdd.n13023 vdd.n9360 2.888
R50402 vdd.n9496 vdd.n9483 2.888
R50403 vdd.n9562 vdd.n9561 2.888
R50404 vdd.n12863 vdd.n9658 2.888
R50405 vdd.n12815 vdd.n9720 2.888
R50406 vdd.n9856 vdd.n9843 2.888
R50407 vdd.n9922 vdd.n9920 2.888
R50408 vdd.n12655 vdd.n10018 2.888
R50409 vdd.n12606 vdd.n10062 2.888
R50410 vdd.n12513 vdd.n10529 2.888
R50411 vdd.n12460 vdd.n12459 2.888
R50412 vdd.n12400 vdd.n10709 2.888
R50413 vdd.n12364 vdd.n10773 2.888
R50414 vdd.n12306 vdd.n12305 2.888
R50415 vdd.n10984 vdd.n10983 2.888
R50416 vdd.n11076 vdd.n11075 2.888
R50417 vdd.n11137 vdd.n11128 2.888
R50418 vdd.n11234 vdd.n11230 2.888
R50419 vdd.n12058 vdd.n11281 2.888
R50420 vdd.n12000 vdd.n11999 2.888
R50421 vdd.n11528 vdd.n11526 2.888
R50422 vdd.n15478 vdd.n15474 2.888
R50423 vdd.n15609 vdd.n15608 2.888
R50424 vdd.n15734 vdd.n15730 2.888
R50425 vdd.n15865 vdd.n15864 2.888
R50426 vdd.n15990 vdd.n15986 2.888
R50427 vdd.n16121 vdd.n16120 2.888
R50428 vdd.n16246 vdd.n16242 2.888
R50429 vdd.n16377 vdd.n16376 2.888
R50430 vdd.n16502 vdd.n16498 2.888
R50431 vdd.n16617 vdd.n16616 2.888
R50432 vdd.n16914 vdd.n16911 2.888
R50433 vdd.n17038 vdd.n17035 2.888
R50434 vdd.n17186 vdd.n17183 2.888
R50435 vdd.n17310 vdd.n17307 2.888
R50436 vdd.n17458 vdd.n17455 2.888
R50437 vdd.n17582 vdd.n17579 2.888
R50438 vdd.n17716 vdd.n17713 2.888
R50439 vdd.n17840 vdd.n17837 2.888
R50440 vdd.n17987 vdd.n17984 2.888
R50441 vdd.n18111 vdd.n18108 2.888
R50442 vdd.n18256 vdd.n18254 2.888
R50443 vdd.n18364 vdd.n18363 2.888
R50444 vdd.n15367 vdd.n15366 2.882
R50445 vdd.n28156 vdd.n28153 2.878
R50446 vdd.n38126 vdd.n38125 2.878
R50447 vdd.n1740 vdd.n1739 2.878
R50448 vdd.n13132 vdd.n9264 2.878
R50449 vdd.n13177 vdd.n9225 2.878
R50450 vdd.n1747 vdd.n1746 2.878
R50451 vdd.n26748 vdd.n26745 2.878
R50452 vdd.n38137 vdd.n38136 2.878
R50453 vdd.n28919 vdd.n28092 2.876
R50454 vdd.n24310 vdd.n22060 2.876
R50455 vdd.n24321 vdd.n22053 2.876
R50456 vdd.n24204 vdd.n22174 2.876
R50457 vdd.n22365 vdd.n22202 2.876
R50458 vdd.n22376 vdd.n22195 2.876
R50459 vdd.n10491 vdd.n10269 2.844
R50460 vdd.n10329 vdd.n10328 2.844
R50461 vdd.n10333 vdd.n10330 2.844
R50462 vdd.n10366 vdd.n10358 2.844
R50463 vdd.n10359 vdd.n9293 2.844
R50464 vdd.n13009 vdd.n9403 2.844
R50465 vdd.n13004 vdd.n9405 2.844
R50466 vdd.n12976 vdd.n9452 2.844
R50467 vdd.n12969 vdd.n9457 2.844
R50468 vdd.n9590 vdd.n9582 2.844
R50469 vdd.n9599 vdd.n9598 2.844
R50470 vdd.n9651 vdd.n9628 2.844
R50471 vdd.n9653 vdd.n9625 2.844
R50472 vdd.n12801 vdd.n9763 2.844
R50473 vdd.n12796 vdd.n9765 2.844
R50474 vdd.n12768 vdd.n9811 2.844
R50475 vdd.n12761 vdd.n9817 2.844
R50476 vdd.n9950 vdd.n9942 2.844
R50477 vdd.n9959 vdd.n9958 2.844
R50478 vdd.n10011 vdd.n9988 2.844
R50479 vdd.n10013 vdd.n9985 2.844
R50480 vdd.n10159 vdd.n10148 2.844
R50481 vdd.n10165 vdd.n10164 2.844
R50482 vdd.n10544 vdd.n10543 2.844
R50483 vdd.n12498 vdd.n12497 2.844
R50484 vdd.n10635 vdd.n10611 2.844
R50485 vdd.n12451 vdd.n12450 2.844
R50486 vdd.n12417 vdd.n10698 2.844
R50487 vdd.n10743 vdd.n10742 2.844
R50488 vdd.n10802 vdd.n10801 2.844
R50489 vdd.n12345 vdd.n10812 2.844
R50490 vdd.n10882 vdd.n10873 2.844
R50491 vdd.n12297 vdd.n12296 2.844
R50492 vdd.n10980 vdd.n10970 2.844
R50493 vdd.n12249 vdd.n10992 2.844
R50494 vdd.n11048 vdd.n11038 2.844
R50495 vdd.n12199 vdd.n11061 2.844
R50496 vdd.n12158 vdd.n11130 2.844
R50497 vdd.n11171 vdd.n11152 2.844
R50498 vdd.n12113 vdd.n11195 2.844
R50499 vdd.n11252 vdd.n11250 2.844
R50500 vdd.n11311 vdd.n11310 2.844
R50501 vdd.n12039 vdd.n11321 2.844
R50502 vdd.n11391 vdd.n11382 2.844
R50503 vdd.n11991 vdd.n11990 2.844
R50504 vdd.n15069 vdd.n15068 2.844
R50505 vdd.n15398 vdd.n15388 2.844
R50506 vdd.n15390 vdd.n15389 2.844
R50507 vdd.n15436 vdd.n15435 2.844
R50508 vdd.n15445 vdd.n15444 2.844
R50509 vdd.n15646 vdd.n15633 2.844
R50510 vdd.n15635 vdd.n15634 2.844
R50511 vdd.n15689 vdd.n15688 2.844
R50512 vdd.n15701 vdd.n15700 2.844
R50513 vdd.n15902 vdd.n15889 2.844
R50514 vdd.n15891 vdd.n15890 2.844
R50515 vdd.n15945 vdd.n15944 2.844
R50516 vdd.n15957 vdd.n15956 2.844
R50517 vdd.n16158 vdd.n16145 2.844
R50518 vdd.n16147 vdd.n16146 2.844
R50519 vdd.n16201 vdd.n16200 2.844
R50520 vdd.n16213 vdd.n16212 2.844
R50521 vdd.n16414 vdd.n16401 2.844
R50522 vdd.n16403 vdd.n16402 2.844
R50523 vdd.n16457 vdd.n16456 2.844
R50524 vdd.n16469 vdd.n16468 2.844
R50525 vdd.n16581 vdd.n16580 2.844
R50526 vdd.n16885 vdd.n16876 2.844
R50527 vdd.n16950 vdd.n16938 2.844
R50528 vdd.n17027 vdd.n17026 2.844
R50529 vdd.n17073 vdd.n17064 2.844
R50530 vdd.n17157 vdd.n17148 2.844
R50531 vdd.n17222 vdd.n17210 2.844
R50532 vdd.n17299 vdd.n17298 2.844
R50533 vdd.n17345 vdd.n17336 2.844
R50534 vdd.n17429 vdd.n17420 2.844
R50535 vdd.n17494 vdd.n17482 2.844
R50536 vdd.n17571 vdd.n17570 2.844
R50537 vdd.n17603 vdd.n16821 2.844
R50538 vdd.n17687 vdd.n17678 2.844
R50539 vdd.n17752 vdd.n17740 2.844
R50540 vdd.n17829 vdd.n17828 2.844
R50541 vdd.n17874 vdd.n17866 2.844
R50542 vdd.n17958 vdd.n17949 2.844
R50543 vdd.n18023 vdd.n18011 2.844
R50544 vdd.n18100 vdd.n18099 2.844
R50545 vdd.n18146 vdd.n18137 2.844
R50546 vdd.n18229 vdd.n18221 2.844
R50547 vdd.n18290 vdd.n18279 2.844
R50548 vdd.n12525 vdd.n10520 2.832
R50549 vdd.n16872 vdd.n16871 2.832
R50550 vdd.n33722 vdd.n33721 2.82
R50551 vdd.n886 vdd.n885 2.82
R50552 vdd.n31545 vdd.n31544 2.82
R50553 vdd.n21544 vdd.n21543 2.814
R50554 vdd.n21494 vdd.n21493 2.814
R50555 vdd.n21285 vdd.n21284 2.814
R50556 vdd.n21235 vdd.n21234 2.814
R50557 vdd.n21026 vdd.n21025 2.814
R50558 vdd.n19127 vdd.n19126 2.814
R50559 vdd.n18919 vdd.n18918 2.814
R50560 vdd.n18869 vdd.n18868 2.814
R50561 vdd.n18660 vdd.n18659 2.814
R50562 vdd.n18610 vdd.n18609 2.814
R50563 vdd.n28166 vdd.n28165 2.77
R50564 vdd.n26738 vdd.n26737 2.77
R50565 vdd.n13336 vdd.n9103 2.752
R50566 vdd.n13335 vdd.n9105 2.752
R50567 vdd.n13426 vdd.n9033 2.752
R50568 vdd.n13481 vdd.t116 2.752
R50569 vdd.n9004 vdd.n8988 2.752
R50570 vdd.n13521 vdd.t316 2.752
R50571 vdd.n13628 vdd.n8882 2.752
R50572 vdd.n13627 vdd.n8884 2.752
R50573 vdd.n13718 vdd.n8812 2.752
R50574 vdd.n13772 vdd.t288 2.752
R50575 vdd.n13803 vdd.n8754 2.752
R50576 vdd.n8695 vdd.n8694 2.752
R50577 vdd.n13927 vdd.t110 2.752
R50578 vdd.n14062 vdd.n8564 2.752
R50579 vdd.n14090 vdd.n8541 2.752
R50580 vdd.n8500 vdd.t132 2.752
R50581 vdd.t326 vdd.n8470 2.752
R50582 vdd.n8472 vdd.n8471 2.752
R50583 vdd.n14217 vdd.n8425 2.752
R50584 vdd.n14337 vdd.n8346 2.752
R50585 vdd.n14361 vdd.n14360 2.752
R50586 vdd.n14354 vdd.t333 2.752
R50587 vdd.t332 vdd.n8287 2.752
R50588 vdd.n14488 vdd.n8222 2.752
R50589 vdd.n14487 vdd.n8224 2.752
R50590 vdd.n14656 vdd.n8145 2.752
R50591 vdd.n14662 vdd.n8141 2.752
R50592 vdd.n99 vdd.n98 2.722
R50593 vdd.n28851 vdd.n28850 2.716
R50594 vdd.n35883 vdd.n35882 2.682
R50595 vdd.n35960 vdd.n35959 2.682
R50596 vdd.n36114 vdd.n36113 2.682
R50597 vdd.n36191 vdd.n36190 2.682
R50598 vdd.n36345 vdd.n36344 2.682
R50599 vdd.n36422 vdd.n36421 2.682
R50600 vdd.n36576 vdd.n36575 2.682
R50601 vdd.n36653 vdd.n36652 2.682
R50602 vdd.n36807 vdd.n36806 2.682
R50603 vdd.n36884 vdd.n36883 2.682
R50604 vdd.n2720 vdd.n2719 2.682
R50605 vdd.n33218 vdd.n33217 2.682
R50606 vdd.n2177 vdd.n2176 2.682
R50607 vdd.n37277 vdd.n37276 2.682
R50608 vdd.n37418 vdd.n37417 2.682
R50609 vdd.n37480 vdd.n37479 2.682
R50610 vdd.n38166 vdd.n38165 2.682
R50611 vdd.n38093 vdd.n38092 2.682
R50612 vdd.n37939 vdd.n37938 2.682
R50613 vdd.n37862 vdd.n37861 2.682
R50614 vdd.n37708 vdd.n37707 2.682
R50615 vdd.n37631 vdd.n37630 2.682
R50616 vdd.n28304 vdd.n28303 2.682
R50617 vdd.n28381 vdd.n28380 2.682
R50618 vdd.n28535 vdd.n28534 2.682
R50619 vdd.n28612 vdd.n28611 2.682
R50620 vdd.n28766 vdd.n28765 2.682
R50621 vdd.n28173 vdd.n28172 2.682
R50622 vdd.n28988 vdd.n28987 2.682
R50623 vdd.n27792 vdd.n27791 2.682
R50624 vdd.n31572 vdd.n31568 2.682
R50625 vdd.n29817 vdd.n29816 2.682
R50626 vdd.n30272 vdd.n30271 2.682
R50627 vdd.n31258 vdd.n31257 2.682
R50628 vdd.n11771 vdd.n11770 2.674
R50629 vdd.n21865 vdd.n21858 2.674
R50630 vdd.n11785 vdd.n11784 2.672
R50631 vdd.n21877 vdd.n21876 2.672
R50632 vdd.n242 vdd.n240 2.67
R50633 vdd.n11922 vdd.n11921 2.666
R50634 vdd.n13084 vdd.n9285 2.666
R50635 vdd.n15003 vdd.n15002 2.666
R50636 vdd.n21745 vdd.n21744 2.666
R50637 vdd.n11901 vdd.n11900 2.646
R50638 vdd.n21992 vdd.n21991 2.646
R50639 vdd.n28176 vdd.n28175 2.645
R50640 vdd.n31261 vdd.n31260 2.645
R50641 ldomc_0.otaldom_0.pcascodeupm_0.vdd vdd.n11906 2.639
R50642 vdd vdd.n21997 2.639
R50643 vdd.n11895 vdd.n11894 2.637
R50644 vdd.n21986 vdd.n21985 2.637
R50645 vdd.n33849 vdd.n33848 2.635
R50646 vdd.n33670 vdd.n33669 2.635
R50647 vdd.n34192 vdd.n34191 2.635
R50648 vdd.n34206 vdd.n34205 2.635
R50649 vdd.n35290 vdd.n35289 2.635
R50650 vdd.n35302 vdd.n35301 2.635
R50651 vdd.n34718 vdd.n34717 2.635
R50652 vdd.n34706 vdd.n34705 2.635
R50653 vdd.n850 vdd.n849 2.635
R50654 vdd.n1063 vdd.n1062 2.635
R50655 vdd.n5907 vdd.n5906 2.635
R50656 vdd.n5893 vdd.n5892 2.635
R50657 vdd.n5465 vdd.n5464 2.635
R50658 vdd.n5453 vdd.n5452 2.635
R50659 vdd.n4292 vdd.n4291 2.635
R50660 vdd.n4280 vdd.n4279 2.635
R50661 vdd.n30242 vdd.n30241 2.635
R50662 vdd.n31504 vdd.n31503 2.635
R50663 vdd.n31527 vdd.n31526 2.635
R50664 vdd.n31516 vdd.n31515 2.635
R50665 vdd.n32292 vdd.n32291 2.635
R50666 vdd.n31527 vdd.n31520 2.635
R50667 vdd.n32182 vdd.n32180 2.635
R50668 vdd.n32160 vdd.n32159 2.635
R50669 vdd.n32180 vdd.n32179 2.635
R50670 vdd.n32151 vdd.n32150 2.635
R50671 vdd.n31664 vdd.n31663 2.635
R50672 vdd.n31919 vdd.n31918 2.635
R50673 vdd.n31947 vdd.n31946 2.635
R50674 vdd.n31923 vdd.n31922 2.635
R50675 vdd.n31920 vdd.n31919 2.635
R50676 vdd.n32439 vdd.n32438 2.635
R50677 vdd.n32451 vdd.n32450 2.635
R50678 vdd.n31066 vdd.n31065 2.635
R50679 vdd.n31068 vdd.n31066 2.635
R50680 vdd.n31041 vdd.n31038 2.635
R50681 vdd.n31031 vdd.n31030 2.635
R50682 vdd.n31270 vdd.n31269 2.635
R50683 vdd.n30512 vdd.n30511 2.635
R50684 vdd.n35864 vdd.n35863 2.635
R50685 vdd.n35969 vdd.n35968 2.635
R50686 vdd.n36095 vdd.n36094 2.635
R50687 vdd.n36200 vdd.n36199 2.635
R50688 vdd.n36326 vdd.n36325 2.635
R50689 vdd.n36431 vdd.n36430 2.635
R50690 vdd.n36557 vdd.n36556 2.635
R50691 vdd.n36662 vdd.n36661 2.635
R50692 vdd.n36788 vdd.n36787 2.635
R50693 vdd.n36893 vdd.n36892 2.635
R50694 vdd.n37036 vdd.n37035 2.635
R50695 vdd.n37109 vdd.n37108 2.635
R50696 vdd.n33110 vdd.n33109 2.635
R50697 vdd.n33031 vdd.n33030 2.635
R50698 vdd.n37402 vdd.n37401 2.635
R50699 vdd.n32864 vdd.n32863 2.635
R50700 vdd.n38178 vdd.n38177 2.635
R50701 vdd.n38074 vdd.n38073 2.635
R50702 vdd.n37948 vdd.n37947 2.635
R50703 vdd.n37843 vdd.n37842 2.635
R50704 vdd.n37717 vdd.n37716 2.635
R50705 vdd.n37612 vdd.n37611 2.635
R50706 vdd.n28285 vdd.n28284 2.635
R50707 vdd.n28390 vdd.n28389 2.635
R50708 vdd.n28516 vdd.n28515 2.635
R50709 vdd.n28621 vdd.n28620 2.635
R50710 vdd.n28747 vdd.n28746 2.635
R50711 vdd.n28142 vdd.n28141 2.635
R50712 vdd.n28961 vdd.n28960 2.635
R50713 vdd.n28974 vdd.n28973 2.635
R50714 vdd.n27820 vdd.n27819 2.635
R50715 vdd.n27811 vdd.n27804 2.635
R50716 vdd.n27814 vdd.n27813 2.635
R50717 vdd.n27813 vdd.n27812 2.635
R50718 vdd.n29875 vdd.n29874 2.635
R50719 vdd.n30011 vdd.n30010 2.635
R50720 vdd.n29776 vdd.n29775 2.635
R50721 vdd.n27330 vdd.n27329 2.635
R50722 vdd.n27342 vdd.n27341 2.635
R50723 vdd.n25782 vdd.n25781 2.635
R50724 vdd.n25794 vdd.n25793 2.635
R50725 vdd.n25503 vdd.n25502 2.635
R50726 vdd.n25618 vdd.n25617 2.635
R50727 vdd.n27232 vdd.n27231 2.635
R50728 vdd.n26153 vdd.n26152 2.635
R50729 vdd.n1277 vdd.n1276 2.635
R50730 vdd.n1699 vdd.n1698 2.635
R50731 vdd.n1601 vdd.n1600 2.635
R50732 vdd.n1518 vdd.n1517 2.635
R50733 vdd.n1420 vdd.n1419 2.635
R50734 vdd.n1337 vdd.n1336 2.635
R50735 vdd.n26803 vdd.n26802 2.635
R50736 vdd.n26886 vdd.n26885 2.635
R50737 vdd.n26984 vdd.n26983 2.635
R50738 vdd.n27067 vdd.n27066 2.635
R50739 vdd.n27165 vdd.n27164 2.635
R50740 vdd.n1199 vdd.n1198 2.635
R50741 vdd.n1932 vdd.n1931 2.635
R50742 vdd.n1933 vdd.n1932 2.635
R50743 vdd.n2651 vdd.n2650 2.635
R50744 vdd.n2639 vdd.n2638 2.635
R50745 vdd.n2042 vdd.n2041 2.635
R50746 vdd.n2385 vdd.n2373 2.635
R50747 vdd.n2029 vdd.n2028 2.635
R50748 vdd.n2044 vdd.n2033 2.635
R50749 vdd.n2030 vdd.n2029 2.635
R50750 vdd.n2199 vdd.n2198 2.635
R50751 vdd.n2180 vdd.n2172 2.635
R50752 vdd.n2189 vdd.n2188 2.635
R50753 vdd.n3817 vdd.n3816 2.635
R50754 vdd.n2016 vdd.n2015 2.635
R50755 vdd.n3758 vdd.n3757 2.635
R50756 vdd.n2018 vdd.n2007 2.635
R50757 vdd.n2059 vdd.n2058 2.635
R50758 vdd.n2723 vdd.n2715 2.635
R50759 vdd.n2756 vdd.n2755 2.635
R50760 vdd.n2839 vdd.n2838 2.635
R50761 vdd.n2937 vdd.n2936 2.635
R50762 vdd.n3020 vdd.n3019 2.635
R50763 vdd.n3118 vdd.n3117 2.635
R50764 vdd.n3201 vdd.n3200 2.635
R50765 vdd.n3299 vdd.n3298 2.635
R50766 vdd.n3382 vdd.n3381 2.635
R50767 vdd.n3480 vdd.n3479 2.635
R50768 vdd.n3563 vdd.n3562 2.635
R50769 vdd.n2049 vdd.n2048 2.635
R50770 vdd.n31721 vdd.n31720 2.635
R50771 vdd.n31713 vdd.n31712 2.635
R50772 vdd.n31715 vdd.n31713 2.635
R50773 vdd.n13196 vdd.n9216 2.635
R50774 vdd.n13191 vdd.n9217 2.635
R50775 vdd.n13291 vdd.n13290 2.635
R50776 vdd.n13301 vdd.n13300 2.635
R50777 vdd.n13490 vdd.n8996 2.635
R50778 vdd.n13485 vdd.n8997 2.635
R50779 vdd.n13583 vdd.n13582 2.635
R50780 vdd.n13593 vdd.n13592 2.635
R50781 vdd.n13770 vdd.n8779 2.635
R50782 vdd.n13765 vdd.n8780 2.635
R50783 vdd.n13851 vdd.n13850 2.635
R50784 vdd.n13897 vdd.n13896 2.635
R50785 vdd.n14054 vdd.n8572 2.635
R50786 vdd.n14047 vdd.n14042 2.635
R50787 vdd.n14140 vdd.n14139 2.635
R50788 vdd.n14186 vdd.n14185 2.635
R50789 vdd.n14329 vdd.n8355 2.635
R50790 vdd.n14322 vdd.n14319 2.635
R50791 vdd.n14456 vdd.n14455 2.635
R50792 vdd.n8259 vdd.n8249 2.635
R50793 vdd.n8158 vdd.n8153 2.635
R50794 vdd.n8158 vdd.n8157 2.635
R50795 vdd.n14756 vdd.n8096 2.635
R50796 vdd.n14756 vdd.n8092 2.635
R50797 vdd.n14814 vdd.n14809 2.635
R50798 vdd.n14814 vdd.n14813 2.635
R50799 vdd.n14934 vdd.n8005 2.635
R50800 vdd.n14934 vdd.n8006 2.635
R50801 vdd.n13158 vdd.n9232 2.635
R50802 vdd.n9233 vdd.n9230 2.635
R50803 vdd.n9121 vdd.n9120 2.635
R50804 vdd.n9113 vdd.n9074 2.635
R50805 vdd.n13452 vdd.n9012 2.635
R50806 vdd.n13459 vdd.n13458 2.635
R50807 vdd.n8900 vdd.n8899 2.635
R50808 vdd.n8892 vdd.n8854 2.635
R50809 vdd.n13742 vdd.n8790 2.635
R50810 vdd.n13753 vdd.n8787 2.635
R50811 vdd.n13919 vdd.n8654 2.635
R50812 vdd.n13938 vdd.n8639 2.635
R50813 vdd.n14026 vdd.n8578 2.635
R50814 vdd.n14031 vdd.n8579 2.635
R50815 vdd.n14209 vdd.n8434 2.635
R50816 vdd.n14228 vdd.n8417 2.635
R50817 vdd.n14316 vdd.n8360 2.635
R50818 vdd.n14370 vdd.n14369 2.635
R50819 vdd.n14479 vdd.n8194 2.635
R50820 vdd.n14535 vdd.n14534 2.635
R50821 vdd.n24261 vdd.n24254 2.635
R50822 vdd.n24263 vdd.n24261 2.635
R50823 vdd.n24159 vdd.n24152 2.635
R50824 vdd.n24021 vdd.n24014 2.635
R50825 vdd.n23927 vdd.n23920 2.635
R50826 vdd.n23789 vdd.n23782 2.635
R50827 vdd.n23695 vdd.n23688 2.635
R50828 vdd.n23101 vdd.n23094 2.635
R50829 vdd.n23239 vdd.n23232 2.635
R50830 vdd.n23333 vdd.n23326 2.635
R50831 vdd.n23471 vdd.n23464 2.635
R50832 vdd.n23565 vdd.n23558 2.635
R50833 vdd.n22522 vdd.n22515 2.635
R50834 vdd.n22660 vdd.n22653 2.635
R50835 vdd.n22754 vdd.n22747 2.635
R50836 vdd.n22892 vdd.n22885 2.635
R50837 vdd.n22986 vdd.n22979 2.635
R50838 vdd.n22433 vdd.n22426 2.635
R50839 vdd.n22435 vdd.n22433 2.635
R50840 vdd.n22289 vdd.n22282 2.635
R50841 vdd.n22291 vdd.n22289 2.635
R50842 vdd.n19360 vdd.n19359 2.635
R50843 vdd.n19473 vdd.n19472 2.635
R50844 vdd.n19566 vdd.n19565 2.635
R50845 vdd.n19673 vdd.n19672 2.635
R50846 vdd.n19768 vdd.n19767 2.635
R50847 vdd.n20965 vdd.n20964 2.635
R50848 vdd.n20870 vdd.n20869 2.635
R50849 vdd.n20774 vdd.n20773 2.635
R50850 vdd.n20682 vdd.n20681 2.635
R50851 vdd.n20569 vdd.n20568 2.635
R50852 vdd.n21585 vdd.n21584 2.635
R50853 vdd.n21439 vdd.n21438 2.635
R50854 vdd.n21326 vdd.n21325 2.635
R50855 vdd.n21180 vdd.n21179 2.635
R50856 vdd.n21067 vdd.n21066 2.635
R50857 vdd.n19073 vdd.n19072 2.635
R50858 vdd.n18960 vdd.n18959 2.635
R50859 vdd.n18814 vdd.n18813 2.635
R50860 vdd.n18701 vdd.n18700 2.635
R50861 vdd.n18555 vdd.n18554 2.635
R50862 vdd.n20463 vdd.n20459 2.635
R50863 vdd.n20316 vdd.n20307 2.635
R50864 vdd.n20234 vdd.n20225 2.635
R50865 vdd.n20080 vdd.n20071 2.635
R50866 vdd.n24692 vdd.n24687 2.635
R50867 vdd.n24805 vdd.n24800 2.635
R50868 vdd.n25223 vdd.n25218 2.635
R50869 vdd.n25110 vdd.n25105 2.635
R50870 vdd.n11877 vdd.n11876 2.608
R50871 vdd.n21968 vdd.n21967 2.608
R50872 vdd.n10470 vdd.n10275 2.607
R50873 vdd.n10284 vdd.n10275 2.607
R50874 vdd.n10425 vdd.n10309 2.607
R50875 vdd.n10316 vdd.n10309 2.607
R50876 vdd.n13057 vdd.n9306 2.607
R50877 vdd.n13057 vdd.n13056 2.607
R50878 vdd.n9371 vdd.n9366 2.607
R50879 vdd.n9388 vdd.n9366 2.607
R50880 vdd.n9502 vdd.n9501 2.607
R50881 vdd.n9503 vdd.n9502 2.607
R50882 vdd.n12922 vdd.n12921 2.607
R50883 vdd.n12921 vdd.n9550 2.607
R50884 vdd.n12849 vdd.n9666 2.607
R50885 vdd.n12849 vdd.n12848 2.607
R50886 vdd.n9731 vdd.n9726 2.607
R50887 vdd.n9748 vdd.n9726 2.607
R50888 vdd.n9862 vdd.n9861 2.607
R50889 vdd.n9863 vdd.n9862 2.607
R50890 vdd.n12714 vdd.n12713 2.607
R50891 vdd.n12713 vdd.n9910 2.607
R50892 vdd.n12641 vdd.n10026 2.607
R50893 vdd.n12641 vdd.n12640 2.607
R50894 vdd.n10081 vdd.n10080 2.607
R50895 vdd.n10550 vdd.n10538 2.607
R50896 vdd.n12499 vdd.n10562 2.607
R50897 vdd.n10610 vdd.n10609 2.607
R50898 vdd.n12450 vdd.n10627 2.607
R50899 vdd.n12409 vdd.n10701 2.607
R50900 vdd.n10741 vdd.n10726 2.607
R50901 vdd.n10794 vdd.n10780 2.607
R50902 vdd.n12345 vdd.n10813 2.607
R50903 vdd.n10890 vdd.n10870 2.607
R50904 vdd.n10907 vdd.n10900 2.607
R50905 vdd.n10975 vdd.n10974 2.607
R50906 vdd.n12249 vdd.n12248 2.607
R50907 vdd.n12213 vdd.n12212 2.607
R50908 vdd.n12201 vdd.n12200 2.607
R50909 vdd.n12165 vdd.n11126 2.607
R50910 vdd.n11172 vdd.n11171 2.607
R50911 vdd.n12107 vdd.n11196 2.607
R50912 vdd.n11251 vdd.n11226 2.607
R50913 vdd.n11303 vdd.n11288 2.607
R50914 vdd.n12039 vdd.n11322 2.607
R50915 vdd.n11399 vdd.n11379 2.607
R50916 vdd.n11416 vdd.n11409 2.607
R50917 vdd.n11505 vdd.n11504 2.607
R50918 vdd.n11942 vdd.n11552 2.607
R50919 vdd.n15275 vdd.n15268 2.607
R50920 vdd.n15277 vdd.n15275 2.607
R50921 vdd.n15356 vdd.n15355 2.607
R50922 vdd.n15355 vdd.n15347 2.607
R50923 vdd.n15497 vdd.n15487 2.607
R50924 vdd.n15499 vdd.n15497 2.607
R50925 vdd.n15595 vdd.n15594 2.607
R50926 vdd.n15594 vdd.n15584 2.607
R50927 vdd.n15753 vdd.n15743 2.607
R50928 vdd.n15755 vdd.n15753 2.607
R50929 vdd.n15851 vdd.n15850 2.607
R50930 vdd.n15850 vdd.n15840 2.607
R50931 vdd.n16009 vdd.n15999 2.607
R50932 vdd.n16011 vdd.n16009 2.607
R50933 vdd.n16107 vdd.n16106 2.607
R50934 vdd.n16106 vdd.n16096 2.607
R50935 vdd.n16265 vdd.n16255 2.607
R50936 vdd.n16267 vdd.n16265 2.607
R50937 vdd.n16363 vdd.n16362 2.607
R50938 vdd.n16362 vdd.n16352 2.607
R50939 vdd.n16521 vdd.n16511 2.607
R50940 vdd.n16523 vdd.n16521 2.607
R50941 vdd.n16710 vdd.n16709 2.607
R50942 vdd.n16902 vdd.n16901 2.607
R50943 vdd.n16924 vdd.n16923 2.607
R50944 vdd.n17016 vdd.n17015 2.607
R50945 vdd.n17075 vdd.n17073 2.607
R50946 vdd.n17174 vdd.n17173 2.607
R50947 vdd.n17196 vdd.n17195 2.607
R50948 vdd.n17288 vdd.n17287 2.607
R50949 vdd.n17347 vdd.n17345 2.607
R50950 vdd.n17446 vdd.n17445 2.607
R50951 vdd.n17468 vdd.n17467 2.607
R50952 vdd.n17560 vdd.n17559 2.607
R50953 vdd.n17605 vdd.n17603 2.607
R50954 vdd.n17704 vdd.n17703 2.607
R50955 vdd.n17726 vdd.n17725 2.607
R50956 vdd.n17818 vdd.n17817 2.607
R50957 vdd.n17876 vdd.n17874 2.607
R50958 vdd.n17975 vdd.n17974 2.607
R50959 vdd.n17997 vdd.n17996 2.607
R50960 vdd.n18089 vdd.n18088 2.607
R50961 vdd.n18148 vdd.n18146 2.607
R50962 vdd.n18245 vdd.n18244 2.607
R50963 vdd.n18266 vdd.n18265 2.607
R50964 vdd.n18337 vdd.n18336 2.607
R50965 vdd.n18400 vdd.n18399 2.607
R50966 vdd.n2423 vdd.n2422 2.598
R50967 vdd.n10477 vdd.n10476 2.581
R50968 vdd.n10416 vdd.n10415 2.581
R50969 vdd.n15261 vdd.n15260 2.581
R50970 vdd.n11765 vdd.n11764 2.578
R50971 vdd.n21846 vdd.n21844 2.578
R50972 vdd.n13072 vdd.n13071 2.567
R50973 vdd.n9399 vdd.n9360 2.567
R50974 vdd.n9483 vdd.n9466 2.567
R50975 vdd.n12929 vdd.t308 2.567
R50976 vdd.n12906 vdd.n9562 2.567
R50977 vdd.n12864 vdd.n12863 2.567
R50978 vdd.n12852 vdd.t304 2.567
R50979 vdd.n9759 vdd.n9720 2.567
R50980 vdd.n12786 vdd.t301 2.567
R50981 vdd.n9843 vdd.n9826 2.567
R50982 vdd.n12698 vdd.n9920 2.567
R50983 vdd.n12656 vdd.n12655 2.567
R50984 vdd.n10105 vdd.n10062 2.567
R50985 vdd.n10512 vdd.t362 2.567
R50986 vdd.t371 vdd.n12535 2.567
R50987 vdd.n12513 vdd.n10528 2.567
R50988 vdd.n12459 vdd.n10615 2.567
R50989 vdd.n12401 vdd.n12400 2.567
R50990 vdd.n12364 vdd.n10774 2.567
R50991 vdd.n12307 vdd.n12306 2.567
R50992 vdd.n10985 vdd.n10984 2.567
R50993 vdd.n12152 vdd.n11137 2.567
R50994 vdd.n11234 vdd.n11221 2.567
R50995 vdd.n11307 vdd.t375 2.567
R50996 vdd.n12058 vdd.n11282 2.567
R50997 vdd.n12001 vdd.n12000 2.567
R50998 vdd.n11987 vdd.t364 2.567
R50999 vdd.n11528 vdd.n11527 2.567
R51000 vdd.n15474 vdd.n15473 2.567
R51001 vdd.n15608 vdd.n15607 2.567
R51002 vdd.n15730 vdd.n15729 2.567
R51003 vdd.n15828 vdd.t251 2.567
R51004 vdd.n15864 vdd.n15863 2.567
R51005 vdd.n15986 vdd.n15985 2.567
R51006 vdd.t261 vdd.n16003 2.567
R51007 vdd.n16120 vdd.n16119 2.567
R51008 vdd.t269 vdd.n15157 2.567
R51009 vdd.n16242 vdd.n16241 2.567
R51010 vdd.n16376 vdd.n16375 2.567
R51011 vdd.n16498 vdd.n16497 2.567
R51012 vdd.n16618 vdd.n16617 2.567
R51013 vdd.n16845 vdd.t6 2.567
R51014 vdd.n16849 vdd.t24 2.567
R51015 vdd.n16915 vdd.n16914 2.567
R51016 vdd.n17039 vdd.n17038 2.567
R51017 vdd.n17187 vdd.n17186 2.567
R51018 vdd.n17311 vdd.n17310 2.567
R51019 vdd.n17459 vdd.n17458 2.567
R51020 vdd.n17583 vdd.n17582 2.567
R51021 vdd.n17841 vdd.n17840 2.567
R51022 vdd.n17988 vdd.n17987 2.567
R51023 vdd.n18096 vdd.t12 2.567
R51024 vdd.n18112 vdd.n18111 2.567
R51025 vdd.n18257 vdd.n18256 2.567
R51026 vdd.n18287 vdd.t32 2.567
R51027 vdd.n18365 vdd.n18364 2.567
R51028 vdd.n15366 vdd.n15365 2.562
R51029 vdd.n1225 vdd.n1221 2.56
R51030 vdd.n9264 vdd.n9239 2.558
R51031 vdd.n9225 vdd.n9224 2.558
R51032 vdd.n2528 vdd.n2527 2.541
R51033 vdd.n1285 vdd.n1284 2.502
R51034 vdd.n31278 vdd.n31277 2.501
R51035 vdd.n31770 vdd.n31769 2.47
R51036 vdd.n25419 vdd.n25418 2.469
R51037 vdd.n35843 vdd.n35842 2.458
R51038 vdd.n36001 vdd.n36000 2.458
R51039 vdd.n36071 vdd.n36070 2.458
R51040 vdd.n36232 vdd.n36231 2.458
R51041 vdd.n36302 vdd.n36301 2.458
R51042 vdd.n36463 vdd.n36462 2.458
R51043 vdd.n36533 vdd.n36532 2.458
R51044 vdd.n36694 vdd.n36693 2.458
R51045 vdd.n36764 vdd.n36763 2.458
R51046 vdd.n36925 vdd.n36924 2.458
R51047 vdd.n3652 vdd.n3651 2.458
R51048 vdd.n33172 vdd.n33171 2.458
R51049 vdd.n33134 vdd.n33133 2.458
R51050 vdd.n2401 vdd.n2400 2.458
R51051 vdd.n37385 vdd.n37384 2.458
R51052 vdd.n32846 vdd.n32845 2.458
R51053 vdd.n38210 vdd.n38209 2.458
R51054 vdd.n38050 vdd.n38049 2.458
R51055 vdd.n37980 vdd.n37979 2.458
R51056 vdd.n37819 vdd.n37818 2.458
R51057 vdd.n37749 vdd.n37748 2.458
R51058 vdd.n28191 vdd.n28190 2.458
R51059 vdd.n28261 vdd.n28260 2.458
R51060 vdd.n28422 vdd.n28421 2.458
R51061 vdd.n28492 vdd.n28491 2.458
R51062 vdd.n28653 vdd.n28652 2.458
R51063 vdd.n28723 vdd.n28722 2.458
R51064 vdd.n26206 vdd.n26205 2.458
R51065 vdd.n31751 vdd.n31750 2.458
R51066 vdd.n27836 vdd.n27835 2.458
R51067 vdd.n27912 vdd.n27911 2.458
R51068 vdd.n31484 vdd.n31483 2.458
R51069 vdd.n30219 vdd.n30218 2.458
R51070 vdd.n30502 vdd.n30501 2.458
R51071 vdd.n13286 vdd.t106 2.446
R51072 vdd.n13304 vdd.n13303 2.446
R51073 vdd.t284 vdd.n13335 2.446
R51074 vdd.n13327 vdd.n9125 2.446
R51075 vdd.n13420 vdd.n9033 2.446
R51076 vdd.n13472 vdd.n9004 2.446
R51077 vdd.n13596 vdd.n13595 2.446
R51078 vdd.n13619 vdd.n8904 2.446
R51079 vdd.n8812 vdd.n8796 2.446
R51080 vdd.n13803 vdd.n8753 2.446
R51081 vdd.n13899 vdd.n8681 2.446
R51082 vdd.n13916 vdd.n13915 2.446
R51083 vdd.n14062 vdd.n8565 2.446
R51084 vdd.n14090 vdd.n8540 2.446
R51085 vdd.n14188 vdd.n8457 2.446
R51086 vdd.n14206 vdd.n14205 2.446
R51087 vdd.n14337 vdd.n8347 2.446
R51088 vdd.n14362 vdd.n14361 2.446
R51089 vdd.n14451 vdd.n8262 2.446
R51090 vdd.n14662 vdd.n8140 2.446
R51091 vdd.n31027 vdd.n31026 2.443
R51092 vdd.n11818 vdd.n11816 2.441
R51093 vdd.n21909 vdd.n21907 2.441
R51094 vdd.n25504 vdd.n25501 2.44
R51095 vdd.n11777 vdd.n11776 2.426
R51096 vdd.n21869 vdd.n21868 2.426
R51097 vdd.n12490 vdd.n10572 2.425
R51098 vdd.n12481 vdd.n10586 2.425
R51099 vdd.n12385 vdd.n10748 2.425
R51100 vdd.n12373 vdd.n10755 2.425
R51101 vdd.n10939 vdd.n10936 2.425
R51102 vdd.n12280 vdd.n10921 2.425
R51103 vdd.n11098 vdd.n11087 2.425
R51104 vdd.n11120 vdd.n11114 2.425
R51105 vdd.n12083 vdd.n11242 2.425
R51106 vdd.n12067 vdd.n11270 2.425
R51107 vdd.n11483 vdd.n11480 2.425
R51108 vdd.n11974 vdd.n11430 2.425
R51109 vdd.n10456 vdd.n10289 2.425
R51110 vdd.n10440 vdd.n10298 2.425
R51111 vdd.n9340 vdd.n9316 2.425
R51112 vdd.n13033 vdd.n9353 2.425
R51113 vdd.n12945 vdd.n9507 2.425
R51114 vdd.n9542 vdd.n9526 2.425
R51115 vdd.n9700 vdd.n9677 2.425
R51116 vdd.n12825 vdd.n9713 2.425
R51117 vdd.n12737 vdd.n9867 2.425
R51118 vdd.n9902 vdd.n9887 2.425
R51119 vdd.n10153 vdd.n10037 2.425
R51120 vdd.n12616 vdd.n10055 2.425
R51121 vdd.n16964 vdd.n16958 2.425
R51122 vdd.n16992 vdd.n16986 2.425
R51123 vdd.n17236 vdd.n17230 2.425
R51124 vdd.n17264 vdd.n17258 2.425
R51125 vdd.n17508 vdd.n17502 2.425
R51126 vdd.n17536 vdd.n17530 2.425
R51127 vdd.n17766 vdd.n17760 2.425
R51128 vdd.n17794 vdd.n17788 2.425
R51129 vdd.n18037 vdd.n18031 2.425
R51130 vdd.n18065 vdd.n18059 2.425
R51131 vdd.n18303 vdd.n18298 2.425
R51132 vdd.n15035 vdd.n15030 2.425
R51133 vdd.n15298 vdd.n15297 2.425
R51134 vdd.n15320 vdd.n15319 2.425
R51135 vdd.n15523 vdd.n15522 2.425
R51136 vdd.n15548 vdd.n15547 2.425
R51137 vdd.n15779 vdd.n15778 2.425
R51138 vdd.n15804 vdd.n15803 2.425
R51139 vdd.n16035 vdd.n16034 2.425
R51140 vdd.n16060 vdd.n16059 2.425
R51141 vdd.n16291 vdd.n16290 2.425
R51142 vdd.n16316 vdd.n16315 2.425
R51143 vdd.n16546 vdd.n16545 2.425
R51144 vdd.n16749 vdd.n16748 2.425
R51145 vdd.n1778 vdd.n1777 2.404
R51146 vdd.n2597 vdd.n2596 2.404
R51147 vdd.n2214 vdd.n2213 2.404
R51148 vdd.n1220 vdd.n1219 2.374
R51149 vdd.n10100 vdd.n10098 2.37
R51150 vdd.n10412 vdd.n10322 2.37
R51151 vdd.n10407 vdd.n10324 2.37
R51152 vdd.n13078 vdd.n13077 2.37
R51153 vdd.n9303 vdd.n9294 2.37
R51154 vdd.n13018 vdd.n13017 2.37
R51155 vdd.n13010 vdd.n9395 2.37
R51156 vdd.n9460 vdd.n9459 2.37
R51157 vdd.n9488 vdd.n9461 2.37
R51158 vdd.n9585 vdd.n9584 2.37
R51159 vdd.n9591 vdd.n9581 2.37
R51160 vdd.n12870 vdd.n12869 2.37
R51161 vdd.n9663 vdd.n9626 2.37
R51162 vdd.n12810 vdd.n12809 2.37
R51163 vdd.n12802 vdd.n9755 2.37
R51164 vdd.n9820 vdd.n9819 2.37
R51165 vdd.n9848 vdd.n9821 2.37
R51166 vdd.n9945 vdd.n9944 2.37
R51167 vdd.n9951 vdd.n9941 2.37
R51168 vdd.n12662 vdd.n12661 2.37
R51169 vdd.n10023 vdd.n9986 2.37
R51170 vdd.n10171 vdd.n10050 2.37
R51171 vdd.n10194 vdd.n10193 2.37
R51172 vdd.n10550 vdd.n10535 2.37
R51173 vdd.n12509 vdd.n10533 2.37
R51174 vdd.n10642 vdd.n10633 2.37
R51175 vdd.n10649 vdd.n10629 2.37
R51176 vdd.n10711 vdd.n10701 2.37
R51177 vdd.n10731 vdd.n10729 2.37
R51178 vdd.n12357 vdd.n10778 2.37
R51179 vdd.n12350 vdd.n10805 2.37
R51180 vdd.n12315 vdd.n10870 2.37
R51181 vdd.n12302 vdd.n12301 2.37
R51182 vdd.n10989 vdd.n10988 2.37
R51183 vdd.n12261 vdd.n12260 2.37
R51184 vdd.n12212 vdd.n11041 2.37
R51185 vdd.n11080 vdd.n11079 2.37
R51186 vdd.n11158 vdd.n11134 2.37
R51187 vdd.n11161 vdd.n11160 2.37
R51188 vdd.n12107 vdd.n11219 2.37
R51189 vdd.n12095 vdd.n12094 2.37
R51190 vdd.n12051 vdd.n11286 2.37
R51191 vdd.n12044 vdd.n11314 2.37
R51192 vdd.n12009 vdd.n11379 2.37
R51193 vdd.n11996 vdd.n11995 2.37
R51194 vdd.n11536 vdd.n11535 2.37
R51195 vdd.n11551 vdd.n11547 2.37
R51196 vdd.n16594 vdd.n16593 2.37
R51197 vdd.n15384 vdd.n15374 2.37
R51198 vdd.n15376 vdd.n15375 2.37
R51199 vdd.n15450 vdd.n15449 2.37
R51200 vdd.n15465 vdd.n15464 2.37
R51201 vdd.n15629 vdd.n15616 2.37
R51202 vdd.n15618 vdd.n15617 2.37
R51203 vdd.n15706 vdd.n15705 2.37
R51204 vdd.n15721 vdd.n15720 2.37
R51205 vdd.n15885 vdd.n15872 2.37
R51206 vdd.n15874 vdd.n15873 2.37
R51207 vdd.n15962 vdd.n15961 2.37
R51208 vdd.n15977 vdd.n15976 2.37
R51209 vdd.n16141 vdd.n16128 2.37
R51210 vdd.n16130 vdd.n16129 2.37
R51211 vdd.n16218 vdd.n16217 2.37
R51212 vdd.n16233 vdd.n16232 2.37
R51213 vdd.n16397 vdd.n16384 2.37
R51214 vdd.n16386 vdd.n16385 2.37
R51215 vdd.n16474 vdd.n16473 2.37
R51216 vdd.n16489 vdd.n16488 2.37
R51217 vdd.n16761 vdd.n16758 2.37
R51218 vdd.n16729 vdd.n16728 2.37
R51219 vdd.n16901 vdd.n16892 2.37
R51220 vdd.n16934 vdd.n16922 2.37
R51221 vdd.n17043 vdd.n17042 2.37
R51222 vdd.n17057 vdd.n17048 2.37
R51223 vdd.n17173 vdd.n17164 2.37
R51224 vdd.n17206 vdd.n17194 2.37
R51225 vdd.n17315 vdd.n17314 2.37
R51226 vdd.n17329 vdd.n17320 2.37
R51227 vdd.n17445 vdd.n17436 2.37
R51228 vdd.n17478 vdd.n17466 2.37
R51229 vdd.n17587 vdd.n17586 2.37
R51230 vdd.n17594 vdd.n16831 2.37
R51231 vdd.n17703 vdd.n17694 2.37
R51232 vdd.n17736 vdd.n17724 2.37
R51233 vdd.n17845 vdd.n17844 2.37
R51234 vdd.n17859 vdd.n17850 2.37
R51235 vdd.n17974 vdd.n17965 2.37
R51236 vdd.n18007 vdd.n17995 2.37
R51237 vdd.n18116 vdd.n18115 2.37
R51238 vdd.n18130 vdd.n18121 2.37
R51239 vdd.n18244 vdd.n18236 2.37
R51240 vdd.n18275 vdd.n18264 2.37
R51241 vdd.n18395 vdd.n18394 2.37
R51242 vdd.n22140 vdd.n22139 2.36
R51243 vdd.n22338 vdd.n22337 2.36
R51244 vdd.n28052 vdd.n28051 2.346
R51245 vdd.n29745 vdd.n29744 2.346
R51246 vdd.n19279 vdd.n19278 2.345
R51247 vdd.n19243 vdd.n19242 2.345
R51248 vdd.n19223 vdd.n19222 2.345
R51249 vdd.n19186 vdd.n19185 2.345
R51250 vdd.n19840 vdd.n19839 2.345
R51251 vdd.n19877 vdd.n19876 2.345
R51252 vdd.n19909 vdd.n19908 2.345
R51253 vdd.n19945 vdd.n19944 2.345
R51254 vdd.n20419 vdd.n20416 2.345
R51255 vdd.n20361 vdd.n20360 2.345
R51256 vdd.n20183 vdd.n20180 2.345
R51257 vdd.n20125 vdd.n20124 2.345
R51258 vdd.n11758 vdd.n11681 2.342
R51259 vdd.n11877 vdd.n11803 2.34
R51260 vdd.n21968 vdd.n21894 2.34
R51261 vdd.n3636 vdd.n3635 2.339
R51262 vdd.n1274 vdd.n1273 2.339
R51263 vdd.n14695 vdd.n8124 2.339
R51264 vdd.n14741 vdd.n8105 2.339
R51265 vdd.n14869 vdd.n8034 2.339
R51266 vdd.n14895 vdd.n14894 2.339
R51267 vdd.n30342 vdd.n30341 2.339
R51268 vdd.n11752 vdd.n11751 2.335
R51269 vdd.n29777 vdd.n29776 2.33
R51270 vdd.n24531 vdd.n24525 2.327
R51271 vdd.n11916 vdd.n11908 2.326
R51272 vdd.n22002 vdd.n21998 2.326
R51273 vdd.n24533 vdd.n24532 2.325
R51274 vdd.n31480 vdd.n31479 2.319
R51275 vdd.n31637 vdd.n31636 2.319
R51276 vdd.n26201 vdd.n26200 2.319
R51277 vdd.n11779 vdd.n11777 2.316
R51278 vdd.n4020 vdd.n1928 2.307
R51279 vdd.n24558 vdd.n24557 2.296
R51280 vdd.n24942 vdd.n24911 2.296
R51281 vdd.n4020 vdd.n1958 2.293
R51282 vdd.n28892 vdd.n28891 2.287
R51283 vdd.n28053 vdd.n28052 2.284
R51284 vdd.n27889 vdd.n27888 2.284
R51285 vdd.n29746 vdd.n29745 2.284
R51286 vdd.n30681 vdd.n30680 2.284
R51287 vdd.n11869 vdd.n11808 2.283
R51288 vdd.n21960 vdd.n21899 2.283
R51289 vdd.n11896 vdd.n11895 2.282
R51290 vdd.n21987 vdd.n21986 2.282
R51291 vdd.n11764 vdd.n11763 2.281
R51292 vdd.n21844 vdd.n21843 2.281
R51293 vdd.n11766 vdd.n11765 2.278
R51294 vdd.n21846 vdd.n21845 2.278
R51295 vdd.n11901 vdd.n11791 2.273
R51296 vdd.n11753 vdd.n11682 2.273
R51297 vdd.n21992 vdd.n21882 2.273
R51298 vdd.n11776 vdd.n11664 2.27
R51299 vdd.n11872 vdd.n11871 2.27
R51300 vdd.n21963 vdd.n21962 2.27
R51301 vdd.n11757 vdd.n11682 2.262
R51302 vdd.n21837 vdd.n21798 2.262
R51303 vdd.n33724 vdd.n33723 2.258
R51304 vdd.n33398 vdd.n33397 2.258
R51305 vdd.n34120 vdd.n34119 2.258
R51306 vdd.n34320 vdd.n34319 2.258
R51307 vdd.n33990 vdd.n33989 2.258
R51308 vdd.n35152 vdd.n35151 2.258
R51309 vdd.n35586 vdd.n35585 2.258
R51310 vdd.n35507 vdd.n35506 2.258
R51311 vdd.n34974 vdd.n34973 2.258
R51312 vdd.n34892 vdd.n34891 2.258
R51313 vdd.n34567 vdd.n34566 2.258
R51314 vdd.n888 vdd.n887 2.258
R51315 vdd.n717 vdd.n716 2.258
R51316 vdd.n376 vdd.n375 2.258
R51317 vdd.n169 vdd.n168 2.258
R51318 vdd.n45 vdd.n44 2.258
R51319 vdd.n448 vdd.n447 2.258
R51320 vdd.n6278 vdd.n6277 2.258
R51321 vdd.n5935 vdd.n5934 2.258
R51322 vdd.n5987 vdd.n5986 2.258
R51323 vdd.n5721 vdd.n5720 2.258
R51324 vdd.n5639 vdd.n5638 2.258
R51325 vdd.n5314 vdd.n5313 2.258
R51326 vdd.n4626 vdd.n4625 2.258
R51327 vdd.n5147 vdd.n5146 2.258
R51328 vdd.n4887 vdd.n4886 2.258
R51329 vdd.n4886 vdd.n4885 2.258
R51330 vdd.n4551 vdd.n4550 2.258
R51331 vdd.n4466 vdd.n4465 2.258
R51332 vdd.n4145 vdd.n4144 2.258
R51333 vdd.n30246 vdd.n30245 2.258
R51334 vdd.n31449 vdd.n31448 2.258
R51335 vdd.n32131 vdd.n32130 2.258
R51336 vdd.n31147 vdd.n31143 2.258
R51337 vdd.n30505 vdd.n30344 2.258
R51338 vdd.n35846 vdd.n35708 2.258
R51339 vdd.n36004 vdd.n35997 2.258
R51340 vdd.n36074 vdd.n36067 2.258
R51341 vdd.n36235 vdd.n36228 2.258
R51342 vdd.n36305 vdd.n36298 2.258
R51343 vdd.n36466 vdd.n36459 2.258
R51344 vdd.n36536 vdd.n36529 2.258
R51345 vdd.n36697 vdd.n36690 2.258
R51346 vdd.n36767 vdd.n36760 2.258
R51347 vdd.n36928 vdd.n36921 2.258
R51348 vdd.n37006 vdd.n37002 2.258
R51349 vdd.n33175 vdd.n33168 2.258
R51350 vdd.n33137 vdd.n33130 2.258
R51351 vdd.n37313 vdd.n37309 2.258
R51352 vdd.n37388 vdd.n37381 2.258
R51353 vdd.n32849 vdd.n32842 2.258
R51354 vdd.n38213 vdd.n38206 2.258
R51355 vdd.n38053 vdd.n38046 2.258
R51356 vdd.n37983 vdd.n37976 2.258
R51357 vdd.n37822 vdd.n37815 2.258
R51358 vdd.n37752 vdd.n37745 2.258
R51359 vdd.n28194 vdd.n28187 2.258
R51360 vdd.n28264 vdd.n28257 2.258
R51361 vdd.n28425 vdd.n28418 2.258
R51362 vdd.n28495 vdd.n28488 2.258
R51363 vdd.n28656 vdd.n28649 2.258
R51364 vdd.n28726 vdd.n28719 2.258
R51365 vdd.n28181 vdd.n28180 2.258
R51366 vdd.n28123 vdd.n28122 2.258
R51367 vdd.n28066 vdd.n28057 2.258
R51368 vdd.n28070 vdd.n28069 2.258
R51369 vdd.n27839 vdd.n27832 2.258
R51370 vdd.n27915 vdd.n27908 2.258
R51371 vdd.n30198 vdd.n30197 2.258
R51372 vdd.n27396 vdd.n27395 2.258
R51373 vdd.n27452 vdd.n27451 2.258
R51374 vdd.n27617 vdd.n27616 2.258
R51375 vdd.n25842 vdd.n25841 2.258
R51376 vdd.n25898 vdd.n25897 2.258
R51377 vdd.n26038 vdd.n26037 2.258
R51378 vdd.n26394 vdd.n26393 2.258
R51379 vdd.n31747 vdd.n31746 2.258
R51380 vdd.n27212 vdd.n27211 2.258
R51381 vdd.n1681 vdd.n1677 2.258
R51382 vdd.n1627 vdd.n1623 2.258
R51383 vdd.n1500 vdd.n1496 2.258
R51384 vdd.n1446 vdd.n1442 2.258
R51385 vdd.n1319 vdd.n1315 2.258
R51386 vdd.n26785 vdd.n26781 2.258
R51387 vdd.n26912 vdd.n26908 2.258
R51388 vdd.n26966 vdd.n26962 2.258
R51389 vdd.n27093 vdd.n27089 2.258
R51390 vdd.n27147 vdd.n27143 2.258
R51391 vdd.n2668 vdd.n2667 2.258
R51392 vdd.n2672 vdd.n2671 2.258
R51393 vdd.n2183 vdd.n2182 2.258
R51394 vdd.n3759 vdd.n3758 2.258
R51395 vdd.n3744 vdd.n3743 2.258
R51396 vdd.n3728 vdd.n3727 2.258
R51397 vdd.n2703 vdd.n2702 2.258
R51398 vdd.n2741 vdd.n2737 2.258
R51399 vdd.n2865 vdd.n2861 2.258
R51400 vdd.n2919 vdd.n2915 2.258
R51401 vdd.n3046 vdd.n3042 2.258
R51402 vdd.n3100 vdd.n3096 2.258
R51403 vdd.n3227 vdd.n3223 2.258
R51404 vdd.n3281 vdd.n3277 2.258
R51405 vdd.n3408 vdd.n3404 2.258
R51406 vdd.n3462 vdd.n3458 2.258
R51407 vdd.n3589 vdd.n3585 2.258
R51408 vdd.n3655 vdd.n3648 2.258
R51409 vdd.n31779 vdd.n31777 2.258
R51410 vdd.n31722 vdd.n31721 2.258
R51411 vdd.n31932 vdd.n31931 2.258
R51412 vdd.n13121 vdd.n13120 2.258
R51413 vdd.n13122 vdd.n13121 2.258
R51414 vdd.n13340 vdd.n9097 2.258
R51415 vdd.n13346 vdd.n9097 2.258
R51416 vdd.n13413 vdd.n13412 2.258
R51417 vdd.n13414 vdd.n13413 2.258
R51418 vdd.n13632 vdd.n8877 2.258
R51419 vdd.n13638 vdd.n8877 2.258
R51420 vdd.n13707 vdd.n13706 2.258
R51421 vdd.n13708 vdd.n13707 2.258
R51422 vdd.n13908 vdd.n8674 2.258
R51423 vdd.n13908 vdd.n8675 2.258
R51424 vdd.n13989 vdd.n13988 2.258
R51425 vdd.n13988 vdd.n8606 2.258
R51426 vdd.n14198 vdd.n8450 2.258
R51427 vdd.n14198 vdd.n8451 2.258
R51428 vdd.n14280 vdd.n14279 2.258
R51429 vdd.n14279 vdd.n8384 2.258
R51430 vdd.n14496 vdd.n8218 2.258
R51431 vdd.n14498 vdd.n14496 2.258
R51432 vdd.n14670 vdd.n8131 2.258
R51433 vdd.n14678 vdd.n14677 2.258
R51434 vdd.n14737 vdd.n8109 2.258
R51435 vdd.n14727 vdd.n14722 2.258
R51436 vdd.n14842 vdd.n8041 2.258
R51437 vdd.n14850 vdd.n14849 2.258
R51438 vdd.n14891 vdd.n14890 2.258
R51439 vdd.n14916 vdd.n8014 2.258
R51440 vdd.n13141 vdd.n9249 2.258
R51441 vdd.n9228 vdd.n9194 2.258
R51442 vdd.n13227 vdd.n9194 2.258
R51443 vdd.n13314 vdd.n13313 2.258
R51444 vdd.n13313 vdd.n9135 2.258
R51445 vdd.n13466 vdd.n8972 2.258
R51446 vdd.n13519 vdd.n8972 2.258
R51447 vdd.n13606 vdd.n13605 2.258
R51448 vdd.n13605 vdd.n8913 2.258
R51449 vdd.n13795 vdd.n8758 2.258
R51450 vdd.n13795 vdd.n8763 2.258
R51451 vdd.n13886 vdd.n8697 2.258
R51452 vdd.n13886 vdd.n8699 2.258
R51453 vdd.n14082 vdd.n8545 2.258
R51454 vdd.n14082 vdd.n8550 2.258
R51455 vdd.n14175 vdd.n8474 2.258
R51456 vdd.n14175 vdd.n8476 2.258
R51457 vdd.n8329 vdd.n8310 2.258
R51458 vdd.n14383 vdd.n8310 2.258
R51459 vdd.n14471 vdd.n14470 2.258
R51460 vdd.n14472 vdd.n14471 2.258
R51461 vdd.n10405 vdd.n10320 2.258
R51462 vdd.n24224 vdd.n24223 2.258
R51463 vdd.n24233 vdd.n24232 2.258
R51464 vdd.n24124 vdd.n24123 2.258
R51465 vdd.n24042 vdd.n24041 2.258
R51466 vdd.n23892 vdd.n23891 2.258
R51467 vdd.n23810 vdd.n23809 2.258
R51468 vdd.n23660 vdd.n23659 2.258
R51469 vdd.n23122 vdd.n23121 2.258
R51470 vdd.n23204 vdd.n23203 2.258
R51471 vdd.n23354 vdd.n23353 2.258
R51472 vdd.n23436 vdd.n23435 2.258
R51473 vdd.n23586 vdd.n23585 2.258
R51474 vdd.n22543 vdd.n22542 2.258
R51475 vdd.n22625 vdd.n22624 2.258
R51476 vdd.n22775 vdd.n22774 2.258
R51477 vdd.n22857 vdd.n22856 2.258
R51478 vdd.n23007 vdd.n23006 2.258
R51479 vdd.n22396 vdd.n22395 2.258
R51480 vdd.n22405 vdd.n22404 2.258
R51481 vdd.n22212 vdd.n22204 2.258
R51482 vdd.n22211 vdd.n22206 2.258
R51483 vdd.n24341 vdd.n24340 2.258
R51484 vdd.n24350 vdd.n24349 2.258
R51485 vdd.n22076 vdd.n22068 2.258
R51486 vdd.n22075 vdd.n22070 2.258
R51487 vdd.n19337 vdd.n19301 2.258
R51488 vdd.n19513 vdd.n19504 2.258
R51489 vdd.n19543 vdd.n19534 2.258
R51490 vdd.n19714 vdd.n19705 2.258
R51491 vdd.n19745 vdd.n19736 2.258
R51492 vdd.n20942 vdd.n20933 2.258
R51493 vdd.n20911 vdd.n20902 2.258
R51494 vdd.n20752 vdd.n20743 2.258
R51495 vdd.n20722 vdd.n20713 2.258
R51496 vdd.n20546 vdd.n19971 2.258
R51497 vdd.n21681 vdd.n21680 2.258
R51498 vdd.n21562 vdd.n21553 2.258
R51499 vdd.n21480 vdd.n21471 2.258
R51500 vdd.n21303 vdd.n21294 2.258
R51501 vdd.n21221 vdd.n21212 2.258
R51502 vdd.n21044 vdd.n21035 2.258
R51503 vdd.n19114 vdd.n19105 2.258
R51504 vdd.n18937 vdd.n18928 2.258
R51505 vdd.n18855 vdd.n18846 2.258
R51506 vdd.n18678 vdd.n18669 2.258
R51507 vdd.n18596 vdd.n18587 2.258
R51508 vdd.n20429 vdd.n20428 2.258
R51509 vdd.n20339 vdd.n20338 2.258
R51510 vdd.n20193 vdd.n20192 2.258
R51511 vdd.n20103 vdd.n20102 2.258
R51512 vdd.n24711 vdd.n24710 2.258
R51513 vdd.n24776 vdd.n24775 2.258
R51514 vdd.n25194 vdd.n25193 2.258
R51515 vdd.n25129 vdd.n25128 2.258
R51516 vdd.n11770 vdd.n11668 2.257
R51517 vdd.n21858 vdd.n21757 2.257
R51518 vdd.n11870 vdd.n11869 2.251
R51519 vdd.n21961 vdd.n21960 2.251
R51520 vdd.n2676 vdd.n2675 2.251
R51521 vdd.n4020 vdd.n4019 2.25
R51522 vdd.n26080 vdd.n26079 2.25
R51523 vdd.n27658 vdd.n27657 2.25
R51524 vdd.n38216 vdd.n35644 2.25
R51525 vdd.n38216 vdd.n35654 2.25
R51526 vdd.n38216 vdd.n35673 2.25
R51527 vdd.n38216 vdd.n37042 2.25
R51528 vdd.n38216 vdd.n33285 2.25
R51529 vdd.n38216 vdd.n37062 2.25
R51530 vdd.n38216 vdd.n33272 2.25
R51531 vdd.n38216 vdd.n37076 2.25
R51532 vdd.n38216 vdd.n33252 2.25
R51533 vdd.n38216 vdd.n37099 2.25
R51534 vdd.n38216 vdd.n33225 2.25
R51535 vdd.n38216 vdd.n37119 2.25
R51536 vdd.n38216 vdd.n33203 2.25
R51537 vdd.n38216 vdd.n37132 2.25
R51538 vdd.n38216 vdd.n33185 2.25
R51539 vdd.n38216 vdd.n37153 2.25
R51540 vdd.n38216 vdd.n33162 2.25
R51541 vdd.n38216 vdd.n37169 2.25
R51542 vdd.n38216 vdd.n37188 2.25
R51543 vdd.n38216 vdd.n33139 2.25
R51544 vdd.n38216 vdd.n37208 2.25
R51545 vdd.n38216 vdd.n33116 2.25
R51546 vdd.n38216 vdd.n37221 2.25
R51547 vdd.n38216 vdd.n33099 2.25
R51548 vdd.n38216 vdd.n37239 2.25
R51549 vdd.n38216 vdd.n33088 2.25
R51550 vdd.n38216 vdd.n37262 2.25
R51551 vdd.n38216 vdd.n33064 2.25
R51552 vdd.n38216 vdd.n37285 2.25
R51553 vdd.n38216 vdd.n33041 2.25
R51554 vdd.n38216 vdd.n37296 2.25
R51555 vdd.n38216 vdd.n33023 2.25
R51556 vdd.n38216 vdd.n37315 2.25
R51557 vdd.n38216 vdd.n33004 2.25
R51558 vdd.n38216 vdd.n37340 2.25
R51559 vdd.n38216 vdd.n37364 2.25
R51560 vdd.n38216 vdd.n32982 2.25
R51561 vdd.n38216 vdd.n37390 2.25
R51562 vdd.n38216 vdd.n32963 2.25
R51563 vdd.n38216 vdd.n37411 2.25
R51564 vdd.n38216 vdd.n32944 2.25
R51565 vdd.n38216 vdd.n37433 2.25
R51566 vdd.n38216 vdd.n32937 2.25
R51567 vdd.n38216 vdd.n37457 2.25
R51568 vdd.n38216 vdd.n32919 2.25
R51569 vdd.n38216 vdd.n37473 2.25
R51570 vdd.n38216 vdd.n32894 2.25
R51571 vdd.n38216 vdd.n37497 2.25
R51572 vdd.n38216 vdd.n32878 2.25
R51573 vdd.n38216 vdd.n37516 2.25
R51574 vdd.n38216 vdd.n32859 2.25
R51575 vdd.n38216 vdd.n37538 2.25
R51576 vdd.n38216 vdd.n37551 2.25
R51577 vdd.n38216 vdd.n32836 2.25
R51578 vdd.n38216 vdd.n37574 2.25
R51579 vdd.n38216 vdd.n38215 2.25
R51580 vdd.n27243 vdd.n27242 2.25
R51581 vdd.n26157 vdd.n26156 2.25
R51582 vdd.n26180 vdd.n26179 2.25
R51583 vdd.n26215 vdd.n26214 2.25
R51584 vdd.n26622 vdd.n26621 2.25
R51585 vdd.n26708 vdd.n26707 2.25
R51586 vdd.n26670 vdd.n26669 2.25
R51587 vdd.n26319 vdd.n26318 2.25
R51588 vdd.n26351 vdd.n26350 2.25
R51589 vdd.n26404 vdd.n26403 2.25
R51590 vdd.n26519 vdd.n26518 2.25
R51591 vdd.n11608 vdd.n11607 2.25
R51592 vdd.n11620 vdd.n11583 2.25
R51593 vdd.n9252 vdd.n9250 2.25
R51594 vdd.n10221 vdd.n10075 2.25
R51595 vdd.n11761 vdd.n11760 2.25
R51596 vdd.n11749 vdd.n11748 2.25
R51597 vdd.n11773 vdd.n11665 2.25
R51598 vdd.n11671 vdd.n11669 2.25
R51599 vdd.n11875 vdd.n11874 2.25
R51600 vdd.n11880 vdd.n11801 2.25
R51601 vdd.n11797 vdd.n11796 2.25
R51602 vdd.n11899 vdd.n11898 2.25
R51603 vdd.n11904 vdd.n11788 2.25
R51604 vdd.n11785 vdd.n11662 2.25
R51605 vdd.n21840 vdd.n21763 2.25
R51606 vdd.n21856 vdd.n21855 2.25
R51607 vdd.n21966 vdd.n21965 2.25
R51608 vdd.n21971 vdd.n21892 2.25
R51609 vdd.n21888 vdd.n21887 2.25
R51610 vdd.n21990 vdd.n21989 2.25
R51611 vdd.n21995 vdd.n21879 2.25
R51612 vdd.n21878 vdd.n21877 2.25
R51613 vdd.n24531 vdd.n24530 2.25
R51614 vdd.n4020 vdd.n2100 2.248
R51615 vdd.n4020 vdd.n2006 2.248
R51616 vdd.n4020 vdd.n2562 2.248
R51617 vdd.n13074 vdd.n9290 2.246
R51618 vdd.n13014 vdd.n13013 2.246
R51619 vdd.n12963 vdd.n9465 2.246
R51620 vdd.n9579 vdd.n9564 2.246
R51621 vdd.n12866 vdd.n9622 2.246
R51622 vdd.n12806 vdd.n12805 2.246
R51623 vdd.n12755 vdd.n9825 2.246
R51624 vdd.n9939 vdd.n9938 2.246
R51625 vdd.n12658 vdd.n9982 2.246
R51626 vdd.n10107 vdd.n10104 2.246
R51627 vdd.n10554 vdd.n10553 2.246
R51628 vdd.n10646 vdd.n10645 2.246
R51629 vdd.n10713 vdd.n10708 2.246
R51630 vdd.n12354 vdd.n12353 2.246
R51631 vdd.n12317 vdd.n10867 2.246
R51632 vdd.n12263 vdd.n10959 2.246
R51633 vdd.n12209 vdd.n11046 2.246
R51634 vdd.n12151 vdd.n12150 2.246
R51635 vdd.n12104 vdd.n12103 2.246
R51636 vdd.n12048 vdd.n12047 2.246
R51637 vdd.n12011 vdd.n11376 2.246
R51638 vdd.n11957 vdd.n11444 2.246
R51639 vdd.n11660 vdd.n11659 2.246
R51640 vdd.n15461 vdd.n15457 2.246
R51641 vdd.n15626 vdd.n15625 2.246
R51642 vdd.n15717 vdd.n15713 2.246
R51643 vdd.n15882 vdd.n15881 2.246
R51644 vdd.n15973 vdd.n15969 2.246
R51645 vdd.n16138 vdd.n16137 2.246
R51646 vdd.n16229 vdd.n16225 2.246
R51647 vdd.n16394 vdd.n16393 2.246
R51648 vdd.n16485 vdd.n16481 2.246
R51649 vdd.n16625 vdd.n16624 2.246
R51650 vdd.n16898 vdd.n16895 2.246
R51651 vdd.n17054 vdd.n17051 2.246
R51652 vdd.n17170 vdd.n17167 2.246
R51653 vdd.n17326 vdd.n17323 2.246
R51654 vdd.n17442 vdd.n17439 2.246
R51655 vdd.n16827 vdd.n16824 2.246
R51656 vdd.n17700 vdd.n17697 2.246
R51657 vdd.n17856 vdd.n17853 2.246
R51658 vdd.n17971 vdd.n17968 2.246
R51659 vdd.n18127 vdd.n18124 2.246
R51660 vdd.n18241 vdd.n18239 2.246
R51661 vdd.n15022 vdd.n15021 2.246
R51662 vdd.n21741 vdd.n21709 2.246
R51663 vdd.n10205 vdd.n10091 2.245
R51664 vdd.n10198 vdd.n10079 2.245
R51665 vdd.n24973 vdd.n24953 2.244
R51666 vdd.n11494 vdd.n11466 2.244
R51667 vdd.n11488 vdd.n11469 2.244
R51668 vdd.n18314 vdd.n15038 2.244
R51669 vdd.n18310 vdd.n16818 2.244
R51670 vdd.n11786 vdd.n11663 2.242
R51671 vdd.n21755 vdd.n21752 2.242
R51672 vdd.n15381 vdd.n15380 2.242
R51673 vdd.n10179 vdd.n10082 2.242
R51674 vdd.n11755 vdd.n11754 2.242
R51675 vdd.n11783 vdd.n11782 2.239
R51676 vdd.n21875 vdd.n21874 2.239
R51677 vdd.n13117 vdd.t319 2.239
R51678 vdd.n13198 vdd.n9212 2.239
R51679 vdd.n13188 vdd.n9222 2.239
R51680 vdd.n11919 vdd.n11918 2.237
R51681 vdd.n35869 vdd.n35868 2.235
R51682 vdd.n35974 vdd.n35973 2.235
R51683 vdd.n36100 vdd.n36099 2.235
R51684 vdd.n36205 vdd.n36204 2.235
R51685 vdd.n36331 vdd.n36330 2.235
R51686 vdd.n36436 vdd.n36435 2.235
R51687 vdd.n36562 vdd.n36561 2.235
R51688 vdd.n36667 vdd.n36666 2.235
R51689 vdd.n36793 vdd.n36792 2.235
R51690 vdd.n36898 vdd.n36897 2.235
R51691 vdd.n2054 vdd.n2053 2.235
R51692 vdd.n2012 vdd.n2011 2.235
R51693 vdd.n2194 vdd.n2193 2.235
R51694 vdd.n2038 vdd.n2037 2.235
R51695 vdd.n37407 vdd.n37406 2.235
R51696 vdd.n1195 vdd.n1194 2.235
R51697 vdd.n1282 vdd.n1281 2.235
R51698 vdd.n38079 vdd.n38078 2.235
R51699 vdd.n37953 vdd.n37952 2.235
R51700 vdd.n37848 vdd.n37847 2.235
R51701 vdd.n37722 vdd.n37721 2.235
R51702 vdd.n37617 vdd.n37616 2.235
R51703 vdd.n28290 vdd.n28289 2.235
R51704 vdd.n28395 vdd.n28394 2.235
R51705 vdd.n28521 vdd.n28520 2.235
R51706 vdd.n28626 vdd.n28625 2.235
R51707 vdd.n28752 vdd.n28751 2.235
R51708 vdd.n28138 vdd.n28137 2.235
R51709 vdd.n28966 vdd.n28965 2.235
R51710 vdd.n27809 vdd.n27808 2.235
R51711 vdd.n32156 vdd.n32155 2.235
R51712 vdd.n31512 vdd.n31508 2.235
R51713 vdd.n32447 vdd.n32443 2.235
R51714 vdd.n31275 vdd.n31274 2.235
R51715 vdd.n1201 vdd.n1197 2.221
R51716 vdd.n2655 vdd.n2651 2.221
R51717 vdd.n2180 vdd.n2179 2.221
R51718 vdd.n2723 vdd.n2722 2.221
R51719 vdd.n29017 vdd.n27769 2.22
R51720 vdd.n3656 vdd.n3655 2.156
R51721 vdd.n35847 vdd.n35846 2.155
R51722 vdd.n30506 vdd.n30505 2.155
R51723 vdd.n2742 vdd.n2741 2.155
R51724 vdd.n31148 vdd.n31147 2.155
R51725 vdd.n13303 vdd.n9142 2.141
R51726 vdd.n13328 vdd.n13327 2.141
R51727 vdd.n13492 vdd.n8992 2.141
R51728 vdd.n13482 vdd.n9002 2.141
R51729 vdd.n13529 vdd.t126 2.141
R51730 vdd.n13595 vdd.n8921 2.141
R51731 vdd.n13608 vdd.t136 2.141
R51732 vdd.n13620 vdd.n13619 2.141
R51733 vdd.n13772 vdd.n8776 2.141
R51734 vdd.n13762 vdd.n8785 2.141
R51735 vdd.n13778 vdd.t104 2.141
R51736 vdd.t104 vdd.n8765 2.141
R51737 vdd.n13809 vdd.t285 2.141
R51738 vdd.n13840 vdd.t112 2.141
R51739 vdd.t330 vdd.n13870 2.141
R51740 vdd.n13899 vdd.n8682 2.141
R51741 vdd.n13917 vdd.n13916 2.141
R51742 vdd.n14052 vdd.n14051 2.141
R51743 vdd.n8576 vdd.n8560 2.141
R51744 vdd.t290 vdd.n14068 2.141
R51745 vdd.n14125 vdd.t329 2.141
R51746 vdd.n14188 vdd.n8458 2.141
R51747 vdd.n14207 vdd.n14206 2.141
R51748 vdd.n14327 vdd.n14326 2.141
R51749 vdd.n14325 vdd.t102 2.141
R51750 vdd.n14372 vdd.n8318 2.141
R51751 vdd.n8262 vdd.n8261 2.141
R51752 vdd.n14480 vdd.n8197 2.141
R51753 vdd.n11625 vdd.n11580 2.133
R51754 vdd.n21646 vdd.n21636 2.133
R51755 vdd.n32059 vdd.n32058 2.133
R51756 vdd.n32069 vdd.n32059 2.133
R51757 vdd.n2522 vdd.n2521 2.133
R51758 vdd.n2416 vdd.n2415 2.133
R51759 vdd.n10420 vdd.n10419 2.133
R51760 vdd.n10419 vdd.n10312 2.133
R51761 vdd.n13069 vdd.n13068 2.133
R51762 vdd.n13068 vdd.n9301 2.133
R51763 vdd.n13021 vdd.n9363 2.133
R51764 vdd.n13021 vdd.n9364 2.133
R51765 vdd.n9494 vdd.n9485 2.133
R51766 vdd.n9494 vdd.n9486 2.133
R51767 vdd.n12910 vdd.n9558 2.133
R51768 vdd.n12910 vdd.n12909 2.133
R51769 vdd.n12861 vdd.n12860 2.133
R51770 vdd.n12860 vdd.n9661 2.133
R51771 vdd.n12813 vdd.n9723 2.133
R51772 vdd.n12813 vdd.n9724 2.133
R51773 vdd.n9854 vdd.n9845 2.133
R51774 vdd.n9854 vdd.n9846 2.133
R51775 vdd.n12702 vdd.n9917 2.133
R51776 vdd.n12702 vdd.n12701 2.133
R51777 vdd.n12653 vdd.n12652 2.133
R51778 vdd.n12652 vdd.n10021 2.133
R51779 vdd.n10170 vdd.n10169 2.133
R51780 vdd.n12623 vdd.n10051 2.133
R51781 vdd.n10558 vdd.n10532 2.133
R51782 vdd.n12511 vdd.n12510 2.133
R51783 vdd.n10637 vdd.n10636 2.133
R51784 vdd.n10650 vdd.n10649 2.133
R51785 vdd.n12404 vdd.n12403 2.133
R51786 vdd.n10730 vdd.n10704 2.133
R51787 vdd.n12362 vdd.n10777 2.133
R51788 vdd.n12350 vdd.n12349 2.133
R51789 vdd.n12309 vdd.n10871 2.133
R51790 vdd.n12303 vdd.n10894 2.133
R51791 vdd.n10981 vdd.n10966 2.133
R51792 vdd.n12260 vdd.n10964 2.133
R51793 vdd.n11072 vdd.n11066 2.133
R51794 vdd.n11078 vdd.n11063 2.133
R51795 vdd.n11133 vdd.n11132 2.133
R51796 vdd.n11161 vdd.n11156 2.133
R51797 vdd.n12099 vdd.n11223 2.133
R51798 vdd.n11232 vdd.n11225 2.133
R51799 vdd.n12056 vdd.n11285 2.133
R51800 vdd.n12044 vdd.n12043 2.133
R51801 vdd.n12003 vdd.n11380 2.133
R51802 vdd.n11997 vdd.n11403 2.133
R51803 vdd.n11530 vdd.n11457 2.133
R51804 vdd.n15370 vdd.n15369 2.133
R51805 vdd.n15369 vdd.n15362 2.133
R51806 vdd.n15480 vdd.n15470 2.133
R51807 vdd.n15482 vdd.n15480 2.133
R51808 vdd.n15612 vdd.n15611 2.133
R51809 vdd.n15611 vdd.n15601 2.133
R51810 vdd.n15736 vdd.n15726 2.133
R51811 vdd.n15738 vdd.n15736 2.133
R51812 vdd.n15868 vdd.n15867 2.133
R51813 vdd.n15867 vdd.n15857 2.133
R51814 vdd.n15992 vdd.n15982 2.133
R51815 vdd.n15994 vdd.n15992 2.133
R51816 vdd.n16124 vdd.n16123 2.133
R51817 vdd.n16123 vdd.n16113 2.133
R51818 vdd.n16248 vdd.n16238 2.133
R51819 vdd.n16250 vdd.n16248 2.133
R51820 vdd.n16380 vdd.n16379 2.133
R51821 vdd.n16379 vdd.n16369 2.133
R51822 vdd.n16504 vdd.n16494 2.133
R51823 vdd.n16506 vdd.n16504 2.133
R51824 vdd.n16767 vdd.n16766 2.133
R51825 vdd.n16745 vdd.n16744 2.133
R51826 vdd.n16918 vdd.n16917 2.133
R51827 vdd.n16908 vdd.n16907 2.133
R51828 vdd.n17032 vdd.n17031 2.133
R51829 vdd.n17059 vdd.n17057 2.133
R51830 vdd.n17190 vdd.n17189 2.133
R51831 vdd.n17180 vdd.n17179 2.133
R51832 vdd.n17304 vdd.n17303 2.133
R51833 vdd.n17331 vdd.n17329 2.133
R51834 vdd.n17462 vdd.n17461 2.133
R51835 vdd.n17452 vdd.n17451 2.133
R51836 vdd.n17576 vdd.n17575 2.133
R51837 vdd.n17594 vdd.n17593 2.133
R51838 vdd.n17720 vdd.n17719 2.133
R51839 vdd.n17710 vdd.n17709 2.133
R51840 vdd.n17834 vdd.n17833 2.133
R51841 vdd.n17861 vdd.n17859 2.133
R51842 vdd.n17991 vdd.n17990 2.133
R51843 vdd.n17981 vdd.n17980 2.133
R51844 vdd.n18105 vdd.n18104 2.133
R51845 vdd.n18132 vdd.n18130 2.133
R51846 vdd.n18260 vdd.n18259 2.133
R51847 vdd.n18251 vdd.n18250 2.133
R51848 vdd.n18360 vdd.n18359 2.133
R51849 vdd.n27783 vdd.n27782 2.129
R51850 vdd.n28178 vdd.n28156 2.113
R51851 vdd.n38139 vdd.n38126 2.113
R51852 vdd.n25513 vdd.n25512 2.113
R51853 vdd.n1748 vdd.n1740 2.113
R51854 vdd.n1748 vdd.n1747 2.113
R51855 vdd.n26755 vdd.n26748 2.113
R51856 vdd.n38139 vdd.n38137 2.113
R51857 vdd.n4020 vdd.n2061 2.111
R51858 vdd.n21610 vdd.n21609 2.111
R51859 vdd.n21516 vdd.t275 2.111
R51860 vdd.n21413 vdd.n21410 2.111
R51861 vdd.n21364 vdd.n21361 2.111
R51862 vdd.n21154 vdd.n21151 2.111
R51863 vdd.n21105 vdd.n21102 2.111
R51864 vdd.n19047 vdd.n19044 2.111
R51865 vdd.n18998 vdd.n18995 2.111
R51866 vdd.n18788 vdd.n18785 2.111
R51867 vdd.n18739 vdd.n18736 2.111
R51868 vdd.n18632 vdd.t352 2.111
R51869 vdd.n18529 vdd.n18526 2.111
R51870 vdd.n4020 vdd.n1188 2.104
R51871 vdd.n4020 vdd.n2020 2.104
R51872 vdd.n4020 vdd.n2032 2.104
R51873 vdd.n31167 vdd.n31131 2.102
R51874 vdd.n31175 vdd.n31169 2.102
R51875 vdd.n30592 vdd.n30285 2.096
R51876 vdd.n28178 vdd.n28166 2.093
R51877 vdd.n26755 vdd.n26738 2.093
R51878 vdd.n2508 vdd.n2507 2.086
R51879 vdd.n31167 vdd.n31164 2.085
R51880 vdd.n31175 vdd.n31171 2.085
R51881 vdd.n3657 vdd.n3646 2.085
R51882 vdd.n28178 vdd.n28176 2.079
R51883 vdd.n31279 vdd.n31261 2.079
R51884 vdd.n4020 vdd.n2046 2.077
R51885 vdd.n30507 vdd.n30506 2.075
R51886 vdd.n35848 vdd.n35847 2.075
R51887 vdd.n2743 vdd.n2742 2.075
R51888 vdd.n31149 vdd.n31148 2.075
R51889 vdd.n3657 vdd.n3656 2.075
R51890 vdd.n1286 vdd.n1285 2.072
R51891 vdd.n31279 vdd.n31278 2.072
R51892 vdd.n31171 vdd.n31170 2.071
R51893 vdd.n31164 vdd.n31163 2.071
R51894 vdd.n30507 vdd.n30342 2.07
R51895 vdd.n1286 vdd.n1274 2.07
R51896 vdd.n3657 vdd.n3636 2.07
R51897 vdd.n2135 vdd.n2134 2.067
R51898 vdd.n4020 vdd.n1181 2.064
R51899 vdd.n4020 vdd.n2025 2.064
R51900 vdd.n4020 vdd.n2047 2.064
R51901 vdd.n30582 vdd.n30302 2.053
R51902 vdd.n11546 vdd.n11545 2.014
R51903 vdd.n35854 vdd.n35853 2.011
R51904 vdd.n35987 vdd.n35986 2.011
R51905 vdd.n36085 vdd.n36084 2.011
R51906 vdd.n36218 vdd.n36217 2.011
R51907 vdd.n36316 vdd.n36315 2.011
R51908 vdd.n36449 vdd.n36448 2.011
R51909 vdd.n36547 vdd.n36546 2.011
R51910 vdd.n36680 vdd.n36679 2.011
R51911 vdd.n36778 vdd.n36777 2.011
R51912 vdd.n36911 vdd.n36910 2.011
R51913 vdd.n3632 vdd.n3631 2.011
R51914 vdd.n33194 vdd.n33193 2.011
R51915 vdd.n37203 vdd.n37202 2.011
R51916 vdd.n2377 vdd.n2376 2.011
R51917 vdd.n32958 vdd.n32957 2.011
R51918 vdd.n1905 vdd.n1904 2.011
R51919 vdd.n1270 vdd.n1269 2.011
R51920 vdd.n38064 vdd.n38063 2.011
R51921 vdd.n37966 vdd.n37965 2.011
R51922 vdd.n37833 vdd.n37832 2.011
R51923 vdd.n37735 vdd.n37734 2.011
R51924 vdd.n37602 vdd.n37601 2.011
R51925 vdd.n28275 vdd.n28274 2.011
R51926 vdd.n28408 vdd.n28407 2.011
R51927 vdd.n28506 vdd.n28505 2.011
R51928 vdd.n28639 vdd.n28638 2.011
R51929 vdd.n28737 vdd.n28736 2.011
R51930 vdd.n28810 vdd.n28809 2.011
R51931 vdd.n28062 vdd.n28061 2.011
R51932 vdd.n31654 vdd.n31653 2.011
R51933 vdd.n32121 vdd.n32120 2.011
R51934 vdd.n29762 vdd.n29761 2.011
R51935 vdd.n30234 vdd.n30233 2.011
R51936 vdd.n30338 vdd.n30337 2.011
R51937 vdd.n27841 vdd.n27840 2.002
R51938 vdd.n35908 vdd.n35907 1.965
R51939 vdd.n35928 vdd.n35927 1.965
R51940 vdd.n36139 vdd.n36138 1.965
R51941 vdd.n36159 vdd.n36158 1.965
R51942 vdd.n36370 vdd.n36369 1.965
R51943 vdd.n36390 vdd.n36389 1.965
R51944 vdd.n36601 vdd.n36600 1.965
R51945 vdd.n36621 vdd.n36620 1.965
R51946 vdd.n36832 vdd.n36831 1.965
R51947 vdd.n36852 vdd.n36851 1.965
R51948 vdd.n33263 vdd.n33262 1.965
R51949 vdd.n33244 vdd.n33243 1.965
R51950 vdd.n33069 vdd.n33068 1.965
R51951 vdd.n37254 vdd.n37253 1.965
R51952 vdd.n37440 vdd.n37439 1.965
R51953 vdd.n32909 vdd.n32908 1.965
R51954 vdd.n38120 vdd.n38119 1.965
R51955 vdd.n38130 vdd.n38129 1.965
R51956 vdd.n37907 vdd.n37906 1.965
R51957 vdd.n37887 vdd.n37886 1.965
R51958 vdd.n37676 vdd.n37675 1.965
R51959 vdd.n37656 vdd.n37655 1.965
R51960 vdd.n28329 vdd.n28328 1.965
R51961 vdd.n28349 vdd.n28348 1.965
R51962 vdd.n28560 vdd.n28559 1.965
R51963 vdd.n28580 vdd.n28579 1.965
R51964 vdd.n28791 vdd.n28790 1.965
R51965 vdd.n28147 vdd.n28146 1.965
R51966 vdd.n27762 vdd.n27761 1.965
R51967 vdd.n31889 vdd.n31888 1.965
R51968 vdd.n32227 vdd.n32226 1.965
R51969 vdd.n29688 vdd.n29687 1.965
R51970 vdd.n30294 vdd.n30293 1.965
R51971 vdd.n30563 vdd.n30562 1.965
R51972 vdd.n2791 vdd.n2790 1.965
R51973 vdd.n2808 vdd.n2807 1.965
R51974 vdd.n2972 vdd.n2971 1.965
R51975 vdd.n2989 vdd.n2988 1.965
R51976 vdd.n3153 vdd.n3152 1.965
R51977 vdd.n3170 vdd.n3169 1.965
R51978 vdd.n3334 vdd.n3333 1.965
R51979 vdd.n3351 vdd.n3350 1.965
R51980 vdd.n3515 vdd.n3514 1.965
R51981 vdd.n3532 vdd.n3531 1.965
R51982 vdd.n3708 vdd.n3707 1.965
R51983 vdd.n4009 vdd.n4008 1.965
R51984 vdd.n2281 vdd.n2280 1.965
R51985 vdd.n2300 vdd.n2299 1.965
R51986 vdd.n1977 vdd.n1976 1.965
R51987 vdd.n1987 vdd.n1986 1.965
R51988 vdd.n1737 vdd.n1736 1.965
R51989 vdd.n1744 vdd.n1743 1.965
R51990 vdd.n1570 vdd.n1569 1.965
R51991 vdd.n1553 vdd.n1552 1.965
R51992 vdd.n1389 vdd.n1388 1.965
R51993 vdd.n1372 vdd.n1371 1.965
R51994 vdd.n26838 vdd.n26837 1.965
R51995 vdd.n26855 vdd.n26854 1.965
R51996 vdd.n27019 vdd.n27018 1.965
R51997 vdd.n27036 vdd.n27035 1.965
R51998 vdd.n27200 vdd.n27199 1.965
R51999 vdd.n26743 vdd.n26742 1.965
R52000 vdd.n31865 vdd.n31864 1.965
R52001 vdd.n31885 vdd.n31884 1.965
R52002 vdd.n32223 vdd.n32222 1.965
R52003 vdd.n32256 vdd.n32255 1.965
R52004 vdd.n31117 vdd.n31116 1.965
R52005 vdd.n31177 vdd.n31176 1.965
R52006 vdd.n13215 vdd.n9203 1.965
R52007 vdd.n13247 vdd.n9177 1.965
R52008 vdd.n13508 vdd.n8982 1.965
R52009 vdd.n13539 vdd.n8956 1.965
R52010 vdd.n13790 vdd.n8768 1.965
R52011 vdd.n13824 vdd.n8737 1.965
R52012 vdd.n14117 vdd.n8513 1.965
R52013 vdd.n14128 vdd.n8506 1.965
R52014 vdd.n14397 vdd.n8302 1.965
R52015 vdd.n14429 vdd.n8276 1.965
R52016 vdd.n14786 vdd.n8071 1.965
R52017 vdd.n8079 vdd.n8065 1.965
R52018 vdd.n11627 vdd.n11575 1.965
R52019 vdd.n13144 vdd.n9247 1.965
R52020 vdd.n13380 vdd.n13379 1.965
R52021 vdd.n13437 vdd.n9023 1.965
R52022 vdd.n13672 vdd.n13671 1.965
R52023 vdd.n13729 vdd.n8803 1.965
R52024 vdd.n13951 vdd.n8633 1.965
R52025 vdd.n13994 vdd.n8587 1.965
R52026 vdd.n14241 vdd.n8411 1.965
R52027 vdd.n14285 vdd.n8367 1.965
R52028 vdd.n14540 vdd.n8180 1.965
R52029 vdd.n14613 vdd.n8168 1.965
R52030 vdd.n19410 vdd.n19409 1.965
R52031 vdd.n19427 vdd.n19426 1.965
R52032 vdd.n19613 vdd.n19612 1.965
R52033 vdd.n19630 vdd.n19629 1.965
R52034 vdd.n19815 vdd.n19814 1.965
R52035 vdd.n19165 vdd.n19164 1.965
R52036 vdd.n20835 vdd.n20834 1.965
R52037 vdd.n20821 vdd.n20820 1.965
R52038 vdd.n20633 vdd.n20632 1.965
R52039 vdd.n20619 vdd.n20618 1.965
R52040 vdd.n21662 vdd.n21661 1.965
R52041 vdd.n21657 vdd.n21656 1.965
R52042 vdd.n21390 vdd.n21389 1.965
R52043 vdd.n21376 vdd.n21375 1.965
R52044 vdd.n21131 vdd.n21130 1.965
R52045 vdd.n21117 vdd.n21116 1.965
R52046 vdd.n19024 vdd.n19023 1.965
R52047 vdd.n19010 vdd.n19009 1.965
R52048 vdd.n18765 vdd.n18764 1.965
R52049 vdd.n18751 vdd.n18750 1.965
R52050 vdd.n18506 vdd.n18505 1.965
R52051 vdd.n18465 vdd.n18464 1.965
R52052 vdd.n19999 vdd.n19993 1.965
R52053 vdd.n20011 vdd.n20005 1.965
R52054 vdd.n24982 vdd.n24981 1.965
R52055 vdd.n3646 vdd.n3645 1.95
R52056 vdd.n24739 vdd.n24738 1.945
R52057 vdd.n25171 vdd.n25170 1.945
R52058 vdd.n25170 vdd.n25169 1.945
R52059 vdd.n24738 vdd.n24737 1.945
R52060 vdd.n1173 vdd.n802 1.94
R52061 vdd.n1173 vdd.n948 1.94
R52062 vdd.n1173 vdd.n882 1.939
R52063 vdd.n1173 vdd.n866 1.938
R52064 vdd.n1173 vdd.n854 1.938
R52065 vdd.n1173 vdd.n913 1.938
R52066 vdd.n1173 vdd.n795 1.936
R52067 vdd.n10277 vdd.n10276 1.936
R52068 vdd.n10319 vdd.n10318 1.936
R52069 vdd.n15272 vdd.n15271 1.936
R52070 vdd.n1173 vdd.n951 1.934
R52071 vdd.n1173 vdd.n812 1.933
R52072 vdd.n587 vdd.n212 1.933
R52073 vdd.n1173 vdd.n842 1.93
R52074 vdd.n33724 vdd.n33722 1.925
R52075 vdd.n888 vdd.n886 1.925
R52076 vdd.n13061 vdd.n13060 1.925
R52077 vdd.n9386 vdd.n9359 1.925
R52078 vdd.n9499 vdd.n9498 1.925
R52079 vdd.n12918 vdd.n12917 1.925
R52080 vdd.n9614 ldomc_0.otaldom_0.pmosrm_0.vdd 1.925
R52081 vdd.n12853 vdd.n12852 1.925
R52082 vdd.n9746 vdd.n9719 1.925
R52083 vdd.n9859 vdd.n9858 1.925
R52084 vdd.n12710 vdd.n12709 1.925
R52085 vdd.n12645 vdd.n12644 1.925
R52086 vdd.n10191 vdd.n10061 1.925
R52087 vdd.n12543 vdd.t359 1.925
R52088 vdd.n12503 vdd.n12502 1.925
R52089 vdd.n12502 vdd.t311 1.925
R52090 vdd.n12461 vdd.n10614 1.925
R52091 vdd.n10738 vdd.n10737 1.925
R52092 vdd.n10798 vdd.n10797 1.925
R52093 vdd.n10909 vdd.n10896 1.925
R52094 vdd.n12269 vdd.n10952 1.925
R52095 vdd.t377 vdd.n11074 1.925
R52096 vdd.n12203 vdd.n11056 1.925
R52097 vdd.n12162 vdd.n12161 1.925
R52098 vdd.n12091 vdd.n12090 1.925
R52099 vdd.n11307 vdd.n11306 1.925
R52100 vdd.n11418 vdd.n11405 1.925
R52101 vdd.n11963 vdd.n11437 1.925
R52102 vdd.n15491 vdd.n15490 1.925
R52103 vdd.n15591 vdd.n15590 1.925
R52104 vdd.n15747 vdd.n15746 1.925
R52105 vdd.n15847 vdd.n15846 1.925
R52106 bandgapmd_0.otam_1.pmosrm_0.vdd vdd.n15196 1.925
R52107 vdd.n16003 vdd.n16002 1.925
R52108 vdd.n16103 vdd.n16102 1.925
R52109 vdd.n16259 vdd.n16258 1.925
R52110 vdd.n16359 vdd.n16358 1.925
R52111 vdd.n16515 vdd.n16514 1.925
R52112 vdd.n16612 vdd.n16611 1.925
R52113 vdd.t22 vdd.n16841 1.925
R52114 vdd.n16931 vdd.n16930 1.925
R52115 vdd.n16930 vdd.t252 1.925
R52116 vdd.n17023 vdd.n17022 1.925
R52117 vdd.n17203 vdd.n17202 1.925
R52118 vdd.n17295 vdd.n17294 1.925
R52119 vdd.n17475 vdd.n17474 1.925
R52120 vdd.n17567 vdd.n17566 1.925
R52121 vdd.n17717 vdd.t10 1.925
R52122 vdd.n17733 vdd.n17732 1.925
R52123 vdd.n17825 vdd.n17824 1.925
R52124 vdd.n18004 vdd.n18003 1.925
R52125 vdd.n18096 vdd.n18095 1.925
R52126 vdd.n18272 vdd.n18271 1.925
R52127 vdd.n18344 vdd.n18343 1.925
R52128 vdd.n15352 vdd.n15351 1.921
R52129 vdd.n13118 vdd.n13117 1.919
R52130 vdd.n13229 vdd.n9190 1.919
R52131 vdd.n33735 vdd.n33733 1.91
R52132 vdd.n936 vdd.n934 1.91
R52133 vdd.n13218 vdd.t323 1.897
R52134 vdd.n10097 vdd.n10096 1.896
R52135 vdd.n12603 vdd.n12602 1.896
R52136 vdd.n10090 vdd.n10065 1.896
R52137 vdd.n10421 vdd.n10420 1.896
R52138 vdd.n10413 vdd.n10312 1.896
R52139 vdd.n13069 vdd.n9300 1.896
R52140 vdd.n13064 vdd.n9301 1.896
R52141 vdd.n9390 vdd.n9363 1.896
R52142 vdd.n9394 vdd.n9364 1.896
R52143 vdd.n9487 vdd.n9485 1.896
R52144 vdd.n9490 vdd.n9486 1.896
R52145 vdd.n12914 vdd.n9558 1.896
R52146 vdd.n12909 vdd.n9560 1.896
R52147 vdd.n12861 vdd.n9660 1.896
R52148 vdd.n12856 vdd.n9661 1.896
R52149 vdd.n9750 vdd.n9723 1.896
R52150 vdd.n9754 vdd.n9724 1.896
R52151 vdd.n9847 vdd.n9845 1.896
R52152 vdd.n9850 vdd.n9846 1.896
R52153 vdd.n12706 vdd.n9917 1.896
R52154 vdd.n12701 vdd.n9919 1.896
R52155 vdd.n12653 vdd.n10020 1.896
R52156 vdd.n12648 vdd.n10021 1.896
R52157 vdd.n10558 vdd.n10557 1.896
R52158 vdd.n12511 vdd.n10532 1.896
R52159 vdd.n10638 vdd.n10637 1.896
R52160 vdd.n10651 vdd.n10650 1.896
R52161 vdd.n12405 vdd.n12404 1.896
R52162 vdd.n12403 vdd.n10704 1.896
R52163 vdd.n12362 vdd.n12361 1.896
R52164 vdd.n12349 vdd.n10809 1.896
R52165 vdd.n12313 vdd.n10871 1.896
R52166 vdd.n12309 vdd.n10894 1.896
R52167 vdd.n10987 vdd.n10966 1.896
R52168 vdd.n12256 vdd.n10964 1.896
R52169 vdd.n11068 vdd.n11066 1.896
R52170 vdd.n11072 vdd.n11063 1.896
R52171 vdd.n12154 vdd.n11133 1.896
R52172 vdd.n11165 vdd.n11156 1.896
R52173 vdd.n12100 vdd.n12099 1.896
R52174 vdd.n11232 vdd.n11223 1.896
R52175 vdd.n12056 vdd.n12055 1.896
R52176 vdd.n12043 vdd.n11318 1.896
R52177 vdd.n12007 vdd.n11380 1.896
R52178 vdd.n12003 vdd.n11403 1.896
R52179 vdd.n11518 vdd.n11459 1.896
R52180 vdd.n11949 vdd.n11546 1.896
R52181 vdd.n16688 vdd.n16687 1.896
R52182 vdd.n16700 vdd.n16697 1.896
R52183 vdd.n16701 vdd.n16696 1.896
R52184 vdd.n15370 vdd.n15360 1.896
R52185 vdd.n15362 vdd.n15361 1.896
R52186 vdd.n15470 vdd.n15469 1.896
R52187 vdd.n15482 vdd.n15481 1.896
R52188 vdd.n15612 vdd.n15599 1.896
R52189 vdd.n15601 vdd.n15600 1.896
R52190 vdd.n15726 vdd.n15725 1.896
R52191 vdd.n15738 vdd.n15737 1.896
R52192 vdd.n15868 vdd.n15855 1.896
R52193 vdd.n15857 vdd.n15856 1.896
R52194 vdd.n15982 vdd.n15981 1.896
R52195 vdd.n15994 vdd.n15993 1.896
R52196 vdd.n16124 vdd.n16111 1.896
R52197 vdd.n16113 vdd.n16112 1.896
R52198 vdd.n16238 vdd.n16237 1.896
R52199 vdd.n16250 vdd.n16249 1.896
R52200 vdd.n16380 vdd.n16367 1.896
R52201 vdd.n16369 vdd.n16368 1.896
R52202 vdd.n16494 vdd.n16493 1.896
R52203 vdd.n16506 vdd.n16505 1.896
R52204 vdd.n16918 vdd.n16906 1.896
R52205 vdd.n16917 vdd.n16908 1.896
R52206 vdd.n17041 vdd.n17032 1.896
R52207 vdd.n17059 vdd.n17058 1.896
R52208 vdd.n17190 vdd.n17178 1.896
R52209 vdd.n17189 vdd.n17180 1.896
R52210 vdd.n17313 vdd.n17304 1.896
R52211 vdd.n17331 vdd.n17330 1.896
R52212 vdd.n17462 vdd.n17450 1.896
R52213 vdd.n17461 vdd.n17452 1.896
R52214 vdd.n17585 vdd.n17576 1.896
R52215 vdd.n17593 vdd.n16832 1.896
R52216 vdd.n17720 vdd.n17708 1.896
R52217 vdd.n17719 vdd.n17710 1.896
R52218 vdd.n17843 vdd.n17834 1.896
R52219 vdd.n17861 vdd.n17860 1.896
R52220 vdd.n17991 vdd.n17979 1.896
R52221 vdd.n17990 vdd.n17981 1.896
R52222 vdd.n18114 vdd.n18105 1.896
R52223 vdd.n18132 vdd.n18131 1.896
R52224 vdd.n18260 vdd.n18249 1.896
R52225 vdd.n18259 vdd.n18251 1.896
R52226 vdd.n18387 vdd.n18385 1.896
R52227 vdd.n33786 vdd.n33785 1.882
R52228 vdd.n33714 vdd.n33713 1.882
R52229 vdd.n33683 vdd.n33682 1.882
R52230 vdd.n33346 vdd.n33345 1.882
R52231 vdd.n34218 vdd.n34217 1.882
R52232 vdd.n34087 vdd.n34086 1.882
R52233 vdd.n34321 vdd.n34320 1.882
R52234 vdd.n33909 vdd.n33908 1.882
R52235 vdd.n35078 vdd.n35077 1.882
R52236 vdd.n35587 vdd.n35586 1.882
R52237 vdd.n35248 vdd.n35247 1.882
R52238 vdd.n35338 vdd.n35337 1.882
R52239 vdd.n34754 vdd.n34753 1.882
R52240 vdd.n34661 vdd.n34660 1.882
R52241 vdd.n34893 vdd.n34892 1.882
R52242 vdd.n34491 vdd.n34490 1.882
R52243 vdd.n862 vdd.n861 1.882
R52244 vdd.n904 vdd.n903 1.882
R52245 vdd.n1148 vdd.n1147 1.882
R52246 vdd.n612 vdd.n611 1.882
R52247 vdd.n231 vdd.n230 1.882
R52248 vdd.n242 vdd.n241 1.882
R52249 vdd.n517 vdd.n516 1.882
R52250 vdd.n6183 vdd.n6182 1.882
R52251 vdd.n5936 vdd.n5935 1.882
R52252 vdd.n5789 vdd.n5788 1.882
R52253 vdd.n5919 vdd.n5918 1.882
R52254 vdd.n5501 vdd.n5500 1.882
R52255 vdd.n5408 vdd.n5407 1.882
R52256 vdd.n5640 vdd.n5639 1.882
R52257 vdd.n5238 vdd.n5237 1.882
R52258 vdd.n4627 vdd.n4626 1.882
R52259 vdd.n4988 vdd.n4987 1.882
R52260 vdd.n4813 vdd.n4812 1.882
R52261 vdd.n4328 vdd.n4327 1.882
R52262 vdd.n4238 vdd.n4237 1.882
R52263 vdd.n4467 vdd.n4466 1.882
R52264 vdd.n4068 vdd.n4067 1.882
R52265 vdd.n30253 vdd.n30251 1.882
R52266 vdd.n30267 vdd.n30266 1.882
R52267 vdd.n30276 vdd.n30275 1.882
R52268 vdd.n31526 vdd.n31525 1.882
R52269 vdd.n32182 vdd.n32181 1.882
R52270 vdd.n32179 vdd.n32178 1.882
R52271 vdd.n31065 vdd.n31064 1.882
R52272 vdd.n31068 vdd.n31067 1.882
R52273 vdd.n31253 vdd.n31252 1.882
R52274 vdd.n30526 vdd.n30525 1.882
R52275 vdd.n35878 vdd.n35877 1.882
R52276 vdd.n35955 vdd.n35954 1.882
R52277 vdd.n36109 vdd.n36108 1.882
R52278 vdd.n36186 vdd.n36185 1.882
R52279 vdd.n36340 vdd.n36339 1.882
R52280 vdd.n36417 vdd.n36416 1.882
R52281 vdd.n36571 vdd.n36570 1.882
R52282 vdd.n36648 vdd.n36647 1.882
R52283 vdd.n36802 vdd.n36801 1.882
R52284 vdd.n36879 vdd.n36878 1.882
R52285 vdd.n33279 vdd.n33278 1.882
R52286 vdd.n33213 vdd.n33212 1.882
R52287 vdd.n37215 vdd.n37214 1.882
R52288 vdd.n37272 vdd.n37271 1.882
R52289 vdd.n37413 vdd.n37412 1.882
R52290 vdd.n37475 vdd.n37474 1.882
R52291 vdd.n38161 vdd.n38160 1.882
R52292 vdd.n38088 vdd.n38087 1.882
R52293 vdd.n37934 vdd.n37933 1.882
R52294 vdd.n37857 vdd.n37856 1.882
R52295 vdd.n37703 vdd.n37702 1.882
R52296 vdd.n37626 vdd.n37625 1.882
R52297 vdd.n28299 vdd.n28298 1.882
R52298 vdd.n28376 vdd.n28375 1.882
R52299 vdd.n28530 vdd.n28529 1.882
R52300 vdd.n28607 vdd.n28606 1.882
R52301 vdd.n28761 vdd.n28760 1.882
R52302 vdd.n28168 vdd.n28167 1.882
R52303 vdd.n28816 vdd.n28813 1.882
R52304 vdd.n28983 vdd.n28982 1.882
R52305 vdd.n28980 vdd.n28979 1.882
R52306 vdd.n27787 vdd.n27786 1.882
R52307 vdd.n27801 vdd.n27800 1.882
R52308 vdd.n29889 vdd.n29888 1.882
R52309 vdd.n29881 vdd.n29879 1.882
R52310 vdd.n29856 vdd.n29855 1.882
R52311 vdd.n29827 vdd.n29826 1.882
R52312 vdd.n29821 vdd.n29820 1.882
R52313 vdd.n29766 vdd.n29756 1.882
R52314 vdd.n27350 vdd.n27349 1.882
R52315 vdd.n27294 vdd.n27293 1.882
R52316 vdd.n27453 vdd.n27452 1.882
R52317 vdd.n27543 vdd.n27542 1.882
R52318 vdd.n25802 vdd.n25801 1.882
R52319 vdd.n25746 vdd.n25745 1.882
R52320 vdd.n25899 vdd.n25898 1.882
R52321 vdd.n25980 vdd.n25979 1.882
R52322 vdd.n25504 vdd.n25503 1.882
R52323 vdd.n26750 vdd.n26749 1.882
R52324 vdd.n27213 vdd.n27212 1.882
R52325 vdd.n1765 vdd.n1764 1.882
R52326 vdd.n1710 vdd.n1709 1.882
R52327 vdd.n1590 vdd.n1589 1.882
R52328 vdd.n1529 vdd.n1528 1.882
R52329 vdd.n1409 vdd.n1408 1.882
R52330 vdd.n1348 vdd.n1347 1.882
R52331 vdd.n26814 vdd.n26813 1.882
R52332 vdd.n26875 vdd.n26874 1.882
R52333 vdd.n26995 vdd.n26994 1.882
R52334 vdd.n27056 vdd.n27055 1.882
R52335 vdd.n27176 vdd.n27175 1.882
R52336 vdd.n1234 vdd.n1233 1.882
R52337 vdd.n1901 vdd.n1900 1.882
R52338 vdd.n1200 vdd.n1199 1.882
R52339 vdd.n1910 vdd.n1909 1.882
R52340 vdd.n1931 vdd.n1930 1.882
R52341 vdd.n1203 vdd.n1190 1.882
R52342 vdd.n1933 vdd.n1929 1.882
R52343 vdd.n2650 vdd.n2649 1.882
R52344 vdd.n2404 vdd.n2397 1.882
R52345 vdd.n2406 vdd.n2394 1.882
R52346 vdd.n2028 vdd.n2027 1.882
R52347 vdd.n2030 vdd.n2026 1.882
R52348 vdd.n2182 vdd.n2181 1.882
R52349 vdd.n2172 vdd.n2171 1.882
R52350 vdd.n3828 vdd.n3826 1.882
R52351 vdd.n3818 vdd.n3817 1.882
R52352 vdd.n3757 vdd.n3756 1.882
R52353 vdd.n3755 vdd.n3754 1.882
R52354 vdd.n3744 vdd.n3740 1.882
R52355 vdd.n2690 vdd.n2689 1.882
R52356 vdd.n2703 vdd.n2700 1.882
R52357 vdd.n2726 vdd.n2723 1.882
R52358 vdd.n2725 vdd.n2724 1.882
R52359 vdd.n2715 vdd.n2714 1.882
R52360 vdd.n2767 vdd.n2766 1.882
R52361 vdd.n2828 vdd.n2827 1.882
R52362 vdd.n2948 vdd.n2947 1.882
R52363 vdd.n3009 vdd.n3008 1.882
R52364 vdd.n3129 vdd.n3128 1.882
R52365 vdd.n3190 vdd.n3189 1.882
R52366 vdd.n3310 vdd.n3309 1.882
R52367 vdd.n3371 vdd.n3370 1.882
R52368 vdd.n3491 vdd.n3490 1.882
R52369 vdd.n3552 vdd.n3551 1.882
R52370 vdd.n31712 vdd.n31711 1.882
R52371 vdd.n31715 vdd.n31714 1.882
R52372 vdd.n31928 vdd.n31927 1.882
R52373 vdd.n13190 vdd.n9220 1.882
R52374 vdd.n13183 vdd.n13180 1.882
R52375 vdd.n13270 vdd.n9161 1.882
R52376 vdd.n13289 vdd.n9148 1.882
R52377 vdd.n13484 vdd.n9000 1.882
R52378 vdd.n13477 vdd.n13475 1.882
R52379 vdd.n13562 vdd.n8939 1.882
R52380 vdd.n13581 vdd.n8927 1.882
R52381 vdd.n13764 vdd.n8783 1.882
R52382 vdd.n13757 vdd.n13755 1.882
R52383 vdd.n13844 vdd.n8723 1.882
R52384 vdd.n13849 vdd.n8724 1.882
R52385 vdd.n14041 vdd.n14040 1.882
R52386 vdd.n14073 vdd.n8557 1.882
R52387 vdd.n14133 vdd.n8502 1.882
R52388 vdd.n14138 vdd.n8503 1.882
R52389 vdd.n14347 vdd.n8340 1.882
R52390 vdd.n14349 vdd.n8336 1.882
R52391 vdd.n8281 vdd.n8244 1.882
R52392 vdd.n8248 vdd.n8245 1.882
R52393 vdd.n14654 vdd.n14653 1.882
R52394 vdd.n14653 vdd.n8150 1.882
R52395 vdd.n14764 vdd.n8086 1.882
R52396 vdd.n14771 vdd.n8086 1.882
R52397 vdd.n14826 vdd.n14825 1.882
R52398 vdd.n14825 vdd.n8059 1.882
R52399 vdd.n14939 vdd.n14938 1.882
R52400 vdd.n14940 vdd.n14939 1.882
R52401 vdd.n9259 vdd.n9256 1.882
R52402 vdd.n13159 vdd.n9235 1.882
R52403 vdd.n13363 vdd.n13362 1.882
R52404 vdd.n9078 vdd.n9075 1.882
R52405 vdd.n9028 vdd.n9014 1.882
R52406 vdd.n13453 vdd.n9011 1.882
R52407 vdd.n13655 vdd.n13654 1.882
R52408 vdd.n8858 vdd.n8855 1.882
R52409 vdd.n8808 vdd.n8794 1.882
R52410 vdd.n13743 vdd.n8792 1.882
R52411 vdd.n13937 vdd.n8637 1.882
R52412 vdd.n13946 vdd.n13942 1.882
R52413 vdd.n14018 vdd.n8584 1.882
R52414 vdd.n14025 vdd.n14024 1.882
R52415 vdd.n14227 vdd.n8415 1.882
R52416 vdd.n14236 vdd.n14232 1.882
R52417 vdd.n14307 vdd.n8362 1.882
R52418 vdd.n14317 vdd.n8359 1.882
R52419 vdd.n14557 vdd.n8191 1.882
R52420 vdd.n14552 vdd.n8192 1.882
R52421 vdd.n24276 vdd.n24269 1.882
R52422 vdd.n24278 vdd.n24276 1.882
R52423 vdd.n24173 vdd.n24166 1.882
R52424 vdd.n24007 vdd.n24000 1.882
R52425 vdd.n23941 vdd.n23934 1.882
R52426 vdd.n23775 vdd.n23768 1.882
R52427 vdd.n23709 vdd.n23702 1.882
R52428 vdd.n23087 vdd.n23080 1.882
R52429 vdd.n23253 vdd.n23246 1.882
R52430 vdd.n23319 vdd.n23312 1.882
R52431 vdd.n23485 vdd.n23478 1.882
R52432 vdd.n23551 vdd.n23544 1.882
R52433 vdd.n22508 vdd.n22501 1.882
R52434 vdd.n22674 vdd.n22667 1.882
R52435 vdd.n22740 vdd.n22733 1.882
R52436 vdd.n22906 vdd.n22899 1.882
R52437 vdd.n22972 vdd.n22965 1.882
R52438 vdd.n22448 vdd.n22441 1.882
R52439 vdd.n22450 vdd.n22448 1.882
R52440 vdd.n22254 vdd.n22253 1.882
R52441 vdd.n22253 vdd.n22245 1.882
R52442 vdd.n22304 vdd.n22297 1.882
R52443 vdd.n22306 vdd.n22304 1.882
R52444 vdd.n22130 vdd.n22129 1.882
R52445 vdd.n22129 vdd.n22121 1.882
R52446 vdd.n19376 vdd.n19375 1.882
R52447 vdd.n19457 vdd.n19456 1.882
R52448 vdd.n19582 vdd.n19581 1.882
R52449 vdd.n19657 vdd.n19656 1.882
R52450 vdd.n19784 vdd.n19783 1.882
R52451 vdd.n20981 vdd.n20980 1.882
R52452 vdd.n19883 vdd.n19882 1.882
R52453 vdd.n20790 vdd.n20789 1.882
R52454 vdd.n20666 vdd.n20665 1.882
R52455 vdd.n20585 vdd.n20584 1.882
R52456 vdd.n21601 vdd.n21600 1.882
R52457 vdd.n21423 vdd.n21422 1.882
R52458 vdd.n21342 vdd.n21341 1.882
R52459 vdd.n21164 vdd.n21163 1.882
R52460 vdd.n21090 vdd.n21089 1.882
R52461 vdd.n19057 vdd.n19056 1.882
R52462 vdd.n18976 vdd.n18975 1.882
R52463 vdd.n18798 vdd.n18797 1.882
R52464 vdd.n18717 vdd.n18716 1.882
R52465 vdd.n18539 vdd.n18538 1.882
R52466 vdd.n20468 vdd.n19982 1.882
R52467 vdd.n20468 vdd.n19985 1.882
R52468 vdd.n20300 vdd.n20291 1.882
R52469 vdd.n20250 vdd.n20241 1.882
R52470 vdd.n20064 vdd.n20028 1.882
R52471 vdd.n24680 vdd.n24675 1.882
R52472 vdd.n24817 vdd.n24812 1.882
R52473 vdd.n25235 vdd.n25230 1.882
R52474 vdd.n25098 vdd.n25093 1.882
R52475 vdd.n11921 vdd.n11920 1.866
R52476 vdd.n11920 vdd.n9285 1.866
R52477 vdd.n21743 vdd.n15003 1.866
R52478 vdd.n21745 vdd.n21743 1.866
R52479 vdd.n25396 vdd.n25381 1.861
R52480 vdd.n25396 vdd.n25386 1.86
R52481 vdd.n24512 vdd.n24511 1.853
R52482 vdd.n25255 vdd.n14975 1.845
R52483 vdd.n35698 vdd.n35697 1.844
R52484 vdd.n35698 vdd.n35696 1.844
R52485 vdd.n35698 vdd.n35695 1.844
R52486 vdd.n35698 vdd.n35694 1.844
R52487 vdd.n27223 vdd.n27222 1.844
R52488 vdd.n27218 vdd.n27217 1.844
R52489 vdd.n28830 vdd.n28829 1.844
R52490 vdd.n28830 vdd.n28828 1.844
R52491 vdd.n28830 vdd.n28827 1.844
R52492 vdd.n28824 vdd.n28822 1.844
R52493 vdd.n28824 vdd.n28821 1.844
R52494 vdd.n28824 vdd.n28823 1.844
R52495 vdd.n25396 vdd.n25382 1.844
R52496 vdd.n3669 vdd.n3666 1.844
R52497 vdd.n3669 vdd.n3665 1.844
R52498 vdd.n3663 vdd.n3660 1.844
R52499 vdd.n3663 vdd.n3659 1.844
R52500 vdd.n27223 vdd.n27221 1.844
R52501 vdd.n27223 vdd.n27220 1.844
R52502 vdd.n27218 vdd.n27216 1.844
R52503 vdd.n27218 vdd.n27215 1.844
R52504 vdd.n25024 vdd.n25023 1.844
R52505 vdd.n35692 vdd.n35688 1.844
R52506 vdd.n35692 vdd.n35689 1.844
R52507 vdd.n35692 vdd.n35690 1.844
R52508 vdd.n35692 vdd.n35691 1.844
R52509 vdd.n32385 vdd.n32384 1.843
R52510 vdd.n9131 vdd.n9103 1.835
R52511 vdd.n9105 vdd.n9104 1.835
R52512 vdd.n13410 vdd.n9032 1.835
R52513 vdd.n13521 vdd.n8969 1.835
R52514 vdd.n8909 vdd.n8882 1.835
R52515 vdd.n8884 vdd.n8883 1.835
R52516 vdd.n13704 vdd.n13703 1.835
R52517 vdd.n13793 vdd.n13792 1.835
R52518 vdd.n13871 vdd.t330 1.835
R52519 vdd.n13888 vdd.n8695 1.835
R52520 vdd.n13927 vdd.n8646 1.835
R52521 vdd.n8600 vdd.n8588 1.835
R52522 vdd.n14080 vdd.n14079 1.835
R52523 vdd.n14177 vdd.n8472 1.835
R52524 vdd.n14217 vdd.n8426 1.835
R52525 vdd.n14277 vdd.n8378 1.835
R52526 vdd.n14381 vdd.n8312 1.835
R52527 vdd.n8233 vdd.n8222 1.835
R52528 vdd.n8224 vdd.n8223 1.835
R52529 vdd.n8141 vdd.t305 1.835
R52530 vdd.n35855 vdd.n35854 1.788
R52531 vdd.n35988 vdd.n35987 1.788
R52532 vdd.n36086 vdd.n36085 1.788
R52533 vdd.n36219 vdd.n36218 1.788
R52534 vdd.n36317 vdd.n36316 1.788
R52535 vdd.n36450 vdd.n36449 1.788
R52536 vdd.n36548 vdd.n36547 1.788
R52537 vdd.n36681 vdd.n36680 1.788
R52538 vdd.n36779 vdd.n36778 1.788
R52539 vdd.n36912 vdd.n36911 1.788
R52540 vdd.n3633 vdd.n3632 1.788
R52541 vdd.n33195 vdd.n33194 1.788
R52542 vdd.n37204 vdd.n37203 1.788
R52543 vdd.n2378 vdd.n2377 1.788
R52544 vdd.n32959 vdd.n32958 1.788
R52545 vdd.n1906 vdd.n1905 1.788
R52546 vdd.n1271 vdd.n1270 1.788
R52547 vdd.n38065 vdd.n38064 1.788
R52548 vdd.n37967 vdd.n37966 1.788
R52549 vdd.n37834 vdd.n37833 1.788
R52550 vdd.n37736 vdd.n37735 1.788
R52551 vdd.n37603 vdd.n37602 1.788
R52552 vdd.n28276 vdd.n28275 1.788
R52553 vdd.n28409 vdd.n28408 1.788
R52554 vdd.n28507 vdd.n28506 1.788
R52555 vdd.n28640 vdd.n28639 1.788
R52556 vdd.n28738 vdd.n28737 1.788
R52557 vdd.n28811 vdd.n28810 1.788
R52558 vdd.n28063 vdd.n28062 1.788
R52559 vdd.n31658 vdd.n31654 1.788
R52560 vdd.n32122 vdd.n32121 1.788
R52561 vdd.n29763 vdd.n29762 1.788
R52562 vdd.n30235 vdd.n30234 1.788
R52563 vdd.n30339 vdd.n30338 1.788
R52564 vdd.n10472 vdd.n10274 1.776
R52565 vdd.n15266 vdd.n15265 1.776
R52566 vdd.n1794 vdd.n1793 1.767
R52567 vdd.n2475 vdd.n2474 1.767
R52568 vdd.n19398 vdd.n19395 1.759
R52569 vdd.t242 vdd.n19417 1.759
R52570 vdd.n19447 vdd.n19444 1.759
R52571 vdd.n19589 vdd.t164 1.759
R52572 vdd.n19604 vdd.n19601 1.759
R52573 vdd.n19647 vdd.n19644 1.759
R52574 vdd.n19806 vdd.n19803 1.759
R52575 vdd.n19156 vdd.n19153 1.759
R52576 vdd.n20855 vdd.n20852 1.759
R52577 vdd.n20812 vdd.n20809 1.759
R52578 vdd.n20797 vdd.t174 1.759
R52579 vdd.n20656 vdd.n20653 1.759
R52580 vdd.n20607 vdd.n20604 1.759
R52581 vdd.n20282 vdd.n20281 1.759
R52582 vdd.n20264 vdd.n20263 1.759
R52583 vdd.n8087 vdd.n8072 1.754
R52584 vdd.n14802 vdd.n14801 1.754
R52585 vdd.n1869 vdd.n1867 1.738
R52586 vdd.n11915 vdd.n11914 1.729
R52587 vdd.n22001 vdd.n22000 1.729
R52588 vdd.n2420 vdd.n2416 1.706
R52589 vdd.n3854 vdd.n3848 1.706
R52590 vdd.n10473 vdd.n10472 1.702
R52591 vdd.n15265 vdd.n15264 1.702
R52592 vdd.n3723 vdd.n3722 1.69
R52593 vdd.n11617 vdd.n11616 1.69
R52594 vdd.n3821 vdd.n3820 1.688
R52595 vdd.n12585 vdd.n12584 1.659
R52596 vdd.n12601 vdd.n10066 1.659
R52597 vdd.n10408 vdd.n10322 1.659
R52598 vdd.n10408 vdd.n10407 1.659
R52599 vdd.n13077 vdd.n13076 1.659
R52600 vdd.n13076 vdd.n9294 1.659
R52601 vdd.n13017 vdd.n13016 1.659
R52602 vdd.n13016 vdd.n9395 1.659
R52603 vdd.n12965 vdd.n9460 1.659
R52604 vdd.n12965 vdd.n9461 1.659
R52605 vdd.n9586 vdd.n9585 1.659
R52606 vdd.n9586 vdd.n9581 1.659
R52607 vdd.n12869 vdd.n12868 1.659
R52608 vdd.n12868 vdd.n9626 1.659
R52609 vdd.n12809 vdd.n12808 1.659
R52610 vdd.n12808 vdd.n9755 1.659
R52611 vdd.n12757 vdd.n9820 1.659
R52612 vdd.n12757 vdd.n9821 1.659
R52613 vdd.n9946 vdd.n9945 1.659
R52614 vdd.n9946 vdd.n9941 1.659
R52615 vdd.n12661 vdd.n12660 1.659
R52616 vdd.n12660 vdd.n9986 1.659
R52617 vdd.n10556 vdd.n10535 1.659
R52618 vdd.n12505 vdd.n10533 1.659
R52619 vdd.n10638 vdd.n10633 1.659
R52620 vdd.n10643 vdd.n10629 1.659
R52621 vdd.n10711 vdd.n10703 1.659
R52622 vdd.n10735 vdd.n10729 1.659
R52623 vdd.n12361 vdd.n10778 1.659
R52624 vdd.n12356 vdd.n10805 1.659
R52625 vdd.n12315 vdd.n12314 1.659
R52626 vdd.n12301 vdd.n10898 1.659
R52627 vdd.n10988 vdd.n10987 1.659
R52628 vdd.n12261 vdd.n10963 1.659
R52629 vdd.n11067 vdd.n11041 1.659
R52630 vdd.n11080 vdd.n11060 1.659
R52631 vdd.n12154 vdd.n11134 1.659
R52632 vdd.n11160 vdd.n11159 1.659
R52633 vdd.n12101 vdd.n11219 1.659
R52634 vdd.n12094 vdd.n12093 1.659
R52635 vdd.n12055 vdd.n11286 1.659
R52636 vdd.n12050 vdd.n11314 1.659
R52637 vdd.n12009 vdd.n12008 1.659
R52638 vdd.n11995 vdd.n11407 1.659
R52639 vdd.n11535 vdd.n11454 1.659
R52640 vdd.n11955 vdd.n11448 1.659
R52641 vdd.n15047 vdd.n15046 1.659
R52642 vdd.n15384 vdd.n15383 1.659
R52643 vdd.n15383 vdd.n15376 1.659
R52644 vdd.n15463 vdd.n15450 1.659
R52645 vdd.n15465 vdd.n15463 1.659
R52646 vdd.n15629 vdd.n15628 1.659
R52647 vdd.n15628 vdd.n15618 1.659
R52648 vdd.n15719 vdd.n15706 1.659
R52649 vdd.n15721 vdd.n15719 1.659
R52650 vdd.n15885 vdd.n15884 1.659
R52651 vdd.n15884 vdd.n15874 1.659
R52652 vdd.n15975 vdd.n15962 1.659
R52653 vdd.n15977 vdd.n15975 1.659
R52654 vdd.n16141 vdd.n16140 1.659
R52655 vdd.n16140 vdd.n16130 1.659
R52656 vdd.n16231 vdd.n16218 1.659
R52657 vdd.n16233 vdd.n16231 1.659
R52658 vdd.n16397 vdd.n16396 1.659
R52659 vdd.n16396 vdd.n16386 1.659
R52660 vdd.n16487 vdd.n16474 1.659
R52661 vdd.n16489 vdd.n16487 1.659
R52662 vdd.n16892 vdd.n16891 1.659
R52663 vdd.n16934 vdd.n16933 1.659
R52664 vdd.n17043 vdd.n17041 1.659
R52665 vdd.n17048 vdd.n17047 1.659
R52666 vdd.n17164 vdd.n17163 1.659
R52667 vdd.n17206 vdd.n17205 1.659
R52668 vdd.n17315 vdd.n17313 1.659
R52669 vdd.n17320 vdd.n17319 1.659
R52670 vdd.n17436 vdd.n17435 1.659
R52671 vdd.n17478 vdd.n17477 1.659
R52672 vdd.n17587 vdd.n17585 1.659
R52673 vdd.n16831 vdd.n16830 1.659
R52674 vdd.n17694 vdd.n17693 1.659
R52675 vdd.n17736 vdd.n17735 1.659
R52676 vdd.n17845 vdd.n17843 1.659
R52677 vdd.n17850 vdd.n17849 1.659
R52678 vdd.n17965 vdd.n17964 1.659
R52679 vdd.n18007 vdd.n18006 1.659
R52680 vdd.n18116 vdd.n18114 1.659
R52681 vdd.n18121 vdd.n18120 1.659
R52682 vdd.n18236 vdd.n18235 1.659
R52683 vdd.n18275 vdd.n18274 1.659
R52684 vdd.n18380 vdd.n18379 1.659
R52685 vdd.n3805 vdd.n3804 1.632
R52686 vdd.n2415 vdd.n2414 1.621
R52687 vdd.n31471 vdd.n31470 1.615
R52688 vdd.n32026 vdd.n32025 1.615
R52689 vdd.n31620 vdd.n31619 1.615
R52690 vdd.n26614 vdd.n26613 1.615
R52691 vdd.n26340 vdd.n26339 1.614
R52692 vdd.n33621 vdd.n33620 1.614
R52693 vdd.n1097 vdd.n1096 1.614
R52694 vdd.n120 vdd.n119 1.614
R52695 vdd.n25426 vdd.n25425 1.614
R52696 vdd.n25665 vdd.n25664 1.614
R52697 vdd.n10403 vdd.n10326 1.613
R52698 vdd.n10368 vdd.n9289 1.604
R52699 vdd.n9407 vdd.n9406 1.604
R52700 vdd.n9434 vdd.t294 1.604
R52701 vdd.n12973 vdd.n12972 1.604
R52702 vdd.n9596 vdd.n9595 1.604
R52703 vdd.n9649 vdd.n9621 1.604
R52704 vdd.n9767 vdd.n9766 1.604
R52705 vdd.n12765 vdd.n12764 1.604
R52706 vdd.n9956 vdd.n9955 1.604
R52707 vdd.n10009 vdd.n9981 1.604
R52708 vdd.n12595 vdd.n10102 1.604
R52709 vdd.n12567 vdd.n10479 1.604
R52710 vdd.n12519 vdd.n10523 1.604
R52711 vdd.t311 vdd.n12501 1.604
R52712 vdd.n12453 vdd.n10622 1.604
R52713 vdd.n12414 vdd.n12413 1.604
R52714 vdd.n10816 vdd.n10807 1.604
R52715 vdd.n10886 vdd.n10885 1.604
R52716 vdd.n12253 ldomc_0.otaldom_0.pmoslm_0.vdd 1.604
R52717 vdd.n12253 vdd.n12252 1.604
R52718 vdd.n11050 vdd.n11045 1.604
R52719 vdd.n11169 vdd.n11168 1.604
R52720 vdd.n12115 vdd.n11192 1.604
R52721 vdd.n11325 vdd.n11316 1.604
R52722 vdd.n11395 vdd.n11394 1.604
R52723 vdd.n11946 vdd.n11945 1.604
R52724 vdd.n15441 vdd.n15440 1.604
R52725 vdd.n15643 vdd.n15642 1.604
R52726 vdd.n15660 vdd.t266 1.604
R52727 vdd.n15697 vdd.n15696 1.604
R52728 vdd.n15899 vdd.n15898 1.604
R52729 vdd.n15953 vdd.n15952 1.604
R52730 vdd.n16155 vdd.n16154 1.604
R52731 vdd.n16209 vdd.n16208 1.604
R52732 vdd.n16411 vdd.n16410 1.604
R52733 vdd.n16465 vdd.n16464 1.604
R52734 vdd.n16633 vdd.n16632 1.604
R52735 vdd.n15116 vdd.n15085 1.604
R52736 vdd.n16882 vdd.n16879 1.604
R52737 vdd.t252 vdd.n16927 1.604
R52738 vdd.n17070 vdd.n17067 1.604
R52739 vdd.n17154 vdd.n17151 1.604
R52740 vdd.n17342 vdd.n17339 1.604
R52741 vdd.n17426 vdd.n17423 1.604
R52742 vdd.n17597 bandgapmd_0.otam_1.pmoslm_0.vdd 1.604
R52743 vdd.n17600 vdd.n17597 1.604
R52744 vdd.n17684 vdd.n17681 1.604
R52745 vdd.n17872 vdd.n17869 1.604
R52746 vdd.n17955 vdd.n17952 1.604
R52747 vdd.n18143 vdd.n18140 1.604
R52748 vdd.n18226 vdd.n18224 1.604
R52749 vdd.n15008 vdd.n15007 1.604
R52750 vdd.n15395 vdd.n15394 1.601
R52751 vdd.n32070 vdd.n32069 1.6
R52752 vdd.n13152 vdd.n9212 1.599
R52753 vdd.n13188 vdd.n13187 1.599
R52754 vdd.n27888 vdd.n27887 1.593
R52755 vdd.n27845 vdd.n27844 1.593
R52756 vdd.n2384 vdd.n2380 1.587
R52757 vdd.n2043 vdd.n2040 1.587
R52758 vdd.n2197 vdd.n2196 1.587
R52759 vdd.n2017 vdd.n2014 1.587
R52760 vdd.n2057 vdd.n2056 1.587
R52761 vdd.n32497 vdd.n32496 1.578
R52762 vdd.n24522 vdd.n24521 1.577
R52763 vdd.n31463 vdd.n31451 1.571
R52764 vdd.n30244 vdd.n30243 1.567
R52765 vdd.n32058 vdd.n32057 1.566
R52766 vdd.n35868 vdd.n35867 1.564
R52767 vdd.n35973 vdd.n35972 1.564
R52768 vdd.n36099 vdd.n36098 1.564
R52769 vdd.n36204 vdd.n36203 1.564
R52770 vdd.n36330 vdd.n36329 1.564
R52771 vdd.n36435 vdd.n36434 1.564
R52772 vdd.n36561 vdd.n36560 1.564
R52773 vdd.n36666 vdd.n36665 1.564
R52774 vdd.n36792 vdd.n36791 1.564
R52775 vdd.n36897 vdd.n36896 1.564
R52776 vdd.n2053 vdd.n2052 1.564
R52777 vdd.n2011 vdd.n2010 1.564
R52778 vdd.n2193 vdd.n2192 1.564
R52779 vdd.n2037 vdd.n2036 1.564
R52780 vdd.n37406 vdd.n37405 1.564
R52781 vdd.n1194 vdd.n1193 1.564
R52782 vdd.n1281 vdd.n1280 1.564
R52783 vdd.n38078 vdd.n38077 1.564
R52784 vdd.n37952 vdd.n37951 1.564
R52785 vdd.n37847 vdd.n37846 1.564
R52786 vdd.n37721 vdd.n37720 1.564
R52787 vdd.n37616 vdd.n37615 1.564
R52788 vdd.n28289 vdd.n28288 1.564
R52789 vdd.n28394 vdd.n28393 1.564
R52790 vdd.n28520 vdd.n28519 1.564
R52791 vdd.n28625 vdd.n28624 1.564
R52792 vdd.n28751 vdd.n28750 1.564
R52793 vdd.n28137 vdd.n28136 1.564
R52794 vdd.n28965 vdd.n28964 1.564
R52795 vdd.n27808 vdd.n27807 1.564
R52796 vdd.n32155 vdd.n32154 1.564
R52797 vdd.n31508 vdd.n31507 1.564
R52798 vdd.n32443 vdd.n32442 1.564
R52799 vdd.n31274 vdd.n31273 1.564
R52800 vdd.n27846 vdd.n27845 1.552
R52801 vdd.n13287 vdd.n9150 1.529
R52802 vdd.t106 vdd.n9151 1.529
R52803 vdd.n13365 vdd.n9071 1.529
R52804 vdd.n13445 vdd.n8992 1.529
R52805 vdd.n13482 vdd.n13481 1.529
R52806 vdd.t126 vdd.n8957 1.529
R52807 vdd.n13568 vdd.t283 1.529
R52808 vdd.n13579 vdd.n8929 1.529
R52809 vdd.n13657 vdd.n8851 1.529
R52810 vdd.n13736 vdd.n8776 1.529
R52811 vdd.n13762 vdd.n13761 1.529
R52812 vdd.n13833 vdd.t285 1.529
R52813 vdd.n13864 vdd.t112 1.529
R52814 vdd.n8721 vdd.n8707 1.529
R52815 vdd.n13935 vdd.n13934 1.529
R52816 vdd.n14052 vdd.n8574 1.529
R52817 vdd.n14068 vdd.n8560 1.529
R52818 vdd.n14069 vdd.t290 1.529
R52819 vdd.n14118 vdd.t122 1.529
R52820 vdd.n8525 vdd.t329 1.529
R52821 vdd.n8500 vdd.n8484 1.529
R52822 vdd.n14225 vdd.n14224 1.529
R52823 vdd.n14327 vdd.n8357 1.529
R52824 vdd.n14345 vdd.n8318 1.529
R52825 vdd.t333 vdd.n8333 1.529
R52826 vdd.n14438 vdd.n14437 1.529
R52827 vdd.n14559 vdd.n8187 1.529
R52828 vdd.n14656 vdd.n8146 1.529
R52829 vdd.n14644 vdd.n8160 1.529
R52830 vdd.n24627 vdd.n24567 1.515
R52831 vdd.n33735 vdd.n33734 1.505
R52832 vdd.n33733 vdd.n33732 1.505
R52833 vdd.n33489 vdd.n33488 1.505
R52834 vdd.n33345 vdd.n33344 1.505
R52835 vdd.n33399 vdd.n33398 1.505
R52836 vdd.n34205 vdd.n34204 1.505
R52837 vdd.n34096 vdd.n34095 1.505
R52838 vdd.n33981 vdd.n33980 1.505
R52839 vdd.n34386 vdd.n34385 1.505
R52840 vdd.n34387 vdd.n34386 1.505
R52841 vdd.n35143 vdd.n35142 1.505
R52842 vdd.n35405 vdd.n35404 1.505
R52843 vdd.n35406 vdd.n35405 1.505
R52844 vdd.n35257 vdd.n35256 1.505
R52845 vdd.n35289 vdd.n35288 1.505
R52846 vdd.n34705 vdd.n34704 1.505
R52847 vdd.n34673 vdd.n34672 1.505
R52848 vdd.n34556 vdd.n34555 1.505
R52849 vdd.n34809 vdd.n34808 1.505
R52850 vdd.n34810 vdd.n34809 1.505
R52851 vdd.n936 vdd.n935 1.505
R52852 vdd.n934 vdd.n933 1.505
R52853 vdd.n976 vdd.n975 1.505
R52854 vdd.n611 vdd.n610 1.505
R52855 vdd.n718 vdd.n717 1.505
R52856 vdd.n315 vdd.n314 1.505
R52857 vdd.n168 vdd.n167 1.505
R52858 vdd.n182 vdd.n181 1.505
R52859 vdd.n449 vdd.n448 1.505
R52860 vdd.n516 vdd.n515 1.505
R52861 vdd.n6266 vdd.n6265 1.505
R52862 vdd.n6099 vdd.n6098 1.505
R52863 vdd.n6100 vdd.n6099 1.505
R52864 vdd.n5801 vdd.n5800 1.505
R52865 vdd.n5906 vdd.n5905 1.505
R52866 vdd.n5452 vdd.n5451 1.505
R52867 vdd.n5420 vdd.n5419 1.505
R52868 vdd.n5303 vdd.n5302 1.505
R52869 vdd.n5556 vdd.n5555 1.505
R52870 vdd.n5557 vdd.n5556 1.505
R52871 vdd.n4751 vdd.n4750 1.505
R52872 vdd.n4750 vdd.n4749 1.505
R52873 vdd.n5160 vdd.n5159 1.505
R52874 vdd.n5079 vdd.n5078 1.505
R52875 vdd.n4932 vdd.n4931 1.505
R52876 vdd.n4279 vdd.n4278 1.505
R52877 vdd.n4250 vdd.n4249 1.505
R52878 vdd.n4133 vdd.n4132 1.505
R52879 vdd.n4382 vdd.n4381 1.505
R52880 vdd.n4383 vdd.n4382 1.505
R52881 vdd.n30200 vdd.n30198 1.505
R52882 vdd.n30229 vdd.n30228 1.505
R52883 vdd.n30253 vdd.n30252 1.505
R52884 vdd.n30243 vdd.n30242 1.505
R52885 vdd.n31450 vdd.n31449 1.505
R52886 vdd.n32291 vdd.n32290 1.505
R52887 vdd.n32102 vdd.n32101 1.505
R52888 vdd.n31922 vdd.n31921 1.505
R52889 vdd.n31041 vdd.n31040 1.505
R52890 vdd.n31285 vdd.n31284 1.505
R52891 vdd.n36018 vdd.n36011 1.505
R52892 vdd.n36060 vdd.n36053 1.505
R52893 vdd.n36249 vdd.n36242 1.505
R52894 vdd.n36291 vdd.n36284 1.505
R52895 vdd.n36480 vdd.n36473 1.505
R52896 vdd.n36522 vdd.n36515 1.505
R52897 vdd.n36711 vdd.n36704 1.505
R52898 vdd.n36753 vdd.n36746 1.505
R52899 vdd.n36942 vdd.n36935 1.505
R52900 vdd.n35686 vdd.n35682 1.505
R52901 vdd.n37150 vdd.n37143 1.505
R52902 vdd.n37178 vdd.n37171 1.505
R52903 vdd.n32991 vdd.n32984 1.505
R52904 vdd.n32977 vdd.n32970 1.505
R52905 vdd.n37525 vdd.n37518 1.505
R52906 vdd.n37571 vdd.n37564 1.505
R52907 vdd.n38039 vdd.n38032 1.505
R52908 vdd.n37997 vdd.n37990 1.505
R52909 vdd.n37808 vdd.n37801 1.505
R52910 vdd.n37766 vdd.n37759 1.505
R52911 vdd.n28208 vdd.n28201 1.505
R52912 vdd.n28250 vdd.n28243 1.505
R52913 vdd.n28439 vdd.n28432 1.505
R52914 vdd.n28481 vdd.n28474 1.505
R52915 vdd.n28670 vdd.n28663 1.505
R52916 vdd.n28712 vdd.n28705 1.505
R52917 vdd.n28115 vdd.n28108 1.505
R52918 vdd.n28089 vdd.n28082 1.505
R52919 vdd.n28071 vdd.n28070 1.505
R52920 vdd.n28968 vdd.n28961 1.505
R52921 vdd.n27800 vdd.n27799 1.505
R52922 vdd.n27916 vdd.n27915 1.505
R52923 vdd.n29860 vdd.n29859 1.505
R52924 vdd.n29723 vdd.n29716 1.505
R52925 vdd.n30192 vdd.n30191 1.505
R52926 vdd.n27341 vdd.n27340 1.505
R52927 vdd.n27371 vdd.n27370 1.505
R52928 vdd.n27497 vdd.n27496 1.505
R52929 vdd.n27498 vdd.n27497 1.505
R52930 vdd.n27259 vdd.n27258 1.505
R52931 vdd.n25793 vdd.n25792 1.505
R52932 vdd.n25739 vdd.n25738 1.505
R52933 vdd.n25934 vdd.n25933 1.505
R52934 vdd.n25935 vdd.n25934 1.505
R52935 vdd.n26027 vdd.n26026 1.505
R52936 vdd.n25522 vdd.n25521 1.505
R52937 vdd.n25620 vdd.n25618 1.505
R52938 vdd.n25402 vdd.n25401 1.505
R52939 vdd.n26300 vdd.n26299 1.505
R52940 vdd.n1670 vdd.n1666 1.505
R52941 vdd.n1638 vdd.n1634 1.505
R52942 vdd.n1489 vdd.n1485 1.505
R52943 vdd.n1457 vdd.n1453 1.505
R52944 vdd.n1308 vdd.n1304 1.505
R52945 vdd.n26774 vdd.n26770 1.505
R52946 vdd.n26923 vdd.n26919 1.505
R52947 vdd.n26955 vdd.n26951 1.505
R52948 vdd.n27104 vdd.n27100 1.505
R52949 vdd.n27136 vdd.n27132 1.505
R52950 vdd.n2876 vdd.n2872 1.505
R52951 vdd.n2908 vdd.n2904 1.505
R52952 vdd.n3057 vdd.n3053 1.505
R52953 vdd.n3089 vdd.n3085 1.505
R52954 vdd.n3238 vdd.n3234 1.505
R52955 vdd.n3270 vdd.n3266 1.505
R52956 vdd.n3419 vdd.n3415 1.505
R52957 vdd.n3451 vdd.n3447 1.505
R52958 vdd.n3600 vdd.n3596 1.505
R52959 vdd.n3645 vdd.n3638 1.505
R52960 vdd.n31726 vdd.n31725 1.505
R52961 vdd.n9123 vdd.n9067 1.505
R52962 vdd.n13393 vdd.n9052 1.505
R52963 vdd.n8902 vdd.n8847 1.505
R52964 vdd.n13685 vdd.n8832 1.505
R52965 vdd.n13913 vdd.n8660 1.505
R52966 vdd.n8611 vdd.n8610 1.505
R52967 vdd.n14203 vdd.n8440 1.505
R52968 vdd.n8389 vdd.n8388 1.505
R52969 vdd.n14693 vdd.n8128 1.505
R52970 vdd.n14688 vdd.n8129 1.505
R52971 vdd.n14718 vdd.n14717 1.505
R52972 vdd.n14739 vdd.n14738 1.505
R52973 vdd.n14867 vdd.n8038 1.505
R52974 vdd.n14862 vdd.n8039 1.505
R52975 vdd.n14902 vdd.n8025 1.505
R52976 vdd.n14892 vdd.n14884 1.505
R52977 vdd.n11615 vdd.n9248 1.505
R52978 vdd.n13136 vdd.n9255 1.505
R52979 vdd.n9256 vdd.n9237 1.505
R52980 vdd.n13221 vdd.n9195 1.505
R52981 vdd.n13221 vdd.n9201 1.505
R52982 vdd.n13306 vdd.n9137 1.505
R52983 vdd.n13307 vdd.n13306 1.505
R52984 vdd.n13513 vdd.n8973 1.505
R52985 vdd.n13513 vdd.n8979 1.505
R52986 vdd.n13598 vdd.n8915 1.505
R52987 vdd.n13599 vdd.n13598 1.505
R52988 vdd.n13812 vdd.n8743 1.505
R52989 vdd.n13812 vdd.n8744 1.505
R52990 vdd.n13877 vdd.n8703 1.505
R52991 vdd.n13877 vdd.n8701 1.505
R52992 vdd.n14099 vdd.n8530 1.505
R52993 vdd.n14099 vdd.n8532 1.505
R52994 vdd.n14166 vdd.n8480 1.505
R52995 vdd.n14166 vdd.n8478 1.505
R52996 vdd.n14392 vdd.n8307 1.505
R52997 vdd.n14392 vdd.n8308 1.505
R52998 vdd.n14449 vdd.n8264 1.505
R52999 vdd.n14449 vdd.n8265 1.505
R53000 vdd.n11742 vdd.n11724 1.505
R53001 vdd.n11717 vdd.n11685 1.505
R53002 vdd.n11705 vdd.n11704 1.505
R53003 vdd.n11826 vdd.n11820 1.505
R53004 vdd.n11864 vdd.n11863 1.505
R53005 vdd.n11848 vdd.n11847 1.505
R53006 vdd.n11913 vdd.n11911 1.505
R53007 vdd.n24212 vdd.n24211 1.505
R53008 vdd.n24209 vdd.n24208 1.505
R53009 vdd.n24110 vdd.n24109 1.505
R53010 vdd.n24056 vdd.n24055 1.505
R53011 vdd.n23878 vdd.n23877 1.505
R53012 vdd.n23824 vdd.n23823 1.505
R53013 vdd.n23646 vdd.n23645 1.505
R53014 vdd.n23136 vdd.n23135 1.505
R53015 vdd.n23190 vdd.n23189 1.505
R53016 vdd.n23368 vdd.n23367 1.505
R53017 vdd.n23422 vdd.n23421 1.505
R53018 vdd.n23600 vdd.n23599 1.505
R53019 vdd.n22557 vdd.n22556 1.505
R53020 vdd.n22611 vdd.n22610 1.505
R53021 vdd.n22789 vdd.n22788 1.505
R53022 vdd.n22843 vdd.n22842 1.505
R53023 vdd.n23021 vdd.n23020 1.505
R53024 vdd.n22384 vdd.n22383 1.505
R53025 vdd.n22381 vdd.n22380 1.505
R53026 vdd.n22348 vdd.n22347 1.505
R53027 vdd.n22352 vdd.n22351 1.505
R53028 vdd.n24329 vdd.n24328 1.505
R53029 vdd.n24326 vdd.n24325 1.505
R53030 vdd.n22064 vdd.n22063 1.505
R53031 vdd.n22081 vdd.n22080 1.505
R53032 vdd.n19281 vdd.n19272 1.505
R53033 vdd.n19245 vdd.n19236 1.505
R53034 vdd.n19225 vdd.n19216 1.505
R53035 vdd.n19188 vdd.n19179 1.505
R53036 vdd.n19842 vdd.n19833 1.505
R53037 vdd.n19879 vdd.n19870 1.505
R53038 vdd.n19911 vdd.n19902 1.505
R53039 vdd.n19947 vdd.n19938 1.505
R53040 vdd.n21546 vdd.n21537 1.505
R53041 vdd.n21496 vdd.n21487 1.505
R53042 vdd.n21287 vdd.n21278 1.505
R53043 vdd.n21237 vdd.n21228 1.505
R53044 vdd.n21028 vdd.n21021 1.505
R53045 vdd.n19129 vdd.n19121 1.505
R53046 vdd.n18921 vdd.n18912 1.505
R53047 vdd.n18871 vdd.n18862 1.505
R53048 vdd.n18662 vdd.n18653 1.505
R53049 vdd.n18612 vdd.n18603 1.505
R53050 vdd.n20413 vdd.n20412 1.505
R53051 vdd.n20355 vdd.n20354 1.505
R53052 vdd.n20177 vdd.n20176 1.505
R53053 vdd.n20119 vdd.n20118 1.505
R53054 vdd.n21806 vdd.n21805 1.505
R53055 vdd.n21768 vdd.n21767 1.505
R53056 vdd.n21917 vdd.n21911 1.505
R53057 vdd.n21955 vdd.n21954 1.505
R53058 vdd.n21939 vdd.n21938 1.505
R53059 vdd.n21754 vdd.n21753 1.505
R53060 vdd.n24724 vdd.n24723 1.505
R53061 vdd.n24764 vdd.n24763 1.505
R53062 vdd.n25182 vdd.n25181 1.505
R53063 vdd.n25142 vdd.n25141 1.505
R53064 vdd.n32536 vdd.n32535 1.5
R53065 vdd.n11493 vdd.n11465 1.5
R53066 vdd.n11500 vdd.n11499 1.5
R53067 vdd.n11510 vdd.n11509 1.5
R53068 vdd.n11512 vdd.n11455 1.5
R53069 vdd.n11540 vdd.n11539 1.5
R53070 vdd.n11544 vdd.n11542 1.5
R53071 vdd.n11590 vdd.n11589 1.5
R53072 vdd.n11585 vdd.n11584 1.5
R53073 vdd.n10175 vdd.n10174 1.5
R53074 vdd.n21700 vdd.n21699 1.5
R53075 vdd.n31239 vdd.n31188 1.5
R53076 vdd.n31290 vdd.n31289 1.499
R53077 vdd.n12572 vdd.n10259 1.492
R53078 vdd.n10135 vdd.n10087 1.492
R53079 vdd.n16794 vdd.n15122 1.492
R53080 vdd.n25640 vdd.n25639 1.472
R53081 vdd.n32030 vdd.n32026 1.444
R53082 vdd.n10193 vdd.n10137 1.422
R53083 vdd.n10471 vdd.n10470 1.422
R53084 vdd.n10285 vdd.n10284 1.422
R53085 vdd.n10426 vdd.n10425 1.422
R53086 vdd.n10316 vdd.n10311 1.422
R53087 vdd.n13063 vdd.n9306 1.422
R53088 vdd.n13056 vdd.n9310 1.422
R53089 vdd.n9380 vdd.n9371 1.422
R53090 vdd.n9389 vdd.n9388 1.422
R53091 vdd.n9501 vdd.n9481 1.422
R53092 vdd.n9503 vdd.n9478 1.422
R53093 vdd.n12923 vdd.n12922 1.422
R53094 vdd.n12915 vdd.n9550 1.422
R53095 vdd.n12855 vdd.n9666 1.422
R53096 vdd.n12848 vdd.n9671 1.422
R53097 vdd.n9740 vdd.n9731 1.422
R53098 vdd.n9749 vdd.n9748 1.422
R53099 vdd.n9861 vdd.n9841 1.422
R53100 vdd.n9863 vdd.n9838 1.422
R53101 vdd.n12715 vdd.n12714 1.422
R53102 vdd.n12707 vdd.n9910 1.422
R53103 vdd.n12647 vdd.n10026 1.422
R53104 vdd.n12640 vdd.n10031 1.422
R53105 vdd.n12619 vdd.n12618 1.422
R53106 vdd.n10194 vdd.n10086 1.422
R53107 vdd.n10546 vdd.n10538 1.422
R53108 vdd.n12505 vdd.n10562 1.422
R53109 vdd.n12463 vdd.n10610 1.422
R53110 vdd.n12446 vdd.n10627 1.422
R53111 vdd.n12410 vdd.n12409 1.422
R53112 vdd.n10735 vdd.n10726 1.422
R53113 vdd.n10800 vdd.n10780 1.422
R53114 vdd.n10835 vdd.n10813 1.422
R53115 vdd.n10890 vdd.n10889 1.422
R53116 vdd.n10907 vdd.n10898 1.422
R53117 vdd.n10976 vdd.n10975 1.422
R53118 vdd.n12248 vdd.n10996 1.422
R53119 vdd.n12214 vdd.n12213 1.422
R53120 vdd.n12201 vdd.n11060 1.422
R53121 vdd.n12159 vdd.n11126 1.422
R53122 vdd.n11173 vdd.n11172 1.422
R53123 vdd.n12111 vdd.n11196 1.422
R53124 vdd.n12093 vdd.n11226 1.422
R53125 vdd.n11309 vdd.n11288 1.422
R53126 vdd.n11344 vdd.n11322 1.422
R53127 vdd.n11399 vdd.n11398 1.422
R53128 vdd.n11416 vdd.n11407 1.422
R53129 vdd.n11954 vdd.n11449 1.422
R53130 vdd.n16728 vdd.n16724 1.422
R53131 vdd.n15268 vdd.n15267 1.422
R53132 vdd.n15277 vdd.n15276 1.422
R53133 vdd.n15356 vdd.n15345 1.422
R53134 vdd.n15347 vdd.n15346 1.422
R53135 vdd.n15487 vdd.n15486 1.422
R53136 vdd.n15499 vdd.n15498 1.422
R53137 vdd.n15595 vdd.n15582 1.422
R53138 vdd.n15584 vdd.n15583 1.422
R53139 vdd.n15743 vdd.n15742 1.422
R53140 vdd.n15755 vdd.n15754 1.422
R53141 vdd.n15851 vdd.n15838 1.422
R53142 vdd.n15840 vdd.n15839 1.422
R53143 vdd.n15999 vdd.n15998 1.422
R53144 vdd.n16011 vdd.n16010 1.422
R53145 vdd.n16107 vdd.n16094 1.422
R53146 vdd.n16096 vdd.n16095 1.422
R53147 vdd.n16255 vdd.n16254 1.422
R53148 vdd.n16267 vdd.n16266 1.422
R53149 vdd.n16363 vdd.n16350 1.422
R53150 vdd.n16352 vdd.n16351 1.422
R53151 vdd.n16511 vdd.n16510 1.422
R53152 vdd.n16523 vdd.n16522 1.422
R53153 vdd.n16751 vdd.n16746 1.422
R53154 vdd.n16729 vdd.n16723 1.422
R53155 vdd.n16902 vdd.n16890 1.422
R53156 vdd.n16933 vdd.n16924 1.422
R53157 vdd.n17025 vdd.n17016 1.422
R53158 vdd.n17075 vdd.n17074 1.422
R53159 vdd.n17174 vdd.n17162 1.422
R53160 vdd.n17205 vdd.n17196 1.422
R53161 vdd.n17297 vdd.n17288 1.422
R53162 vdd.n17347 vdd.n17346 1.422
R53163 vdd.n17446 vdd.n17434 1.422
R53164 vdd.n17477 vdd.n17468 1.422
R53165 vdd.n17569 vdd.n17560 1.422
R53166 vdd.n17605 vdd.n17604 1.422
R53167 vdd.n17704 vdd.n17692 1.422
R53168 vdd.n17735 vdd.n17726 1.422
R53169 vdd.n17827 vdd.n17818 1.422
R53170 vdd.n17876 vdd.n17875 1.422
R53171 vdd.n17975 vdd.n17963 1.422
R53172 vdd.n18006 vdd.n17997 1.422
R53173 vdd.n18098 vdd.n18089 1.422
R53174 vdd.n18148 vdd.n18147 1.422
R53175 vdd.n18245 vdd.n18234 1.422
R53176 vdd.n18274 vdd.n18266 1.422
R53177 vdd.n24926 vdd.n24925 1.414
R53178 vdd.n21572 vdd.t246 1.407
R53179 vdd.n21528 vdd.n21527 1.407
R53180 vdd.n21510 vdd.n21509 1.407
R53181 vdd.t278 vdd.n21297 1.407
R53182 vdd.n21269 vdd.n21268 1.407
R53183 vdd.n21251 vdd.n21250 1.407
R53184 vdd.n19151 vdd.n19147 1.407
R53185 vdd.n21003 vdd.n21001 1.407
R53186 vdd.n18903 vdd.n18902 1.407
R53187 vdd.n18885 vdd.n18884 1.407
R53188 vdd.t346 vdd.n18849 1.407
R53189 vdd.n18644 vdd.n18643 1.407
R53190 vdd.n18626 vdd.n18625 1.407
R53191 vdd.n18574 vdd.t247 1.407
R53192 vdd.n24964 vdd.n24963 1.393
R53193 vdd.n24542 vdd.n24541 1.393
R53194 vdd.n24891 vdd.n24890 1.375
R53195 vdd.n33863 vdd.n33780 1.356
R53196 vdd.n35612 vdd.n35357 1.356
R53197 vdd.n35026 vdd.n34773 1.356
R53198 vdd.n5775 vdd.n5520 1.356
R53199 vdd.n4605 vdd.n4347 1.356
R53200 vdd.n6358 vdd.n5848 1.356
R53201 vdd.n33863 vdd.n33852 1.355
R53202 vdd.n33863 vdd.n33789 1.355
R53203 vdd.n587 vdd.n306 1.355
R53204 vdd.n587 vdd.n319 1.354
R53205 vdd.n6358 vdd.n5859 1.354
R53206 vdd.n6358 vdd.n5923 1.354
R53207 vdd.n587 vdd.n380 1.354
R53208 vdd.n587 vdd.n388 1.353
R53209 vdd.n33863 vdd.n33860 1.353
R53210 vdd.n1173 vdd.n961 1.353
R53211 vdd.n35844 vdd.n35843 1.341
R53212 vdd.n36002 vdd.n36001 1.341
R53213 vdd.n36072 vdd.n36071 1.341
R53214 vdd.n36233 vdd.n36232 1.341
R53215 vdd.n36303 vdd.n36302 1.341
R53216 vdd.n36464 vdd.n36463 1.341
R53217 vdd.n36534 vdd.n36533 1.341
R53218 vdd.n36695 vdd.n36694 1.341
R53219 vdd.n36765 vdd.n36764 1.341
R53220 vdd.n36926 vdd.n36925 1.341
R53221 vdd.n3653 vdd.n3652 1.341
R53222 vdd.n33173 vdd.n33172 1.341
R53223 vdd.n33135 vdd.n33134 1.341
R53224 vdd.n2402 vdd.n2401 1.341
R53225 vdd.n37386 vdd.n37385 1.341
R53226 vdd.n32847 vdd.n32846 1.341
R53227 vdd.n38211 vdd.n38210 1.341
R53228 vdd.n38051 vdd.n38050 1.341
R53229 vdd.n37981 vdd.n37980 1.341
R53230 vdd.n37820 vdd.n37819 1.341
R53231 vdd.n37750 vdd.n37749 1.341
R53232 vdd.n28192 vdd.n28191 1.341
R53233 vdd.n28262 vdd.n28261 1.341
R53234 vdd.n28423 vdd.n28422 1.341
R53235 vdd.n28493 vdd.n28492 1.341
R53236 vdd.n28654 vdd.n28653 1.341
R53237 vdd.n28724 vdd.n28723 1.341
R53238 vdd.n26210 vdd.n26206 1.341
R53239 vdd.n31755 vdd.n31751 1.341
R53240 vdd.n27837 vdd.n27836 1.341
R53241 vdd.n27913 vdd.n27912 1.341
R53242 vdd.n31488 vdd.n31484 1.341
R53243 vdd.n30220 vdd.n30219 1.341
R53244 vdd.n30503 vdd.n30502 1.341
R53245 bandgapmd_0.vdd vdd.n25256 1.325
R53246 vdd.n24882 vdd.n24881 1.313
R53247 vdd.n10466 vdd.n10465 1.29
R53248 vdd.n10430 vdd.n10429 1.29
R53249 vdd.n15286 vdd.n15285 1.29
R53250 vdd.n15337 vdd.n15336 1.29
R53251 vdd.n9319 vdd.n9317 1.283
R53252 vdd.n9383 vdd.n9368 1.283
R53253 vdd.t360 vdd.n9414 1.283
R53254 vdd.n12955 vdd.n9475 1.283
R53255 vdd.n9554 vdd.n9525 1.283
R53256 ldomc_0.otaldom_0.pmosrm_0.vdd vdd.n9610 1.283
R53257 vdd.n9679 vdd.n9678 1.283
R53258 vdd.n9743 vdd.n9728 1.283
R53259 vdd.n12747 vdd.n9835 1.283
R53260 vdd.n9914 vdd.n9886 1.283
R53261 vdd.n10039 vdd.n10038 1.283
R53262 vdd.n10188 vdd.n10139 1.283
R53263 vdd.n10577 vdd.n10564 1.283
R53264 vdd.n12471 vdd.n12470 1.283
R53265 vdd.n10688 vdd.t314 1.283
R53266 vdd.n12394 vdd.n10719 1.283
R53267 vdd.n12370 vdd.n10764 1.283
R53268 vdd.n12293 vdd.n12292 1.283
R53269 vdd.n12271 vdd.n10922 1.283
R53270 vdd.n12193 vdd.n12192 1.283
R53271 vdd.n12173 vdd.n11106 1.283
R53272 vdd.n11259 vdd.n11258 1.283
R53273 vdd.n12064 vdd.n11274 1.283
R53274 vdd.n11987 vdd.n11986 1.283
R53275 vdd.n11965 vdd.n11431 1.283
R53276 vdd.n15508 vdd.n15507 1.283
R53277 vdd.n15574 vdd.n15573 1.283
R53278 vdd.t28 vdd.n15228 1.283
R53279 vdd.n15764 vdd.n15763 1.283
R53280 vdd.n15830 vdd.n15829 1.283
R53281 vdd.n15199 bandgapmd_0.otam_1.pmosrm_0.vdd 1.283
R53282 vdd.n16020 vdd.n16019 1.283
R53283 vdd.n16086 vdd.n16085 1.283
R53284 vdd.n16276 vdd.n16275 1.283
R53285 vdd.n16342 vdd.n16341 1.283
R53286 vdd.n16532 vdd.n16531 1.283
R53287 vdd.n16550 vdd.n16549 1.283
R53288 vdd.n16947 vdd.n16946 1.283
R53289 vdd.n17007 vdd.n17006 1.283
R53290 vdd.n17123 vdd.t257 1.283
R53291 vdd.n17219 vdd.n17218 1.283
R53292 vdd.n17279 vdd.n17278 1.283
R53293 vdd.n17491 vdd.n17490 1.283
R53294 vdd.n17551 vdd.n17550 1.283
R53295 vdd.n17749 vdd.n17748 1.283
R53296 vdd.n17809 vdd.n17808 1.283
R53297 vdd.n18020 vdd.n18019 1.283
R53298 vdd.n18080 vdd.n18079 1.283
R53299 vdd.n18287 vdd.n18286 1.283
R53300 vdd.n18327 vdd.n18326 1.283
R53301 vdd.n13219 vdd.n13218 1.279
R53302 vdd.n28118 vdd.n28117 1.249
R53303 vdd.n11833 vdd.n11814 1.233
R53304 vdd.n21924 vdd.n21905 1.233
R53305 vdd.n11734 vdd.n11733 1.233
R53306 vdd.n21810 vdd.n21808 1.233
R53307 vdd.n25158 vdd.n25157 1.226
R53308 vdd.n24756 vdd.n24755 1.226
R53309 vdd.n13316 vdd.n9132 1.223
R53310 vdd.n13348 vdd.n9093 1.223
R53311 vdd.n13391 vdd.n13390 1.223
R53312 vdd.n13511 vdd.n8949 1.223
R53313 vdd.n8920 vdd.t136 1.223
R53314 vdd.n13608 vdd.n8910 1.223
R53315 vdd.n13640 vdd.n8873 1.223
R53316 vdd.n13683 vdd.n13682 1.223
R53317 vdd.n13810 vdd.n13809 1.223
R53318 vdd.n13889 vdd.n8693 1.223
R53319 vdd.n13905 vdd.n8677 1.223
R53320 vdd.n8601 vdd.n8594 1.223
R53321 vdd.n14097 vdd.n14096 1.223
R53322 vdd.n14178 vdd.n8470 1.223
R53323 vdd.n14195 vdd.n8453 1.223
R53324 vdd.n14207 vdd.t130 1.223
R53325 vdd.n8379 vdd.n8372 1.223
R53326 vdd.n14394 vdd.n8297 1.223
R53327 vdd.n14468 vdd.n8234 1.223
R53328 vdd.n14500 vdd.n8215 1.223
R53329 vdd.n27233 vdd.n27232 1.215
R53330 vdd.n31514 vdd.n31504 1.214
R53331 vdd.n32160 vdd.n32158 1.214
R53332 vdd.n32158 vdd.n32151 1.214
R53333 vdd.n31668 vdd.n31664 1.214
R53334 vdd.n32449 vdd.n32439 1.214
R53335 vdd.n32451 vdd.n32449 1.214
R53336 vdd.n10663 vdd.n10657 1.212
R53337 vdd.n10691 vdd.n10679 1.212
R53338 vdd.n10846 vdd.n10843 1.212
R53339 vdd.n10859 vdd.n10856 1.212
R53340 vdd.n11005 vdd.n11002 1.212
R53341 vdd.n12233 vdd.n11014 1.212
R53342 vdd.n12135 vdd.n11177 1.212
R53343 vdd.n11200 vdd.n11183 1.212
R53344 vdd.n11355 vdd.n11352 1.212
R53345 vdd.n11368 vdd.n11365 1.212
R53346 vdd.n10386 vdd.n10337 1.212
R53347 vdd.n10378 vdd.n10343 1.212
R53348 vdd.n9438 vdd.n9433 1.212
R53349 vdd.n12988 vdd.n9417 1.212
R53350 vdd.n12890 vdd.n9607 1.212
R53351 vdd.n12882 vdd.n9613 1.212
R53352 vdd.n9797 vdd.n9793 1.212
R53353 vdd.n12780 vdd.n9778 1.212
R53354 vdd.n12682 vdd.n9967 1.212
R53355 vdd.n12674 vdd.n9973 1.212
R53356 vdd.n10483 vdd.n10121 1.212
R53357 vdd.n17098 vdd.n17097 1.212
R53358 vdd.n17115 vdd.n17114 1.212
R53359 vdd.n17370 vdd.n17369 1.212
R53360 vdd.n17387 vdd.n17386 1.212
R53361 vdd.n17628 vdd.n17627 1.212
R53362 vdd.n17645 vdd.n17644 1.212
R53363 vdd.n17899 vdd.n17898 1.212
R53364 vdd.n17916 vdd.n17915 1.212
R53365 vdd.n18171 vdd.n18170 1.212
R53366 vdd.n18188 vdd.n18187 1.212
R53367 vdd.n15253 vdd.n15249 1.212
R53368 vdd.n15242 vdd.n15238 1.212
R53369 vdd.n15231 vdd.n15224 1.212
R53370 vdd.n15217 vdd.n15210 1.212
R53371 vdd.n15203 vdd.n15184 1.212
R53372 vdd.n15193 vdd.n15189 1.212
R53373 vdd.n15175 vdd.n15168 1.212
R53374 vdd.n15161 vdd.n15154 1.212
R53375 vdd.n15147 vdd.n15140 1.212
R53376 vdd.n15133 vdd.n15126 1.212
R53377 vdd.n16655 vdd.n16654 1.212
R53378 vdd.n12569 vdd.n10269 1.185
R53379 vdd.n12584 vdd.n10123 1.185
R53380 vdd.n12599 vdd.n12598 1.185
R53381 vdd.n10401 vdd.n10329 1.185
R53382 vdd.n10401 vdd.n10330 1.185
R53383 vdd.n10366 vdd.n10365 1.185
R53384 vdd.n10365 vdd.n10359 1.185
R53385 vdd.n13005 vdd.n9403 1.185
R53386 vdd.n13005 vdd.n13004 1.185
R53387 vdd.n12970 vdd.n9452 1.185
R53388 vdd.n12970 vdd.n12969 1.185
R53389 vdd.n9582 vdd.n9577 1.185
R53390 vdd.n9598 vdd.n9577 1.185
R53391 vdd.n9652 vdd.n9651 1.185
R53392 vdd.n9653 vdd.n9652 1.185
R53393 vdd.n12797 vdd.n9763 1.185
R53394 vdd.n12797 vdd.n12796 1.185
R53395 vdd.n12762 vdd.n9811 1.185
R53396 vdd.n12762 vdd.n12761 1.185
R53397 vdd.n9942 vdd.n9936 1.185
R53398 vdd.n9958 vdd.n9936 1.185
R53399 vdd.n10012 vdd.n10011 1.185
R53400 vdd.n10013 vdd.n10012 1.185
R53401 vdd.n10545 vdd.n10544 1.185
R53402 vdd.n12497 vdd.n10566 1.185
R53403 vdd.n12463 vdd.n10611 1.185
R53404 vdd.n12451 vdd.n10626 1.185
R53405 vdd.n12411 vdd.n10698 1.185
R53406 vdd.n10743 vdd.n10723 1.185
R53407 vdd.n10801 vdd.n10800 1.185
R53408 vdd.n10812 vdd.n10811 1.185
R53409 vdd.n10888 vdd.n10873 1.185
R53410 vdd.n12296 vdd.n12295 1.185
R53411 vdd.n10976 vdd.n10970 1.185
R53412 vdd.n12255 vdd.n10992 1.185
R53413 vdd.n11048 vdd.n11040 1.185
R53414 vdd.n12195 vdd.n11061 1.185
R53415 vdd.n12159 vdd.n12158 1.185
R53416 vdd.n11166 vdd.n11152 1.185
R53417 vdd.n12113 vdd.n12112 1.185
R53418 vdd.n11256 vdd.n11250 1.185
R53419 vdd.n11310 vdd.n11309 1.185
R53420 vdd.n11321 vdd.n11320 1.185
R53421 vdd.n11397 vdd.n11382 1.185
R53422 vdd.n11990 vdd.n11989 1.185
R53423 vdd.n11522 vdd.n11459 1.185
R53424 vdd.n11948 vdd.n11547 1.185
R53425 vdd.n15118 vdd.n15069 1.185
R53426 vdd.n15398 vdd.n15397 1.185
R53427 vdd.n15397 vdd.n15390 1.185
R53428 vdd.n15443 vdd.n15436 1.185
R53429 vdd.n15445 vdd.n15443 1.185
R53430 vdd.n15646 vdd.n15645 1.185
R53431 vdd.n15645 vdd.n15635 1.185
R53432 vdd.n15699 vdd.n15689 1.185
R53433 vdd.n15701 vdd.n15699 1.185
R53434 vdd.n15902 vdd.n15901 1.185
R53435 vdd.n15901 vdd.n15891 1.185
R53436 vdd.n15955 vdd.n15945 1.185
R53437 vdd.n15957 vdd.n15955 1.185
R53438 vdd.n16158 vdd.n16157 1.185
R53439 vdd.n16157 vdd.n16147 1.185
R53440 vdd.n16211 vdd.n16201 1.185
R53441 vdd.n16213 vdd.n16211 1.185
R53442 vdd.n16414 vdd.n16413 1.185
R53443 vdd.n16413 vdd.n16403 1.185
R53444 vdd.n16467 vdd.n16457 1.185
R53445 vdd.n16469 vdd.n16467 1.185
R53446 vdd.n16876 vdd.n16875 1.185
R53447 vdd.n16950 vdd.n16949 1.185
R53448 vdd.n17027 vdd.n17025 1.185
R53449 vdd.n17064 vdd.n17063 1.185
R53450 vdd.n17148 vdd.n17147 1.185
R53451 vdd.n17222 vdd.n17221 1.185
R53452 vdd.n17299 vdd.n17297 1.185
R53453 vdd.n17336 vdd.n17335 1.185
R53454 vdd.n17420 vdd.n17419 1.185
R53455 vdd.n17494 vdd.n17493 1.185
R53456 vdd.n17571 vdd.n17569 1.185
R53457 vdd.n16821 vdd.n16820 1.185
R53458 vdd.n17678 vdd.n17677 1.185
R53459 vdd.n17752 vdd.n17751 1.185
R53460 vdd.n17829 vdd.n17827 1.185
R53461 vdd.n17866 vdd.n17865 1.185
R53462 vdd.n17949 vdd.n17948 1.185
R53463 vdd.n18023 vdd.n18022 1.185
R53464 vdd.n18100 vdd.n18098 1.185
R53465 vdd.n18137 vdd.n18136 1.185
R53466 vdd.n18221 vdd.n18220 1.185
R53467 vdd.n18290 vdd.n18289 1.185
R53468 vdd.n18346 vdd.n18338 1.185
R53469 vdd.n11782 vdd.n11781 1.179
R53470 vdd.n21874 vdd.n21873 1.179
R53471 vdd.n19267 vdd.n19266 1.172
R53472 vdd.n19255 vdd.n19254 1.172
R53473 vdd.n19211 vdd.n19210 1.172
R53474 vdd.n19199 vdd.n19198 1.172
R53475 vdd.n19853 vdd.n19852 1.172
R53476 vdd.n19865 vdd.n19864 1.172
R53477 vdd.n19921 vdd.n19920 1.172
R53478 vdd.n19933 vdd.n19932 1.172
R53479 vdd.n20400 vdd.n20397 1.172
R53480 vdd.n20380 vdd.n20379 1.172
R53481 vdd.n20346 vdd.t253 1.172
R53482 vdd.n20200 vdd.t267 1.172
R53483 vdd.n20164 vdd.n20161 1.172
R53484 vdd.n20144 vdd.n20143 1.172
R53485 vdd.n14685 vdd.n14684 1.169
R53486 vdd.n14714 vdd.n14713 1.169
R53487 vdd.n14731 vdd.t307 1.169
R53488 vdd.n14846 vdd.t292 1.169
R53489 vdd.n14859 vdd.n14858 1.169
R53490 vdd.n14906 vdd.n8021 1.169
R53491 vdd.n32128 vdd.n32127 1.166
R53492 vdd.n1819 vdd.n1818 1.161
R53493 vdd.n13139 vdd.n13138 1.161
R53494 vdd.n21689 vdd.n21688 1.161
R53495 vdd.n2510 vdd.n2508 1.16
R53496 vdd.n4657 vdd.n4656 1.156
R53497 vdd.n34011 vdd.n34010 1.153
R53498 vdd.n35174 vdd.n35173 1.153
R53499 vdd.n34599 vdd.n34598 1.153
R53500 vdd.n6311 vdd.n6310 1.153
R53501 vdd.n5346 vdd.n5345 1.153
R53502 vdd.n4177 vdd.n4176 1.153
R53503 vdd.n10240 vdd.n10236 1.147
R53504 vdd.n16668 vdd.n16667 1.147
R53505 vdd.n11900 vdd.n11793 1.143
R53506 vdd.n21991 vdd.n21884 1.143
R53507 vdd.n11772 vdd.n11771 1.141
R53508 vdd.n11876 vdd.n11804 1.141
R53509 vdd.n21865 vdd.n21864 1.141
R53510 vdd.n21967 vdd.n21895 1.141
R53511 vdd.n11906 vdd.n11905 1.141
R53512 vdd.n21997 vdd.n21996 1.141
R53513 vdd.n14975 ldomc_0.otaldom_0.pmosbm_0.vdd 1.136
R53514 vdd.n25257 vdd.n21747 1.133
R53515 vdd.n1813 vdd.n1812 1.13
R53516 vdd.n33777 vdd.n33776 1.129
R53517 vdd.n33707 vdd.n33706 1.129
R53518 vdd.n33694 vdd.n33693 1.129
R53519 vdd.n33480 vdd.n33479 1.129
R53520 vdd.n33359 vdd.n33358 1.129
R53521 vdd.n34229 vdd.n34228 1.129
R53522 vdd.n34080 vdd.n34079 1.129
R53523 vdd.n34336 vdd.n34335 1.129
R53524 vdd.n33869 vdd.n33867 1.129
R53525 vdd.n33897 vdd.n33896 1.129
R53526 vdd.n34349 vdd.n34348 1.129
R53527 vdd.n35120 vdd.n35118 1.129
R53528 vdd.n35091 vdd.n35090 1.129
R53529 vdd.n35367 vdd.n35366 1.129
R53530 vdd.n35602 vdd.n35601 1.129
R53531 vdd.n35239 vdd.n35238 1.129
R53532 vdd.n35350 vdd.n35349 1.129
R53533 vdd.n34766 vdd.n34765 1.129
R53534 vdd.n34652 vdd.n34651 1.129
R53535 vdd.n35014 vdd.n35013 1.129
R53536 vdd.n34533 vdd.n34531 1.129
R53537 vdd.n34504 vdd.n34503 1.129
R53538 vdd.n34777 vdd.n34776 1.129
R53539 vdd.n872 vdd.n871 1.129
R53540 vdd.n791 vdd.n790 1.129
R53541 vdd.n1160 vdd.n1159 1.129
R53542 vdd.n965 vdd.n964 1.129
R53543 vdd.n677 vdd.n676 1.129
R53544 vdd.n224 vdd.n223 1.129
R53545 vdd.n253 vdd.n252 1.129
R53546 vdd.n251 vdd.n250 1.129
R53547 vdd.n3 vdd.n2 1.129
R53548 vdd.n12 vdd.n11 1.129
R53549 vdd.n46 vdd.n45 1.129
R53550 vdd.n569 vdd.n568 1.129
R53551 vdd.n6143 vdd.n6141 1.129
R53552 vdd.n6171 vdd.n6170 1.129
R53553 vdd.n6055 vdd.n6054 1.129
R53554 vdd.n6037 vdd.n6036 1.129
R53555 vdd.n5782 vdd.n5781 1.129
R53556 vdd.n5856 vdd.n5855 1.129
R53557 vdd.n5513 vdd.n5512 1.129
R53558 vdd.n5399 vdd.n5398 1.129
R53559 vdd.n5761 vdd.n5760 1.129
R53560 vdd.n5280 vdd.n5278 1.129
R53561 vdd.n5251 vdd.n5250 1.129
R53562 vdd.n5524 vdd.n5523 1.129
R53563 vdd.n4701 vdd.n4700 1.129
R53564 vdd.n4793 vdd.n4791 1.129
R53565 vdd.n4979 vdd.n4978 1.129
R53566 vdd.n4955 vdd.n4954 1.129
R53567 vdd.n5080 vdd.n5079 1.129
R53568 vdd.n4822 vdd.n4821 1.129
R53569 vdd.n4824 vdd.n4823 1.129
R53570 vdd.n4804 vdd.n4803 1.129
R53571 vdd.n4340 vdd.n4339 1.129
R53572 vdd.n4229 vdd.n4228 1.129
R53573 vdd.n4591 vdd.n4590 1.129
R53574 vdd.n4110 vdd.n4108 1.129
R53575 vdd.n4081 vdd.n4080 1.129
R53576 vdd.n4351 vdd.n4350 1.129
R53577 vdd.n30284 vdd.n30283 1.129
R53578 vdd.n31517 vdd.n31516 1.129
R53579 vdd.n31535 vdd.n31534 1.129
R53580 vdd.n31560 vdd.n31559 1.129
R53581 vdd.n31557 vdd.n31556 1.129
R53582 vdd.n31037 vdd.n31036 1.129
R53583 vdd.n31040 vdd.n31039 1.129
R53584 vdd.n31264 vdd.n31263 1.129
R53585 vdd.n30540 vdd.n30539 1.129
R53586 vdd.n35892 vdd.n35891 1.129
R53587 vdd.n35941 vdd.n35940 1.129
R53588 vdd.n36123 vdd.n36122 1.129
R53589 vdd.n36172 vdd.n36171 1.129
R53590 vdd.n36354 vdd.n36353 1.129
R53591 vdd.n36403 vdd.n36402 1.129
R53592 vdd.n36585 vdd.n36584 1.129
R53593 vdd.n36634 vdd.n36633 1.129
R53594 vdd.n36816 vdd.n36815 1.129
R53595 vdd.n36865 vdd.n36864 1.129
R53596 vdd.n37051 vdd.n37050 1.129
R53597 vdd.n37090 vdd.n37089 1.129
R53598 vdd.n37224 vdd.n37223 1.129
R53599 vdd.n33052 vdd.n33051 1.129
R53600 vdd.n32922 vdd.n32921 1.129
R53601 vdd.n37463 vdd.n37462 1.129
R53602 vdd.n38145 vdd.n38144 1.129
R53603 vdd.n38102 vdd.n38101 1.129
R53604 vdd.n37920 vdd.n37919 1.129
R53605 vdd.n37871 vdd.n37870 1.129
R53606 vdd.n37689 vdd.n37688 1.129
R53607 vdd.n37640 vdd.n37639 1.129
R53608 vdd.n28313 vdd.n28312 1.129
R53609 vdd.n28362 vdd.n28361 1.129
R53610 vdd.n28544 vdd.n28543 1.129
R53611 vdd.n28593 vdd.n28592 1.129
R53612 vdd.n28775 vdd.n28774 1.129
R53613 vdd.n28158 vdd.n28157 1.129
R53614 vdd.n28132 vdd.n28131 1.129
R53615 vdd.n28816 vdd.n28815 1.129
R53616 vdd.n28124 vdd.n28123 1.129
R53617 vdd.n27747 vdd.n27746 1.129
R53618 vdd.n29032 vdd.n29031 1.129
R53619 vdd.n27821 vdd.n27820 1.129
R53620 vdd.n27814 vdd.n27811 1.129
R53621 vdd.n29865 vdd.n29864 1.129
R53622 vdd.n29945 vdd.n29944 1.129
R53623 vdd.n29845 vdd.n29844 1.129
R53624 vdd.n29844 vdd.n29843 1.129
R53625 vdd.n29831 vdd.n29830 1.129
R53626 vdd.n29812 vdd.n29811 1.129
R53627 vdd.n29766 vdd.n29765 1.129
R53628 vdd.n30205 vdd.n30204 1.129
R53629 vdd.n27356 vdd.n27355 1.129
R53630 vdd.n27653 vdd.n27652 1.129
R53631 vdd.n27300 vdd.n27299 1.129
R53632 vdd.n27462 vdd.n27461 1.129
R53633 vdd.n27277 vdd.n27276 1.129
R53634 vdd.n27554 vdd.n27553 1.129
R53635 vdd.n27587 vdd.n27585 1.129
R53636 vdd.n25808 vdd.n25807 1.129
R53637 vdd.n26075 vdd.n26074 1.129
R53638 vdd.n25752 vdd.n25751 1.129
R53639 vdd.n25908 vdd.n25907 1.129
R53640 vdd.n25723 vdd.n25722 1.129
R53641 vdd.n25991 vdd.n25990 1.129
R53642 vdd.n26003 vdd.n26001 1.129
R53643 vdd.n25445 vdd.n25444 1.129
R53644 vdd.n25487 vdd.n25486 1.129
R53645 vdd.n25578 vdd.n25577 1.129
R53646 vdd.n1754 vdd.n1753 1.129
R53647 vdd.n1721 vdd.n1720 1.129
R53648 vdd.n1579 vdd.n1578 1.129
R53649 vdd.n1540 vdd.n1539 1.129
R53650 vdd.n1398 vdd.n1397 1.129
R53651 vdd.n1359 vdd.n1358 1.129
R53652 vdd.n26825 vdd.n26824 1.129
R53653 vdd.n26864 vdd.n26863 1.129
R53654 vdd.n27006 vdd.n27005 1.129
R53655 vdd.n27045 vdd.n27044 1.129
R53656 vdd.n27187 vdd.n27186 1.129
R53657 vdd.n26733 vdd.n26732 1.129
R53658 vdd.n1909 vdd.n1908 1.129
R53659 vdd.n1908 vdd.n1901 1.129
R53660 vdd.n1910 vdd.n1898 1.129
R53661 vdd.n1202 vdd.n1201 1.129
R53662 vdd.n1184 vdd.n1183 1.129
R53663 vdd.n1186 vdd.n1182 1.129
R53664 vdd.n2671 vdd.n2670 1.129
R53665 vdd.n2641 vdd.n2640 1.129
R53666 vdd.n2640 vdd.n2639 1.129
R53667 vdd.n2445 vdd.n2443 1.129
R53668 vdd.n2423 vdd.n2413 1.129
R53669 vdd.n2043 vdd.n2042 1.129
R53670 vdd.n2044 vdd.n2043 1.129
R53671 vdd.n2113 vdd.n2112 1.129
R53672 vdd.n2111 vdd.n2110 1.129
R53673 vdd.n2151 vdd.n2150 1.129
R53674 vdd.n2197 vdd.n2189 1.129
R53675 vdd.n3923 vdd.n3922 1.129
R53676 vdd.n2017 vdd.n2016 1.129
R53677 vdd.n2018 vdd.n2017 1.129
R53678 vdd.n3742 vdd.n3741 1.129
R53679 vdd.n3740 vdd.n3739 1.129
R53680 vdd.n2702 vdd.n2701 1.129
R53681 vdd.n2699 vdd.n2698 1.129
R53682 vdd.n2059 vdd.n2057 1.129
R53683 vdd.n2778 vdd.n2777 1.129
R53684 vdd.n2817 vdd.n2816 1.129
R53685 vdd.n2959 vdd.n2958 1.129
R53686 vdd.n2998 vdd.n2997 1.129
R53687 vdd.n3140 vdd.n3139 1.129
R53688 vdd.n3179 vdd.n3178 1.129
R53689 vdd.n3321 vdd.n3320 1.129
R53690 vdd.n3360 vdd.n3359 1.129
R53691 vdd.n3502 vdd.n3501 1.129
R53692 vdd.n3541 vdd.n3540 1.129
R53693 vdd.n2057 vdd.n2049 1.129
R53694 vdd.n31723 vdd.n31722 1.129
R53695 vdd.n31724 vdd.n31723 1.129
R53696 vdd.n31726 vdd.n31724 1.129
R53697 vdd.n31701 vdd.n31700 1.129
R53698 vdd.n31704 vdd.n31703 1.129
R53699 vdd.n31927 vdd.n31926 1.129
R53700 vdd.n13179 vdd.n9206 1.129
R53701 vdd.n13209 vdd.n13208 1.129
R53702 vdd.n13250 vdd.n13249 1.129
R53703 vdd.n13269 vdd.n13268 1.129
R53704 vdd.n13474 vdd.n8986 1.129
R53705 vdd.n13561 vdd.n13560 1.129
R53706 vdd.n13780 vdd.n8771 1.129
R53707 vdd.n13843 vdd.n13842 1.129
R53708 vdd.n14072 vdd.n8554 1.129
R53709 vdd.n14132 vdd.n14131 1.129
R53710 vdd.n14358 vdd.n14357 1.129
R53711 vdd.n8338 vdd.n8337 1.129
R53712 vdd.n14426 vdd.n8278 1.129
R53713 vdd.n8283 vdd.n8282 1.129
R53714 vdd.n8090 vdd.n8089 1.129
R53715 vdd.n8089 vdd.n8069 1.129
R53716 vdd.n14804 vdd.n8061 1.129
R53717 vdd.n14805 vdd.n14804 1.129
R53718 vdd.n9255 vdd.n9249 1.129
R53719 vdd.n13135 vdd.n9261 1.129
R53720 vdd.n9087 vdd.n9086 1.129
R53721 vdd.n9080 vdd.n9079 1.129
R53722 vdd.n13434 vdd.n9025 1.129
R53723 vdd.n9030 vdd.n9029 1.129
R53724 vdd.n8867 vdd.n8866 1.129
R53725 vdd.n8860 vdd.n8859 1.129
R53726 vdd.n13726 vdd.n8805 1.129
R53727 vdd.n8810 vdd.n8809 1.129
R53728 vdd.n13945 vdd.n8634 1.129
R53729 vdd.n13954 vdd.n8635 1.129
R53730 vdd.n13997 vdd.n8586 1.129
R53731 vdd.n14019 vdd.n8583 1.129
R53732 vdd.n14235 vdd.n8412 1.129
R53733 vdd.n14244 vdd.n8413 1.129
R53734 vdd.n14288 vdd.n8366 1.129
R53735 vdd.n14308 vdd.n8364 1.129
R53736 vdd.n14551 vdd.n14538 1.129
R53737 vdd.n14544 vdd.n14542 1.129
R53738 vdd.n24292 vdd.n24285 1.129
R53739 vdd.n24293 vdd.n24292 1.129
R53740 vdd.n24187 vdd.n24180 1.129
R53741 vdd.n23993 vdd.n23986 1.129
R53742 vdd.n23955 vdd.n23948 1.129
R53743 vdd.n23761 vdd.n23754 1.129
R53744 vdd.n23723 vdd.n23716 1.129
R53745 vdd.n23073 vdd.n23066 1.129
R53746 vdd.n23267 vdd.n23260 1.129
R53747 vdd.n23305 vdd.n23298 1.129
R53748 vdd.n23499 vdd.n23492 1.129
R53749 vdd.n23537 vdd.n23530 1.129
R53750 vdd.n22494 vdd.n22487 1.129
R53751 vdd.n22688 vdd.n22681 1.129
R53752 vdd.n22726 vdd.n22719 1.129
R53753 vdd.n22920 vdd.n22913 1.129
R53754 vdd.n22958 vdd.n22951 1.129
R53755 vdd.n22464 vdd.n22457 1.129
R53756 vdd.n22465 vdd.n22464 1.129
R53757 vdd.n22320 vdd.n22313 1.129
R53758 vdd.n22321 vdd.n22320 1.129
R53759 vdd.n19392 vdd.n19391 1.129
R53760 vdd.n19441 vdd.n19440 1.129
R53761 vdd.n19598 vdd.n19597 1.129
R53762 vdd.n19641 vdd.n19640 1.129
R53763 vdd.n19800 vdd.n19799 1.129
R53764 vdd.n19160 vdd.n19159 1.129
R53765 vdd.n20849 vdd.n20848 1.129
R53766 vdd.n20806 vdd.n20805 1.129
R53767 vdd.n20650 vdd.n20649 1.129
R53768 vdd.n20601 vdd.n20600 1.129
R53769 vdd.n21680 vdd.n21679 1.129
R53770 vdd.n21407 vdd.n21406 1.129
R53771 vdd.n21358 vdd.n21357 1.129
R53772 vdd.n21148 vdd.n21147 1.129
R53773 vdd.n21099 vdd.n21098 1.129
R53774 vdd.n19041 vdd.n19040 1.129
R53775 vdd.n18992 vdd.n18991 1.129
R53776 vdd.n18782 vdd.n18781 1.129
R53777 vdd.n18733 vdd.n18732 1.129
R53778 vdd.n18523 vdd.n18522 1.129
R53779 vdd.n20284 vdd.n20275 1.129
R53780 vdd.n20266 vdd.n20257 1.129
R53781 vdd.n24829 vdd.n24824 1.129
R53782 vdd.n25247 vdd.n25242 1.129
R53783 vdd.n11489 vdd.n11488 1.125
R53784 vdd.n18310 vdd.n16809 1.125
R53785 vdd.n35882 vdd.n35881 1.117
R53786 vdd.n35959 vdd.n35958 1.117
R53787 vdd.n36113 vdd.n36112 1.117
R53788 vdd.n36190 vdd.n36189 1.117
R53789 vdd.n36344 vdd.n36343 1.117
R53790 vdd.n36421 vdd.n36420 1.117
R53791 vdd.n36575 vdd.n36574 1.117
R53792 vdd.n36652 vdd.n36651 1.117
R53793 vdd.n36806 vdd.n36805 1.117
R53794 vdd.n36883 vdd.n36882 1.117
R53795 vdd.n2719 vdd.n2718 1.117
R53796 vdd.n33217 vdd.n33216 1.117
R53797 vdd.n2176 vdd.n2175 1.117
R53798 vdd.n37276 vdd.n37275 1.117
R53799 vdd.n37417 vdd.n37416 1.117
R53800 vdd.n37479 vdd.n37478 1.117
R53801 vdd.n38165 vdd.n38164 1.117
R53802 vdd.n38092 vdd.n38091 1.117
R53803 vdd.n37938 vdd.n37937 1.117
R53804 vdd.n37861 vdd.n37860 1.117
R53805 vdd.n37707 vdd.n37706 1.117
R53806 vdd.n37630 vdd.n37629 1.117
R53807 vdd.n28303 vdd.n28302 1.117
R53808 vdd.n28380 vdd.n28379 1.117
R53809 vdd.n28534 vdd.n28533 1.117
R53810 vdd.n28611 vdd.n28610 1.117
R53811 vdd.n28765 vdd.n28764 1.117
R53812 vdd.n28172 vdd.n28171 1.117
R53813 vdd.n28987 vdd.n28986 1.117
R53814 vdd.n27791 vdd.n27790 1.117
R53815 vdd.n31568 vdd.n31567 1.117
R53816 vdd.n29816 vdd.n29815 1.117
R53817 vdd.n30271 vdd.n30270 1.117
R53818 vdd.n31257 vdd.n31256 1.117
R53819 vdd.n1178 vdd.n1177 1.108
R53820 vdd.n25257 vdd.n22004 1.104
R53821 vdd.n1236 vdd.n1235 1.101
R53822 vdd.n25146 vdd.n25145 1.081
R53823 vdd.n24768 vdd.n24767 1.081
R53824 vdd.n25669 vdd.n25397 1.075
R53825 vdd.n25439 vdd.n25438 1.07
R53826 vdd.n2422 vdd.n2421 1.068
R53827 vdd.n32405 vdd.n32395 1.066
R53828 vdd.n31462 vdd.n31452 1.066
R53829 vdd.n31599 vdd.n31595 1.066
R53830 vdd.n26312 vdd.n26302 1.066
R53831 vdd.n10247 vdd.n10246 1.066
R53832 vdd.n10246 vdd.n10231 1.066
R53833 vdd.n16669 vdd.n16649 1.066
R53834 vdd.n16669 vdd.n16646 1.066
R53835 vdd.n32093 vdd.n32092 1.059
R53836 vdd.n27226 vdd.n27219 1.05
R53837 vdd.n3820 vdd.n3819 1.043
R53838 vdd.n5189 vdd.n4951 1.038
R53839 vdd.n1173 vdd.n1172 1.038
R53840 vdd.n587 vdd.n210 1.038
R53841 vdd.n31600 vdd.n31594 1.038
R53842 vdd.n34443 vdd.n34232 1.036
R53843 vdd.n25258 vdd.n25257 1.027
R53844 vdd.n25465 vdd.n25464 1.01
R53845 vdd.n32387 vdd.n32385 1.009
R53846 vdd.n10540 vdd.n10520 1.009
R53847 vdd.n16873 vdd.n16872 1.009
R53848 vdd.n28832 vdd.n28831 1.005
R53849 vdd.n28102 vdd.n28101 1.005
R53850 vdd.n3672 vdd.n3664 1.001
R53851 vdd.n28092 vdd.n28089 0.985
R53852 vdd.n2521 vdd.n2520 0.985
R53853 vdd.n35693 vdd.n35692 0.981
R53854 vdd.n35699 vdd.n35698 0.981
R53855 vdd.n32485 vdd.n32481 0.978
R53856 vdd.n25416 vdd.n25415 0.976
R53857 vdd.n27225 vdd.n27224 0.975
R53858 vdd.n10394 vdd.n10393 0.968
R53859 vdd.n25422 vdd.n25419 0.964
R53860 vdd.n10370 vdd.n10357 0.962
R53861 vdd.n9435 vdd.n9434 0.962
R53862 vdd.n12984 vdd.n9421 0.962
R53863 vdd.n12919 vdd.t366 0.962
R53864 vdd.n12898 vdd.n9571 0.962
R53865 vdd.n9646 vdd.n9630 0.962
R53866 vdd.t304 vdd.n12851 0.962
R53867 vdd.n9794 vdd.n9769 0.962
R53868 vdd.n12690 vdd.n9930 0.962
R53869 vdd.n10006 vdd.n9990 0.962
R53870 vdd.n10239 vdd.n10103 0.962
R53871 vdd.n10487 vdd.n10480 0.962
R53872 vdd.n12521 vdd.n10518 0.962
R53873 vdd.n12443 vdd.n12442 0.962
R53874 vdd.n12425 vdd.n10672 0.962
R53875 vdd.n12413 vdd.t357 0.962
R53876 vdd.n12342 vdd.n12341 0.962
R53877 vdd.n12323 vdd.n10862 0.962
R53878 vdd.n11003 vdd.n10994 0.962
R53879 vdd.n12223 vdd.n12222 0.962
R53880 vdd.n12144 vdd.n11145 0.962
R53881 vdd.n11211 vdd.n11210 0.962
R53882 vdd.n12036 vdd.n12035 0.962
R53883 vdd.n12017 vdd.n11371 0.962
R53884 vdd.n11933 vdd.n11549 0.962
R53885 vdd.n15427 vdd.n15426 0.962
R53886 vdd.n15660 vdd.n15659 0.962
R53887 vdd.n15680 vdd.n15679 0.962
R53888 vdd.n15848 vdd.t34 0.962
R53889 vdd.n15916 vdd.n15915 0.962
R53890 vdd.n15936 vdd.n15935 0.962
R53891 vdd.n16007 vdd.t261 0.962
R53892 vdd.n16172 vdd.n16171 0.962
R53893 vdd.n16428 vdd.n16427 0.962
R53894 vdd.n16448 vdd.n16447 0.962
R53895 vdd.n16643 vdd.n16642 0.962
R53896 vdd.n15079 vdd.n15075 0.962
R53897 vdd.n16868 vdd.n16865 0.962
R53898 vdd.n17086 vdd.n17083 0.962
R53899 vdd.n17138 vdd.n17135 0.962
R53900 vdd.n17151 vdd.t8 0.962
R53901 vdd.n17358 vdd.n17355 0.962
R53902 vdd.n17410 vdd.n17407 0.962
R53903 vdd.n17616 vdd.n17613 0.962
R53904 vdd.n17668 vdd.n17665 0.962
R53905 vdd.n17887 vdd.n17884 0.962
R53906 vdd.n17939 vdd.n17936 0.962
R53907 vdd.n18159 vdd.n18156 0.962
R53908 vdd.n18211 vdd.n18208 0.962
R53909 vdd.n15011 vdd.n15010 0.962
R53910 vdd.n15410 vdd.n15409 0.96
R53911 vdd.n13133 vdd.n13132 0.959
R53912 vdd.n12598 vdd.n12597 0.948
R53913 vdd.n10463 vdd.n10281 0.948
R53914 vdd.n10458 vdd.n10282 0.948
R53915 vdd.n10437 vdd.n10300 0.948
R53916 vdd.n10427 vdd.n10305 0.948
R53917 vdd.n9313 vdd.n9312 0.948
R53918 vdd.n9337 vdd.n9314 0.948
R53919 vdd.n9374 vdd.n9373 0.948
R53920 vdd.n9381 vdd.n9370 0.948
R53921 vdd.n12953 vdd.n12952 0.948
R53922 vdd.n9513 vdd.n9479 0.948
R53923 vdd.n9545 vdd.n9528 0.948
R53924 vdd.n9549 vdd.n9529 0.948
R53925 vdd.n9674 vdd.n9673 0.948
R53926 vdd.n9697 vdd.n9675 0.948
R53927 vdd.n9734 vdd.n9733 0.948
R53928 vdd.n9741 vdd.n9730 0.948
R53929 vdd.n12745 vdd.n12744 0.948
R53930 vdd.n9873 vdd.n9839 0.948
R53931 vdd.n9905 vdd.n9889 0.948
R53932 vdd.n9909 vdd.n9890 0.948
R53933 vdd.n10034 vdd.n10033 0.948
R53934 vdd.n10150 vdd.n10035 0.948
R53935 vdd.n10171 vdd.n10170 0.948
R53936 vdd.n10183 vdd.n10080 0.948
R53937 vdd.n10186 vdd.n10185 0.948
R53938 vdd.n10542 vdd.n10521 0.948
R53939 vdd.n10575 vdd.n10566 0.948
R53940 vdd.n12468 vdd.n10603 0.948
R53941 vdd.n12438 vdd.n10658 0.948
R53942 vdd.n12421 vdd.n10676 0.948
R53943 vdd.n12392 vdd.n10723 0.948
R53944 vdd.n10789 vdd.n10788 0.948
R53945 vdd.n10837 vdd.n10833 0.948
R53946 vdd.n10878 vdd.n10876 0.948
R53947 vdd.n12295 vdd.n10901 0.948
R53948 vdd.n12274 vdd.n12273 0.948
R53949 vdd.n11022 vdd.n11000 0.948
R53950 vdd.n12219 vdd.n12218 0.948
R53951 vdd.n12195 vdd.n11084 0.948
R53952 vdd.n12171 vdd.n12170 0.948
R53953 vdd.n12137 vdd.n11150 0.948
R53954 vdd.n11215 vdd.n11214 0.948
R53955 vdd.n11256 vdd.n11247 0.948
R53956 vdd.n11298 vdd.n11297 0.948
R53957 vdd.n11346 vdd.n11342 0.948
R53958 vdd.n11387 vdd.n11385 0.948
R53959 vdd.n11989 vdd.n11410 0.948
R53960 vdd.n11968 vdd.n11967 0.948
R53961 vdd.n11504 vdd.n11458 0.948
R53962 vdd.n11518 vdd.n11517 0.948
R53963 vdd.n11517 vdd.n11516 0.948
R53964 vdd.n11531 vdd.n11530 0.948
R53965 vdd.n11531 vdd.n11454 0.948
R53966 vdd.n11955 vdd.n11954 0.948
R53967 vdd.n11938 vdd.n11552 0.948
R53968 vdd.n11597 vdd.n11586 0.948
R53969 vdd.n15282 vdd.n15281 0.948
R53970 vdd.n15291 vdd.n15290 0.948
R53971 vdd.n15341 vdd.n15331 0.948
R53972 vdd.n15333 vdd.n15332 0.948
R53973 vdd.n15504 vdd.n15503 0.948
R53974 vdd.n15516 vdd.n15515 0.948
R53975 vdd.n15578 vdd.n15565 0.948
R53976 vdd.n15567 vdd.n15566 0.948
R53977 vdd.n15760 vdd.n15759 0.948
R53978 vdd.n15772 vdd.n15771 0.948
R53979 vdd.n15834 vdd.n15821 0.948
R53980 vdd.n15823 vdd.n15822 0.948
R53981 vdd.n16016 vdd.n16015 0.948
R53982 vdd.n16028 vdd.n16027 0.948
R53983 vdd.n16090 vdd.n16077 0.948
R53984 vdd.n16079 vdd.n16078 0.948
R53985 vdd.n16272 vdd.n16271 0.948
R53986 vdd.n16284 vdd.n16283 0.948
R53987 vdd.n16346 vdd.n16333 0.948
R53988 vdd.n16335 vdd.n16334 0.948
R53989 vdd.n16528 vdd.n16527 0.948
R53990 vdd.n16540 vdd.n16539 0.948
R53991 vdd.n16711 vdd.n16710 0.948
R53992 vdd.n16715 vdd.n16712 0.948
R53993 vdd.n16886 vdd.n16874 0.948
R53994 vdd.n16949 vdd.n16940 0.948
R53995 vdd.n17009 vdd.n17000 0.948
R53996 vdd.n17091 vdd.n17090 0.948
R53997 vdd.n17158 vdd.n17146 0.948
R53998 vdd.n17221 vdd.n17212 0.948
R53999 vdd.n17281 vdd.n17272 0.948
R54000 vdd.n17363 vdd.n17362 0.948
R54001 vdd.n17430 vdd.n17418 0.948
R54002 vdd.n17493 vdd.n17484 0.948
R54003 vdd.n17553 vdd.n17544 0.948
R54004 vdd.n17621 vdd.n17620 0.948
R54005 vdd.n17688 vdd.n17676 0.948
R54006 vdd.n17751 vdd.n17742 0.948
R54007 vdd.n17811 vdd.n17802 0.948
R54008 vdd.n17892 vdd.n17891 0.948
R54009 vdd.n17959 vdd.n17947 0.948
R54010 vdd.n18022 vdd.n18013 0.948
R54011 vdd.n18082 vdd.n18073 0.948
R54012 vdd.n18164 vdd.n18163 0.948
R54013 vdd.n18230 vdd.n18219 0.948
R54014 vdd.n18289 vdd.n18281 0.948
R54015 vdd.n18329 vdd.n18320 0.948
R54016 vdd.n18347 vdd.n18337 0.948
R54017 vdd.n18354 vdd.n18353 0.948
R54018 vdd.n18355 vdd.n18354 0.948
R54019 vdd.n18368 vdd.n18360 0.948
R54020 vdd.n18368 vdd.n18367 0.948
R54021 vdd.n18381 vdd.n18380 0.948
R54022 vdd.n18402 vdd.n18400 0.948
R54023 vdd.n18413 vdd.n18412 0.948
R54024 vdd.n28826 vdd.n28825 0.942
R54025 vdd.n24622 vdd.n24619 0.942
R54026 vdd.n11747 vdd.n11746 0.938
R54027 vdd.n21829 vdd.n21828 0.938
R54028 vdd.n2685 vdd.n2684 0.937
R54029 vdd.n24780 vdd.n24779 0.932
R54030 vdd.n25133 vdd.n25132 0.932
R54031 vdd.n3671 vdd.n3670 0.93
R54032 vdd.n31617 vdd.n31616 0.924
R54033 vdd.n26705 vdd.n26704 0.924
R54034 vdd.n13257 vdd.t323 0.917
R54035 vdd.n13266 vdd.n13265 0.917
R54036 vdd.n13354 vdd.n9062 0.917
R54037 vdd.n13427 vdd.n13426 0.917
R54038 vdd.n13420 vdd.t334 0.917
R54039 vdd.t116 vdd.n13480 0.917
R54040 vdd.n13498 vdd.n8988 0.917
R54041 vdd.n13558 vdd.n13557 0.917
R54042 vdd.n13646 vdd.n8842 0.917
R54043 vdd.n13719 vdd.n13718 0.917
R54044 vdd.n13778 vdd.n8754 0.917
R54045 vdd.n13840 vdd.n13839 0.917
R54046 vdd.n13943 vdd.n8629 0.917
R54047 vdd.n14011 vdd.n8564 0.917
R54048 vdd.n8552 vdd.n8541 0.917
R54049 vdd.n8498 vdd.n8490 0.917
R54050 vdd.n14233 vdd.n8407 0.917
R54051 vdd.n14301 vdd.n8346 0.917
R54052 vdd.n14360 vdd.n8333 0.917
R54053 vdd.n14419 vdd.t332 0.917
R54054 vdd.n8287 vdd.n8286 0.917
R54055 vdd.n14530 vdd.n8187 0.917
R54056 vdd.n14549 vdd.n14548 0.917
R54057 vdd.n8173 vdd.n8145 0.917
R54058 vdd.n31611 vdd.n31610 0.911
R54059 vdd.n26693 vdd.n26692 0.911
R54060 vdd.n26302 vdd.n26301 0.91
R54061 vdd.n6358 vdd.n6137 0.898
R54062 vdd.n24843 vdd.n24842 0.897
R54063 vdd.n32737 vdd.n30013 0.894
R54064 vdd.n27660 vdd.n25355 0.894
R54065 vdd.n36016 vdd.n36015 0.894
R54066 vdd.n36058 vdd.n36057 0.894
R54067 vdd.n36247 vdd.n36246 0.894
R54068 vdd.n36289 vdd.n36288 0.894
R54069 vdd.n36478 vdd.n36477 0.894
R54070 vdd.n36520 vdd.n36519 0.894
R54071 vdd.n36709 vdd.n36708 0.894
R54072 vdd.n36751 vdd.n36750 0.894
R54073 vdd.n36940 vdd.n36939 0.894
R54074 vdd.n3643 vdd.n3642 0.894
R54075 vdd.n37148 vdd.n37147 0.894
R54076 vdd.n37176 vdd.n37175 0.894
R54077 vdd.n32989 vdd.n32988 0.894
R54078 vdd.n32975 vdd.n32974 0.894
R54079 vdd.n37523 vdd.n37522 0.894
R54080 vdd.n37569 vdd.n37568 0.894
R54081 vdd.n38037 vdd.n38036 0.894
R54082 vdd.n37995 vdd.n37994 0.894
R54083 vdd.n37806 vdd.n37805 0.894
R54084 vdd.n37764 vdd.n37763 0.894
R54085 vdd.n28206 vdd.n28205 0.894
R54086 vdd.n28248 vdd.n28247 0.894
R54087 vdd.n28437 vdd.n28436 0.894
R54088 vdd.n28479 vdd.n28478 0.894
R54089 vdd.n28668 vdd.n28667 0.894
R54090 vdd.n28710 vdd.n28709 0.894
R54091 vdd.n28113 vdd.n28112 0.894
R54092 vdd.n28087 vdd.n28086 0.894
R54093 vdd.n31629 vdd.n31625 0.894
R54094 vdd.n32067 vdd.n32063 0.894
R54095 vdd.n29721 vdd.n29720 0.894
R54096 vdd.n30189 vdd.n30188 0.894
R54097 vdd.n32737 vdd.n30699 0.892
R54098 vdd.n31451 vdd.n31447 0.886
R54099 vdd.n24934 vdd.n24933 0.874
R54100 vdd.n29023 vdd.n29022 0.872
R54101 vdd.n385 vdd.n384 0.862
R54102 vdd.n31593 vdd.n31592 0.861
R54103 vdd.n1241 vdd.n1237 0.853
R54104 vdd.n2496 vdd.n2492 0.853
R54105 vdd.n2526 vdd.n2522 0.853
R54106 vdd.n3815 vdd.n3811 0.853
R54107 vdd.n3898 vdd.n3894 0.853
R54108 vdd.n3937 vdd.n3933 0.853
R54109 vdd.n33854 vdd.n33853 0.847
R54110 vdd.n954 vdd.n953 0.847
R54111 vdd.n28101 vdd.n28100 0.841
R54112 vdd.n28095 vdd.n28094 0.841
R54113 vdd.n30695 vdd.n30694 0.841
R54114 vdd.n30680 vdd.n30679 0.84
R54115 vdd.n33863 vdd.n33701 0.839
R54116 vdd.n28096 vdd.n28095 0.82
R54117 vdd.n30696 vdd.n30695 0.82
R54118 vdd.n35680 vdd.n35679 0.818
R54119 vdd.n33256 vdd.n33255 0.818
R54120 vdd.n37192 vdd.n37191 0.818
R54121 vdd.n32948 vdd.n32947 0.818
R54122 vdd.n37592 vdd.n37591 0.818
R54123 vdd.n35678 vdd.n35677 0.818
R54124 vdd.n33254 vdd.n33253 0.818
R54125 vdd.n37190 vdd.n37189 0.818
R54126 vdd.n37232 vdd.n37231 0.818
R54127 vdd.n32946 vdd.n32945 0.818
R54128 vdd.n32933 vdd.n32932 0.818
R54129 vdd.n37590 vdd.n37589 0.818
R54130 vdd.n37237 vdd.n37236 0.818
R54131 vdd.n32935 vdd.n32934 0.818
R54132 vdd.n30314 vdd.n30313 0.818
R54133 vdd.n30556 vdd.n30555 0.818
R54134 vdd.n1833 vdd.n1832 0.813
R54135 vdd.n32394 vdd.n32393 0.813
R54136 vdd.n27656 vdd.n27655 0.812
R54137 vdd.n26078 vdd.n26077 0.812
R54138 vdd.n32102 vdd.n32100 0.801
R54139 vdd.n32128 vdd.n32124 0.782
R54140 vdd.n10167 vdd.n10144 0.778
R54141 vdd.n16770 vdd.n16769 0.778
R54142 vdd.n24792 vdd.n24791 0.777
R54143 vdd.n25121 vdd.n25120 0.777
R54144 vdd.n32131 vdd.n32129 0.765
R54145 vdd.t200 vdd.n24498 0.753
R54146 vdd.n33743 vdd.n33742 0.752
R54147 vdd.n33669 vdd.n33668 0.752
R54148 vdd.n33500 vdd.n33499 0.752
R54149 vdd.n33522 vdd.n33521 0.752
R54150 vdd.n33468 vdd.n33467 0.752
R54151 vdd.n33450 vdd.n33449 0.752
R54152 vdd.n34191 vdd.n34190 0.752
R54153 vdd.n34105 vdd.n34104 0.752
R54154 vdd.n34121 vdd.n34120 0.752
R54155 vdd.n34059 vdd.n34058 0.752
R54156 vdd.n33908 vdd.n33907 0.752
R54157 vdd.n34375 vdd.n34374 0.752
R54158 vdd.n34362 vdd.n34361 0.752
R54159 vdd.n33989 vdd.n33988 0.752
R54160 vdd.n35151 vdd.n35150 0.752
R54161 vdd.n35220 vdd.n35219 0.752
R54162 vdd.n35077 vdd.n35076 0.752
R54163 vdd.n35398 vdd.n35397 0.752
R54164 vdd.n35378 vdd.n35377 0.752
R54165 vdd.n35508 vdd.n35507 0.752
R54166 vdd.n35484 vdd.n35483 0.752
R54167 vdd.n35301 vdd.n35300 0.752
R54168 vdd.n34717 vdd.n34716 0.752
R54169 vdd.n34956 vdd.n34955 0.752
R54170 vdd.n34975 vdd.n34974 0.752
R54171 vdd.n34633 vdd.n34632 0.752
R54172 vdd.n34490 vdd.n34489 0.752
R54173 vdd.n34801 vdd.n34800 0.752
R54174 vdd.n34788 vdd.n34787 0.752
R54175 vdd.n34566 vdd.n34565 0.752
R54176 vdd.n917 vdd.n916 0.752
R54177 vdd.n1062 vdd.n1061 0.752
R54178 vdd.n990 vdd.n989 0.752
R54179 vdd.n1003 vdd.n1002 0.752
R54180 vdd.n708 vdd.n707 0.752
R54181 vdd.n769 vdd.n768 0.752
R54182 vdd.n363 vdd.n362 0.752
R54183 vdd.n218 vdd.n217 0.752
R54184 vdd.n194 vdd.n193 0.752
R54185 vdd.n464 vdd.n463 0.752
R54186 vdd.n482 vdd.n481 0.752
R54187 vdd.n6277 vdd.n6276 0.752
R54188 vdd.n6344 vdd.n6343 0.752
R54189 vdd.n6182 vdd.n6181 0.752
R54190 vdd.n6089 vdd.n6088 0.752
R54191 vdd.n6068 vdd.n6067 0.752
R54192 vdd.n5988 vdd.n5987 0.752
R54193 vdd.n5813 vdd.n5812 0.752
R54194 vdd.n5892 vdd.n5891 0.752
R54195 vdd.n5464 vdd.n5463 0.752
R54196 vdd.n5703 vdd.n5702 0.752
R54197 vdd.n5722 vdd.n5721 0.752
R54198 vdd.n5380 vdd.n5379 0.752
R54199 vdd.n5237 vdd.n5236 0.752
R54200 vdd.n5548 vdd.n5547 0.752
R54201 vdd.n5535 vdd.n5534 0.752
R54202 vdd.n5313 vdd.n5312 0.752
R54203 vdd.n4781 vdd.n4779 0.752
R54204 vdd.n4764 vdd.n4763 0.752
R54205 vdd.n4987 vdd.n4986 0.752
R54206 vdd.n5174 vdd.n5173 0.752
R54207 vdd.n5146 vdd.n5145 0.752
R54208 vdd.n4944 vdd.n4943 0.752
R54209 vdd.n4291 vdd.n4290 0.752
R54210 vdd.n4530 vdd.n4529 0.752
R54211 vdd.n4552 vdd.n4551 0.752
R54212 vdd.n4210 vdd.n4209 0.752
R54213 vdd.n4067 vdd.n4066 0.752
R54214 vdd.n4375 vdd.n4374 0.752
R54215 vdd.n4362 vdd.n4361 0.752
R54216 vdd.n4144 vdd.n4143 0.752
R54217 vdd.n30200 vdd.n30199 0.752
R54218 vdd.n31174 vdd.n31173 0.752
R54219 vdd.n32272 vdd.n32271 0.752
R54220 vdd.n32127 vdd.n32126 0.752
R54221 vdd.n32073 vdd.n32072 0.752
R54222 vdd.n31946 vdd.n31945 0.752
R54223 vdd.n32490 vdd.n32489 0.752
R54224 vdd.n36032 vdd.n36025 0.752
R54225 vdd.n36046 vdd.n36039 0.752
R54226 vdd.n36263 vdd.n36256 0.752
R54227 vdd.n36277 vdd.n36270 0.752
R54228 vdd.n36494 vdd.n36487 0.752
R54229 vdd.n36508 vdd.n36501 0.752
R54230 vdd.n36725 vdd.n36718 0.752
R54231 vdd.n36739 vdd.n36732 0.752
R54232 vdd.n36956 vdd.n36949 0.752
R54233 vdd.n36970 vdd.n36963 0.752
R54234 vdd.n33148 vdd.n33141 0.752
R54235 vdd.n35642 vdd.n35635 0.752
R54236 vdd.n37324 vdd.n37317 0.752
R54237 vdd.n37354 vdd.n37347 0.752
R54238 vdd.n35669 vdd.n35662 0.752
R54239 vdd.n32831 vdd.n32824 0.752
R54240 vdd.n38025 vdd.n38018 0.752
R54241 vdd.n38011 vdd.n38004 0.752
R54242 vdd.n37794 vdd.n37787 0.752
R54243 vdd.n37780 vdd.n37773 0.752
R54244 vdd.n28222 vdd.n28215 0.752
R54245 vdd.n28236 vdd.n28229 0.752
R54246 vdd.n28453 vdd.n28446 0.752
R54247 vdd.n28467 vdd.n28460 0.752
R54248 vdd.n28684 vdd.n28677 0.752
R54249 vdd.n28698 vdd.n28691 0.752
R54250 vdd.n28091 vdd.n28090 0.752
R54251 vdd.n28066 vdd.n28065 0.752
R54252 vdd.n28975 vdd.n28974 0.752
R54253 vdd.n27752 vdd.n27751 0.752
R54254 vdd.n27987 vdd.n27986 0.752
R54255 vdd.n27986 vdd.n27979 0.752
R54256 vdd.n27883 vdd.n27875 0.752
R54257 vdd.n27883 vdd.n27876 0.752
R54258 vdd.n27916 vdd.n27907 0.752
R54259 vdd.n27939 vdd.n27938 0.752
R54260 vdd.n29881 vdd.n29880 0.752
R54261 vdd.n30010 vdd.n30009 0.752
R54262 vdd.n30193 vdd.n30192 0.752
R54263 vdd.n27329 vdd.n27328 0.752
R54264 vdd.n27379 vdd.n27378 0.752
R54265 vdd.n27397 vdd.n27396 0.752
R54266 vdd.n27474 vdd.n27473 0.752
R54267 vdd.n27269 vdd.n27268 0.752
R54268 vdd.n27542 vdd.n27541 0.752
R54269 vdd.n27599 vdd.n27598 0.752
R54270 vdd.n27616 vdd.n27615 0.752
R54271 vdd.n25781 vdd.n25780 0.752
R54272 vdd.n25822 vdd.n25821 0.752
R54273 vdd.n25843 vdd.n25842 0.752
R54274 vdd.n25712 vdd.n25711 0.752
R54275 vdd.n25924 vdd.n25923 0.752
R54276 vdd.n25979 vdd.n25978 0.752
R54277 vdd.n26015 vdd.n26014 0.752
R54278 vdd.n26037 vdd.n26036 0.752
R54279 vdd.n25392 vdd.n25391 0.752
R54280 vdd.n25529 vdd.n25528 0.752
R54281 vdd.n25440 vdd.n25439 0.752
R54282 vdd.n25542 vdd.n25540 0.752
R54283 vdd.n25606 vdd.n25605 0.752
R54284 vdd.n25380 vdd.n25379 0.752
R54285 vdd.n26395 vdd.n26394 0.752
R54286 vdd.n26299 vdd.n26298 0.752
R54287 vdd.n1659 vdd.n1655 0.752
R54288 vdd.n1649 vdd.n1645 0.752
R54289 vdd.n1478 vdd.n1474 0.752
R54290 vdd.n1468 vdd.n1464 0.752
R54291 vdd.n1297 vdd.n1293 0.752
R54292 vdd.n26763 vdd.n26759 0.752
R54293 vdd.n26934 vdd.n26930 0.752
R54294 vdd.n26944 vdd.n26940 0.752
R54295 vdd.n27115 vdd.n27111 0.752
R54296 vdd.n27125 vdd.n27121 0.752
R54297 vdd.n1201 vdd.n1200 0.752
R54298 vdd.n1203 vdd.n1202 0.752
R54299 vdd.n2573 vdd.n2572 0.752
R54300 vdd.n2384 vdd.n2383 0.752
R54301 vdd.n2200 vdd.n2199 0.752
R54302 vdd.n3787 vdd.n3785 0.752
R54303 vdd.n2726 vdd.n2725 0.752
R54304 vdd.n2887 vdd.n2883 0.752
R54305 vdd.n2897 vdd.n2893 0.752
R54306 vdd.n3068 vdd.n3064 0.752
R54307 vdd.n3078 vdd.n3074 0.752
R54308 vdd.n3249 vdd.n3245 0.752
R54309 vdd.n3259 vdd.n3255 0.752
R54310 vdd.n3430 vdd.n3426 0.752
R54311 vdd.n3440 vdd.n3436 0.752
R54312 vdd.n3611 vdd.n3607 0.752
R54313 vdd.n3621 vdd.n3617 0.752
R54314 vdd.n31779 vdd.n31778 0.752
R54315 vdd.n13357 vdd.n13356 0.752
R54316 vdd.n13402 vdd.n13401 0.752
R54317 vdd.n13649 vdd.n13648 0.752
R54318 vdd.n13695 vdd.n13694 0.752
R54319 vdd.n13965 vdd.n8624 0.752
R54320 vdd.n8625 vdd.n8613 0.752
R54321 vdd.n14255 vdd.n8402 0.752
R54322 vdd.n8403 vdd.n8391 0.752
R54323 vdd.n14687 vdd.n14682 0.752
R54324 vdd.n14716 vdd.n8111 0.752
R54325 vdd.n14861 vdd.n14853 0.752
R54326 vdd.n14904 vdd.n14903 0.752
R54327 vdd.n13240 vdd.n9182 0.752
R54328 vdd.n13241 vdd.n13240 0.752
R54329 vdd.n13279 vdd.n13278 0.752
R54330 vdd.n13279 vdd.n9153 0.752
R54331 vdd.n13532 vdd.n8961 0.752
R54332 vdd.n13533 vdd.n13532 0.752
R54333 vdd.n13571 vdd.n13570 0.752
R54334 vdd.n13571 vdd.n8932 0.752
R54335 vdd.n13817 vdd.n13816 0.752
R54336 vdd.n13818 vdd.n13817 0.752
R54337 vdd.n13859 vdd.n13858 0.752
R54338 vdd.n13859 vdd.n8705 0.752
R54339 vdd.n14105 vdd.n14103 0.752
R54340 vdd.n14105 vdd.n14104 0.752
R54341 vdd.n14148 vdd.n14147 0.752
R54342 vdd.n14148 vdd.n8482 0.752
R54343 vdd.n14411 vdd.n8293 0.752
R54344 vdd.n14411 vdd.n8294 0.752
R54345 vdd.n14414 vdd.n14413 0.752
R54346 vdd.n14414 vdd.n8267 0.752
R54347 vdd.n11741 vdd.n11726 0.752
R54348 vdd.n11736 vdd.n11731 0.752
R54349 vdd.n11697 vdd.n11694 0.752
R54350 vdd.n11710 vdd.n11709 0.752
R54351 vdd.n11825 vdd.n11821 0.752
R54352 vdd.n11831 vdd.n11830 0.752
R54353 vdd.n11859 vdd.n11838 0.752
R54354 vdd.n11853 vdd.n11852 0.752
R54355 vdd.n22166 vdd.n22165 0.752
R54356 vdd.n24096 vdd.n24095 0.752
R54357 vdd.n24070 vdd.n24069 0.752
R54358 vdd.n23864 vdd.n23863 0.752
R54359 vdd.n23838 vdd.n23837 0.752
R54360 vdd.n23632 vdd.n23631 0.752
R54361 vdd.n23150 vdd.n23149 0.752
R54362 vdd.n23176 vdd.n23175 0.752
R54363 vdd.n23382 vdd.n23381 0.752
R54364 vdd.n23408 vdd.n23407 0.752
R54365 vdd.n23614 vdd.n23613 0.752
R54366 vdd.n22571 vdd.n22570 0.752
R54367 vdd.n22597 vdd.n22596 0.752
R54368 vdd.n22803 vdd.n22802 0.752
R54369 vdd.n22829 vdd.n22828 0.752
R54370 vdd.n23035 vdd.n23034 0.752
R54371 vdd.n22187 vdd.n22186 0.752
R54372 vdd.n22201 vdd.n22197 0.752
R54373 vdd.n22045 vdd.n22044 0.752
R54374 vdd.n22059 vdd.n22055 0.752
R54375 vdd.n19269 vdd.n19260 0.752
R54376 vdd.n19257 vdd.n19248 0.752
R54377 vdd.n19213 vdd.n19204 0.752
R54378 vdd.n19201 vdd.n19192 0.752
R54379 vdd.n19855 vdd.n19846 0.752
R54380 vdd.n19867 vdd.n19858 0.752
R54381 vdd.n19923 vdd.n19914 0.752
R54382 vdd.n19935 vdd.n19926 0.752
R54383 vdd.n21530 vdd.n21521 0.752
R54384 vdd.n21512 vdd.n21503 0.752
R54385 vdd.n21271 vdd.n21262 0.752
R54386 vdd.n21253 vdd.n21244 0.752
R54387 vdd.n21014 vdd.n21013 0.752
R54388 vdd.n19139 vdd.n19135 0.752
R54389 vdd.n18905 vdd.n18896 0.752
R54390 vdd.n18887 vdd.n18878 0.752
R54391 vdd.n18646 vdd.n18637 0.752
R54392 vdd.n18628 vdd.n18619 0.752
R54393 vdd.n20394 vdd.n20393 0.752
R54394 vdd.n20371 vdd.n20370 0.752
R54395 vdd.n20158 vdd.n20157 0.752
R54396 vdd.n20135 vdd.n20134 0.752
R54397 vdd.n21814 vdd.n21813 0.752
R54398 vdd.n21916 vdd.n21912 0.752
R54399 vdd.n21922 vdd.n21921 0.752
R54400 vdd.n21950 vdd.n21929 0.752
R54401 vdd.n21944 vdd.n21943 0.752
R54402 vdd.n24736 vdd.n24735 0.752
R54403 vdd.n24752 vdd.n24751 0.752
R54404 vdd.n25168 vdd.n25167 0.752
R54405 vdd.n25154 vdd.n25153 0.752
R54406 vdd.n2294 vdd.n2133 0.75
R54407 vdd.n34443 vdd.n34440 0.75
R54408 vdd.n32737 vdd.n29953 0.738
R54409 vdd.n587 vdd.n586 0.737
R54410 vdd.n33863 vdd.n33474 0.736
R54411 vdd.n1173 vdd.n787 0.736
R54412 vdd.n5189 vdd.n4800 0.734
R54413 vdd.n4016 vdd.n2678 0.718
R54414 vdd.n10490 vdd.n10123 0.711
R54415 vdd.n10397 vdd.n10396 0.711
R54416 vdd.n10396 vdd.n10334 0.711
R54417 vdd.n10372 vdd.n10353 0.711
R54418 vdd.n10372 vdd.n10354 0.711
R54419 vdd.n9430 vdd.n9429 0.711
R54420 vdd.n9431 vdd.n9430 0.711
R54421 vdd.n12982 vdd.n12981 0.711
R54422 vdd.n12981 vdd.n9424 0.711
R54423 vdd.n12896 vdd.n9574 0.711
R54424 vdd.n12896 vdd.n9575 0.711
R54425 vdd.n9644 vdd.n9632 0.711
R54426 vdd.n9644 vdd.n9633 0.711
R54427 vdd.n9790 vdd.n9789 0.711
R54428 vdd.n9791 vdd.n9790 0.711
R54429 vdd.n12774 vdd.n12773 0.711
R54430 vdd.n12773 vdd.n9784 0.711
R54431 vdd.n12688 vdd.n9933 0.711
R54432 vdd.n12688 vdd.n9934 0.711
R54433 vdd.n10004 vdd.n9992 0.711
R54434 vdd.n10004 vdd.n9993 0.711
R54435 vdd.n10163 vdd.n10148 0.711
R54436 vdd.n12524 vdd.n12523 0.711
R54437 vdd.n12492 vdd.n12491 0.711
R54438 vdd.n12468 vdd.n12467 0.711
R54439 vdd.n12445 vdd.n10654 0.711
R54440 vdd.n12423 vdd.n12422 0.711
R54441 vdd.n12386 vdd.n10724 0.711
R54442 vdd.n10789 vdd.n10784 0.711
R54443 vdd.n10834 vdd.n10832 0.711
R54444 vdd.n10877 vdd.n10854 0.711
R54445 vdd.n10935 vdd.n10929 0.711
R54446 vdd.n12273 vdd.n10925 0.711
R54447 vdd.n10999 vdd.n10998 0.711
R54448 vdd.n12220 vdd.n11035 0.711
R54449 vdd.n12187 vdd.n11088 0.711
R54450 vdd.n12170 vdd.n11110 0.711
R54451 vdd.n12142 vdd.n11149 0.711
R54452 vdd.n11213 vdd.n11198 0.711
R54453 vdd.n11264 vdd.n11244 0.711
R54454 vdd.n11298 vdd.n11292 0.711
R54455 vdd.n11343 vdd.n11341 0.711
R54456 vdd.n11386 vdd.n11363 0.711
R54457 vdd.n11479 vdd.n11473 0.711
R54458 vdd.n11967 vdd.n11434 0.711
R54459 vdd.n11936 vdd.n11935 0.711
R54460 vdd.n15413 vdd.n15412 0.711
R54461 vdd.n15412 vdd.n15404 0.711
R54462 vdd.n15429 vdd.n15422 0.711
R54463 vdd.n15431 vdd.n15429 0.711
R54464 vdd.n15663 vdd.n15662 0.711
R54465 vdd.n15662 vdd.n15652 0.711
R54466 vdd.n15682 vdd.n15672 0.711
R54467 vdd.n15684 vdd.n15682 0.711
R54468 vdd.n15919 vdd.n15918 0.711
R54469 vdd.n15918 vdd.n15908 0.711
R54470 vdd.n15938 vdd.n15928 0.711
R54471 vdd.n15940 vdd.n15938 0.711
R54472 vdd.n16175 vdd.n16174 0.711
R54473 vdd.n16174 vdd.n16164 0.711
R54474 vdd.n16194 vdd.n16184 0.711
R54475 vdd.n16196 vdd.n16194 0.711
R54476 vdd.n16431 vdd.n16430 0.711
R54477 vdd.n16430 vdd.n16420 0.711
R54478 vdd.n16450 vdd.n16440 0.711
R54479 vdd.n16452 vdd.n16450 0.711
R54480 vdd.n16579 vdd.n16578 0.711
R54481 vdd.n16834 vdd.n16833 0.711
R54482 vdd.n16966 vdd.n16965 0.711
R54483 vdd.n17011 vdd.n17009 0.711
R54484 vdd.n17080 vdd.n17079 0.711
R54485 vdd.n17132 vdd.n17131 0.711
R54486 vdd.n17238 vdd.n17237 0.711
R54487 vdd.n17283 vdd.n17281 0.711
R54488 vdd.n17352 vdd.n17351 0.711
R54489 vdd.n17404 vdd.n17403 0.711
R54490 vdd.n17510 vdd.n17509 0.711
R54491 vdd.n17555 vdd.n17553 0.711
R54492 vdd.n17610 vdd.n17609 0.711
R54493 vdd.n17662 vdd.n17661 0.711
R54494 vdd.n17768 vdd.n17767 0.711
R54495 vdd.n17813 vdd.n17811 0.711
R54496 vdd.n17881 vdd.n17880 0.711
R54497 vdd.n17933 vdd.n17932 0.711
R54498 vdd.n18039 vdd.n18038 0.711
R54499 vdd.n18084 vdd.n18082 0.711
R54500 vdd.n18153 vdd.n18152 0.711
R54501 vdd.n18205 vdd.n18204 0.711
R54502 vdd.n18305 vdd.n18304 0.711
R54503 vdd.n18329 vdd.n18321 0.711
R54504 vdd.n18410 vdd.n18409 0.711
R54505 vdd.n21660 vdd.n21658 0.703
R54506 vdd.n21672 vdd.n21669 0.703
R54507 vdd.n21394 vdd.n21391 0.703
R54508 vdd.n21380 vdd.n21377 0.703
R54509 vdd.n21135 vdd.n21132 0.703
R54510 vdd.n21121 vdd.n21118 0.703
R54511 vdd.n19028 vdd.n19025 0.703
R54512 vdd.n19014 vdd.n19011 0.703
R54513 vdd.n18769 vdd.n18766 0.703
R54514 vdd.n18755 vdd.n18752 0.703
R54515 vdd.n18510 vdd.n18507 0.703
R54516 vdd.n18496 vdd.n18493 0.703
R54517 vdd.n3663 vdd.n3662 0.7
R54518 vdd.n3669 vdd.n3668 0.7
R54519 vdd.n35687 vdd.n35686 0.697
R54520 vdd.n37151 vdd.n37150 0.697
R54521 vdd.n37179 vdd.n37178 0.697
R54522 vdd.n32992 vdd.n32991 0.697
R54523 vdd.n32978 vdd.n32977 0.697
R54524 vdd.n37526 vdd.n37525 0.697
R54525 vdd.n37572 vdd.n37571 0.697
R54526 vdd.n29724 vdd.n29723 0.697
R54527 vdd.n9123 vdd.n9098 0.697
R54528 vdd.n13394 vdd.n13393 0.697
R54529 vdd.n8902 vdd.n8878 0.697
R54530 vdd.n13686 vdd.n13685 0.697
R54531 vdd.n13913 vdd.n13912 0.697
R54532 vdd.n8610 vdd.n8607 0.697
R54533 vdd.n14203 vdd.n14202 0.697
R54534 vdd.n8388 vdd.n8385 0.697
R54535 vdd.n19282 vdd.n19281 0.697
R54536 vdd.n19246 vdd.n19245 0.697
R54537 vdd.n19226 vdd.n19225 0.697
R54538 vdd.n19189 vdd.n19188 0.697
R54539 vdd.n19843 vdd.n19842 0.697
R54540 vdd.n19880 vdd.n19879 0.697
R54541 vdd.n19912 vdd.n19911 0.697
R54542 vdd.n19948 vdd.n19947 0.697
R54543 vdd.n27208 vdd.n27207 0.689
R54544 vdd.n4016 vdd.n2683 0.687
R54545 vdd.n25551 vdd.n25550 0.677
R54546 vdd.n35896 vdd.n35895 0.67
R54547 vdd.n35945 vdd.n35944 0.67
R54548 vdd.n36127 vdd.n36126 0.67
R54549 vdd.n36176 vdd.n36175 0.67
R54550 vdd.n36358 vdd.n36357 0.67
R54551 vdd.n36407 vdd.n36406 0.67
R54552 vdd.n36589 vdd.n36588 0.67
R54553 vdd.n36638 vdd.n36637 0.67
R54554 vdd.n36820 vdd.n36819 0.67
R54555 vdd.n36869 vdd.n36868 0.67
R54556 vdd.n37055 vdd.n37054 0.67
R54557 vdd.n37094 vdd.n37093 0.67
R54558 vdd.n2155 vdd.n2154 0.67
R54559 vdd.n33056 vdd.n33055 0.67
R54560 vdd.n32926 vdd.n32925 0.67
R54561 vdd.n37467 vdd.n37466 0.67
R54562 vdd.n38149 vdd.n38148 0.67
R54563 vdd.n38106 vdd.n38105 0.67
R54564 vdd.n37924 vdd.n37923 0.67
R54565 vdd.n37875 vdd.n37874 0.67
R54566 vdd.n37693 vdd.n37692 0.67
R54567 vdd.n37644 vdd.n37643 0.67
R54568 vdd.n28317 vdd.n28316 0.67
R54569 vdd.n28366 vdd.n28365 0.67
R54570 vdd.n28548 vdd.n28547 0.67
R54571 vdd.n28597 vdd.n28596 0.67
R54572 vdd.n28779 vdd.n28778 0.67
R54573 vdd.n28162 vdd.n28161 0.67
R54574 vdd.n31842 vdd.n31841 0.67
R54575 vdd.n29027 vdd.n29026 0.67
R54576 vdd.n29869 vdd.n29868 0.67
R54577 vdd.n29835 vdd.n29834 0.67
R54578 vdd.n31090 vdd.n31089 0.67
R54579 vdd.n30544 vdd.n30543 0.67
R54580 vdd.n36973 vdd.n35699 0.658
R54581 vdd.n36973 vdd.n35693 0.658
R54582 vdd.n11819 vdd.n11818 0.649
R54583 vdd.n21910 vdd.n21909 0.649
R54584 vdd.n10455 vdd.n10454 0.645
R54585 vdd.n10441 vdd.n10297 0.645
R54586 vdd.n15301 vdd.n15300 0.645
R54587 vdd.n15323 vdd.n15322 0.645
R54588 vdd.n11784 vdd.n11783 0.645
R54589 vdd.n21876 vdd.n21875 0.645
R54590 vdd.n25563 vdd.n25562 0.643
R54591 vdd.n9341 vdd.n9318 0.641
R54592 vdd.t225 vdd.n13042 0.641
R54593 vdd.n13032 vdd.n13031 0.641
R54594 vdd.n12947 vdd.n12946 0.641
R54595 vdd.n9541 vdd.n9540 0.641
R54596 vdd.n9701 vdd.n9680 0.641
R54597 vdd.n12824 vdd.n12823 0.641
R54598 vdd.t301 vdd.n12785 0.641
R54599 vdd.n12776 vdd.t387 0.641
R54600 vdd.n12739 vdd.n12738 0.641
R54601 vdd.n9901 vdd.n9885 0.641
R54602 vdd.n12697 vdd.t353 0.641
R54603 vdd.n10154 vdd.t299 0.641
R54604 vdd.n12615 vdd.n12614 0.641
R54605 vdd.n10487 vdd.t80 0.641
R54606 vdd.n12489 vdd.n12488 0.641
R54607 vdd.n12482 vdd.n10584 0.641
R54608 vdd.n12384 vdd.n12383 0.641
R54609 vdd.n12372 vdd.n10763 0.641
R54610 vdd.n10937 vdd.t306 0.641
R54611 vdd.n10938 vdd.n10937 0.641
R54612 vdd.n12279 vdd.n12278 0.641
R54613 vdd.n11075 vdd.t377 0.641
R54614 vdd.n11099 vdd.n11086 0.641
R54615 vdd.n11119 vdd.n11118 0.641
R54616 vdd.n12084 vdd.n11240 0.641
R54617 vdd.n12066 vdd.n11273 0.641
R54618 vdd.n11482 vdd.n11481 0.641
R54619 vdd.n11973 vdd.n11972 0.641
R54620 vdd.n11945 vdd.t190 0.641
R54621 vdd.n15526 vdd.n15525 0.641
R54622 vdd.n15551 vdd.t195 0.641
R54623 vdd.n15557 vdd.n15556 0.641
R54624 vdd.n15782 vdd.n15781 0.641
R54625 vdd.n15813 vdd.n15812 0.641
R54626 vdd.n16038 vdd.n16037 0.641
R54627 vdd.n16069 vdd.n16068 0.641
R54628 vdd.n15158 vdd.t269 0.641
R54629 vdd.t2 vdd.n16191 0.641
R54630 vdd.n16294 vdd.n16293 0.641
R54631 vdd.n16325 vdd.n16324 0.641
R54632 vdd.t16 vdd.n16391 0.641
R54633 vdd.n16548 vdd.t259 0.641
R54634 vdd.n16556 vdd.n16555 0.641
R54635 vdd.n15075 vdd.t336 0.641
R54636 vdd.n16963 vdd.n16962 0.641
R54637 vdd.n16991 vdd.n16990 0.641
R54638 vdd.n17235 vdd.n17234 0.641
R54639 vdd.n17263 vdd.n17262 0.641
R54640 vdd.n17507 vdd.t254 0.641
R54641 vdd.n17507 vdd.n17506 0.641
R54642 vdd.n17535 vdd.n17534 0.641
R54643 vdd.t10 vdd.n17716 0.641
R54644 vdd.n17765 vdd.n17764 0.641
R54645 vdd.n17793 vdd.n17792 0.641
R54646 vdd.n18036 vdd.n18035 0.641
R54647 vdd.n18064 vdd.n18063 0.641
R54648 vdd.n18302 vdd.n18301 0.641
R54649 vdd.n15034 vdd.n15033 0.641
R54650 vdd.t220 vdd.n15008 0.641
R54651 vdd.n5189 vdd.n5186 0.64
R54652 vdd.n13177 vdd.t320 0.639
R54653 vdd.n10389 vdd.n9297 0.637
R54654 vdd.n15408 vdd.n15407 0.637
R54655 vdd.n12571 vdd.n12570 0.636
R54656 vdd.n34443 vdd.n34072 0.63
R54657 vdd.n35612 vdd.n35234 0.63
R54658 vdd.n35026 vdd.n34647 0.63
R54659 vdd.n6358 vdd.n6357 0.63
R54660 vdd.n5775 vdd.n5394 0.63
R54661 vdd.n4605 vdd.n4224 0.63
R54662 vdd.n29684 vdd.n29683 0.623
R54663 vdd.n24804 vdd.n24803 0.615
R54664 vdd.n25109 vdd.n25108 0.615
R54665 vdd.n33798 vdd.n33797 0.614
R54666 vdd.n829 vdd.n828 0.614
R54667 vdd.n323 vdd.n322 0.613
R54668 vdd.n34162 vdd.n34161 0.613
R54669 vdd.n35311 vdd.n35310 0.613
R54670 vdd.n34735 vdd.n34734 0.613
R54671 vdd.n5863 vdd.n5862 0.613
R54672 vdd.n5482 vdd.n5481 0.613
R54673 vdd.n4309 vdd.n4308 0.613
R54674 vdd.n4905 vdd.n4904 0.612
R54675 vdd.n13238 vdd.n9185 0.611
R54676 vdd.n13238 vdd.n13237 0.611
R54677 vdd.n13246 vdd.n13245 0.611
R54678 vdd.n9179 vdd.n9165 0.611
R54679 vdd.n13276 vdd.n9158 0.611
R54680 vdd.n9151 vdd.n9140 0.611
R54681 vdd.n13304 vdd.n9140 0.611
R54682 vdd.n9132 vdd.n9131 0.611
R54683 vdd.n9104 vdd.n9093 0.611
R54684 vdd.n9125 vdd.n9122 0.611
R54685 vdd.n9122 vdd.n9070 0.611
R54686 vdd.n13359 vdd.n9089 0.611
R54687 vdd.n13376 vdd.n13375 0.611
R54688 vdd.n13378 vdd.n13377 0.611
R54689 vdd.n13404 vdd.n9046 0.611
R54690 vdd.n9056 vdd.n9046 0.611
R54691 vdd.n8981 vdd.t316 0.611
R54692 vdd.n13530 vdd.n8964 0.611
R54693 vdd.n13530 vdd.n13529 0.611
R54694 vdd.n13538 vdd.n13537 0.611
R54695 vdd.n8958 vdd.n8944 0.611
R54696 vdd.n13568 vdd.n8936 0.611
R54697 vdd.n8930 vdd.n8918 0.611
R54698 vdd.n13596 vdd.n8918 0.611
R54699 vdd.n8910 vdd.n8909 0.611
R54700 vdd.n8883 vdd.n8873 0.611
R54701 vdd.n8904 vdd.n8901 0.611
R54702 vdd.n8901 vdd.n8850 0.611
R54703 vdd.n13651 vdd.n8869 0.611
R54704 vdd.n13668 vdd.n13667 0.611
R54705 vdd.n13670 vdd.n13669 0.611
R54706 vdd.n13697 vdd.n8825 0.611
R54707 vdd.n8836 vdd.n8825 0.611
R54708 vdd.n8739 vdd.n8738 0.611
R54709 vdd.n13820 vdd.n8739 0.611
R54710 vdd.n13823 vdd.n13822 0.611
R54711 vdd.n13864 vdd.n8712 0.611
R54712 vdd.n13856 vdd.n8719 0.611
R54713 vdd.n13870 vdd.n8708 0.611
R54714 vdd.n8708 vdd.n8681 0.611
R54715 vdd.n13889 vdd.n13888 0.611
R54716 vdd.n8677 vdd.n8646 0.611
R54717 vdd.n13915 vdd.n8657 0.611
R54718 vdd.n8663 vdd.n8657 0.611
R54719 vdd.n13967 vdd.n8619 0.611
R54720 vdd.n13961 vdd.n13960 0.611
R54721 vdd.n8632 vdd.n8631 0.611
R54722 vdd.n13976 vdd.n13974 0.611
R54723 vdd.n13976 vdd.n13975 0.611
R54724 vdd.n14108 vdd.n14107 0.611
R54725 vdd.n14107 vdd.n8525 0.611
R54726 vdd.n14127 vdd.n14126 0.611
R54727 vdd.n14153 vdd.n8489 0.611
R54728 vdd.n14145 vdd.n8497 0.611
R54729 vdd.n14159 vdd.n8485 0.611
R54730 vdd.n8485 vdd.n8457 0.611
R54731 vdd.n14168 vdd.t326 0.611
R54732 vdd.n14178 vdd.n14177 0.611
R54733 vdd.n8453 vdd.n8426 0.611
R54734 vdd.n14205 vdd.n8436 0.611
R54735 vdd.n8438 vdd.n8436 0.611
R54736 vdd.n14257 vdd.n8397 0.611
R54737 vdd.n14251 vdd.n14250 0.611
R54738 vdd.n8410 vdd.n8408 0.611
R54739 vdd.n14266 vdd.n14264 0.611
R54740 vdd.n14266 vdd.n14265 0.611
R54741 vdd.t317 vdd.n14407 0.611
R54742 vdd.n14409 vdd.n14408 0.611
R54743 vdd.n14409 vdd.n8273 0.611
R54744 vdd.n8285 vdd.n8274 0.611
R54745 vdd.n14420 vdd.n14419 0.611
R54746 vdd.n14461 vdd.n8241 0.611
R54747 vdd.n14452 vdd.n14451 0.611
R54748 vdd.n8234 vdd.n8233 0.611
R54749 vdd.t321 vdd.n14487 0.611
R54750 vdd.n8223 vdd.n8215 0.611
R54751 vdd.n14645 vdd.n14644 0.611
R54752 vdd.n11675 vdd.n11674 0.605
R54753 vdd.n21851 vdd.n21850 0.605
R54754 vdd.n258 vdd.n257 0.586
R54755 vdd.n19367 vdd.t244 0.586
R54756 vdd.n19414 vdd.n19411 0.586
R54757 vdd.n19431 vdd.n19428 0.586
R54758 vdd.n19617 vdd.n19614 0.586
R54759 vdd.n19634 vdd.n19631 0.586
R54760 vdd.n19819 vdd.n19816 0.586
R54761 vdd.n19169 vdd.n19166 0.586
R54762 vdd.n20839 vdd.n20836 0.586
R54763 vdd.n20825 vdd.n20822 0.586
R54764 vdd.n20637 vdd.n20634 0.586
R54765 vdd.n20623 vdd.n20620 0.586
R54766 vdd.n20576 vdd.t241 0.586
R54767 vdd.n20403 vdd.t265 0.586
R54768 vdd.n19998 vdd.n19997 0.586
R54769 vdd.n20010 vdd.n20009 0.586
R54770 vdd.n20140 vdd.t268 0.586
R54771 vdd.n11605 vdd.n11604 0.585
R54772 vdd.n21698 vdd.n21697 0.585
R54773 vdd.n14702 vdd.t297 0.584
R54774 vdd.n14788 vdd.n14787 0.584
R54775 vdd.n14780 vdd.n8064 0.584
R54776 vdd.n14876 vdd.t293 0.584
R54777 vdd.n35026 vdd.n35025 0.563
R54778 vdd.n5775 vdd.n5772 0.563
R54779 vdd.n4605 vdd.n4602 0.563
R54780 vdd.n35612 vdd.n35611 0.56
R54781 vdd.n3663 vdd.t89 0.553
R54782 vdd.n3663 vdd.t230 0.553
R54783 vdd.n3669 vdd.t231 0.553
R54784 vdd.n33853 vdd.t78 0.553
R54785 vdd.n33853 vdd.t75 0.553
R54786 vdd.n34010 vdd.t65 0.553
R54787 vdd.n34010 vdd.t81 0.553
R54788 vdd.n35173 vdd.t44 0.553
R54789 vdd.n35173 vdd.t69 0.553
R54790 vdd.n34598 vdd.t58 0.553
R54791 vdd.n34598 vdd.t48 0.553
R54792 vdd.n953 vdd.t74 0.553
R54793 vdd.n953 vdd.t91 0.553
R54794 vdd.n384 vdd.t52 0.553
R54795 vdd.n384 vdd.t41 0.553
R54796 vdd.n6310 vdd.t67 0.553
R54797 vdd.n6310 vdd.t57 0.553
R54798 vdd.n5345 vdd.t86 0.553
R54799 vdd.n5345 vdd.t98 0.553
R54800 vdd.n4656 vdd.t96 0.553
R54801 vdd.n4656 vdd.t51 0.553
R54802 vdd.n4176 vdd.t40 0.553
R54803 vdd.n4176 vdd.t93 0.553
R54804 vdd.n35692 vdd.t209 0.553
R54805 vdd.n35698 vdd.t210 0.553
R54806 vdd.n35698 vdd.t61 0.553
R54807 vdd.n27223 vdd.t234 0.553
R54808 vdd.n27218 vdd.t90 0.553
R54809 vdd.n27218 vdd.t233 0.553
R54810 vdd.n28830 vdd.t218 0.553
R54811 vdd.n28830 vdd.t64 0.553
R54812 vdd.n28824 vdd.t217 0.553
R54813 vdd.n27655 vdd.t79 0.553
R54814 vdd.n27655 vdd.t77 0.553
R54815 vdd.n26077 vdd.t76 0.553
R54816 vdd.n26077 vdd.t92 0.553
R54817 vdd.n25396 vdd.t55 0.553
R54818 vdd.n25396 vdd.t45 0.553
R54819 vdd.n32737 vdd.n29039 0.548
R54820 vdd.n32406 vdd.n32405 0.533
R54821 vdd.n32100 vdd.n32099 0.533
R54822 vdd.n32510 vdd.n32509 0.533
R54823 vdd.n26342 vdd.n26341 0.533
R54824 vdd.n1836 vdd.n1251 0.531
R54825 vdd.n3997 vdd.n3747 0.53
R54826 vdd.n31463 vdd.n31462 0.505
R54827 vdd.n31600 vdd.n31599 0.505
R54828 vdd.n26313 vdd.n26312 0.505
R54829 vdd.n11884 vdd.n11881 0.503
R54830 vdd.n21975 vdd.n21972 0.503
R54831 vdd.n3683 vdd.n2711 0.5
R54832 vdd.n2248 vdd.n2206 0.5
R54833 vdd.n1827 vdd.n1255 0.5
R54834 vdd.n11783 vdd.n11778 0.5
R54835 vdd.n21875 vdd.n21871 0.5
R54836 vdd.n3680 vdd.n2712 0.499
R54837 vdd.n12570 vdd.n12569 0.488
R54838 vdd.n15119 vdd.n15118 0.488
R54839 vdd.n27657 vdd.n27656 0.484
R54840 vdd.n26079 vdd.n26078 0.484
R54841 vdd.n12597 vdd.n10098 0.474
R54842 vdd.n10096 vdd.n10066 0.474
R54843 vdd.n12603 vdd.n10065 0.474
R54844 vdd.n10457 vdd.n10288 0.474
R54845 vdd.n10450 vdd.n10292 0.474
R54846 vdd.n10301 vdd.n10295 0.474
R54847 vdd.n10439 vdd.n10438 0.474
R54848 vdd.n9336 vdd.n9335 0.474
R54849 vdd.n9348 vdd.n9346 0.474
R54850 vdd.n13039 vdd.n9333 0.474
R54851 vdd.n13034 vdd.n9352 0.474
R54852 vdd.n12944 vdd.n9510 0.474
R54853 vdd.n12939 vdd.n9511 0.474
R54854 vdd.n9535 vdd.n9532 0.474
R54855 vdd.n9544 vdd.n9543 0.474
R54856 vdd.n9696 vdd.n9695 0.474
R54857 vdd.n9708 vdd.n9706 0.474
R54858 vdd.n12831 vdd.n9693 0.474
R54859 vdd.n12826 vdd.n9712 0.474
R54860 vdd.n12736 vdd.n9870 0.474
R54861 vdd.n12731 vdd.n9871 0.474
R54862 vdd.n9896 vdd.n9893 0.474
R54863 vdd.n9904 vdd.n9903 0.474
R54864 vdd.n10152 vdd.n10151 0.474
R54865 vdd.n10164 vdd.n10163 0.474
R54866 vdd.n12619 vdd.n10051 0.474
R54867 vdd.n12617 vdd.n10054 0.474
R54868 vdd.n10184 vdd.n10183 0.474
R54869 vdd.n12491 vdd.n10569 0.474
R54870 vdd.n12480 vdd.n12479 0.474
R54871 vdd.n10682 vdd.n10662 0.474
R54872 vdd.n10694 vdd.n10693 0.474
R54873 vdd.n12386 vdd.n10747 0.474
R54874 vdd.n12374 vdd.n10753 0.474
R54875 vdd.n10849 vdd.n10828 0.474
R54876 vdd.n12328 vdd.n12327 0.474
R54877 vdd.n10935 vdd.n10927 0.474
R54878 vdd.n12281 vdd.n10920 0.474
R54879 vdd.n11020 vdd.n11018 0.474
R54880 vdd.n12230 vdd.n11016 0.474
R54881 vdd.n11097 vdd.n11088 0.474
R54882 vdd.n11121 vdd.n11112 0.474
R54883 vdd.n12129 vdd.n11179 0.474
R54884 vdd.n11203 vdd.n11201 0.474
R54885 vdd.n12082 vdd.n11244 0.474
R54886 vdd.n12069 vdd.n12068 0.474
R54887 vdd.n11358 vdd.n11337 0.474
R54888 vdd.n12022 vdd.n12021 0.474
R54889 vdd.n11479 vdd.n11471 0.474
R54890 vdd.n11975 vdd.n11429 0.474
R54891 vdd.n11522 vdd.n11458 0.474
R54892 vdd.n11537 vdd.n11536 0.474
R54893 vdd.n11942 vdd.n11551 0.474
R54894 vdd.n11938 vdd.n11937 0.474
R54895 vdd.n16594 vdd.n16592 0.474
R54896 vdd.n16688 vdd.n16686 0.474
R54897 vdd.n16701 vdd.n16700 0.474
R54898 vdd.n15296 vdd.n15295 0.474
R54899 vdd.n15307 vdd.n15306 0.474
R54900 vdd.n15327 vdd.n15315 0.474
R54901 vdd.n15317 vdd.n15316 0.474
R54902 vdd.n15521 vdd.n15520 0.474
R54903 vdd.n15535 vdd.n15534 0.474
R54904 vdd.n15561 vdd.n15543 0.474
R54905 vdd.n15545 vdd.n15544 0.474
R54906 vdd.n15777 vdd.n15776 0.474
R54907 vdd.n15791 vdd.n15790 0.474
R54908 vdd.n15817 vdd.n15799 0.474
R54909 vdd.n15801 vdd.n15800 0.474
R54910 vdd.n16033 vdd.n16032 0.474
R54911 vdd.n16047 vdd.n16046 0.474
R54912 vdd.n16073 vdd.n16055 0.474
R54913 vdd.n16057 vdd.n16056 0.474
R54914 vdd.n16289 vdd.n16288 0.474
R54915 vdd.n16303 vdd.n16302 0.474
R54916 vdd.n16329 vdd.n16311 0.474
R54917 vdd.n16313 vdd.n16312 0.474
R54918 vdd.n16544 vdd.n16543 0.474
R54919 vdd.n16580 vdd.n16579 0.474
R54920 vdd.n16746 vdd.n16745 0.474
R54921 vdd.n16750 vdd.n16747 0.474
R54922 vdd.n16716 vdd.n16711 0.474
R54923 vdd.n16965 vdd.n16956 0.474
R54924 vdd.n16993 vdd.n16984 0.474
R54925 vdd.n17107 vdd.n17106 0.474
R54926 vdd.n17142 vdd.n17130 0.474
R54927 vdd.n17237 vdd.n17228 0.474
R54928 vdd.n17265 vdd.n17256 0.474
R54929 vdd.n17379 vdd.n17378 0.474
R54930 vdd.n17414 vdd.n17402 0.474
R54931 vdd.n17509 vdd.n17500 0.474
R54932 vdd.n17537 vdd.n17528 0.474
R54933 vdd.n17637 vdd.n17636 0.474
R54934 vdd.n17672 vdd.n17660 0.474
R54935 vdd.n17767 vdd.n17758 0.474
R54936 vdd.n17795 vdd.n17786 0.474
R54937 vdd.n17908 vdd.n17907 0.474
R54938 vdd.n17943 vdd.n17931 0.474
R54939 vdd.n18038 vdd.n18029 0.474
R54940 vdd.n18066 vdd.n18057 0.474
R54941 vdd.n18180 vdd.n18179 0.474
R54942 vdd.n18215 vdd.n18203 0.474
R54943 vdd.n18304 vdd.n18296 0.474
R54944 vdd.n15036 vdd.n15028 0.474
R54945 vdd.n18347 vdd.n18346 0.474
R54946 vdd.n18375 vdd.n18374 0.474
R54947 vdd.n18399 vdd.n18395 0.474
R54948 vdd.n18402 vdd.n18401 0.474
R54949 vdd.n2706 vdd.n2705 0.472
R54950 vdd.n2164 vdd.n2163 0.472
R54951 vdd.n2569 vdd.n2568 0.472
R54952 vdd.n35675 vdd.n35674 0.472
R54953 vdd.n33101 vdd.n33100 0.472
R54954 vdd.n37400 vdd.n37399 0.472
R54955 vdd.n37595 vdd.n37594 0.472
R54956 vdd.n26148 vdd.n26147 0.472
R54957 vdd.n31957 vdd.n31956 0.472
R54958 vdd.n32313 vdd.n32312 0.472
R54959 vdd.n27780 vdd.n27779 0.472
R54960 vdd.n29698 vdd.n29697 0.472
R54961 vdd.n30319 vdd.n30318 0.472
R54962 vdd.n30322 vdd.n30321 0.472
R54963 vdd.n33090 vdd.n33089 0.471
R54964 vdd.n37045 vdd.n37044 0.471
R54965 vdd.n37431 vdd.n37430 0.471
R54966 vdd.n31662 vdd.n31661 0.471
R54967 vdd.n31502 vdd.n31501 0.471
R54968 vdd.n28021 vdd.n28020 0.471
R54969 vdd.n29772 vdd.n29771 0.471
R54970 vdd.n2708 vdd.n2707 0.471
R54971 vdd.n2166 vdd.n2165 0.471
R54972 vdd.n2571 vdd.n2570 0.471
R54973 vdd.n26150 vdd.n26149 0.471
R54974 vdd.n24963 vdd.n24960 0.471
R54975 vdd.n24925 vdd.n24922 0.471
R54976 vdd.n24541 vdd.n24538 0.471
R54977 vdd.n24890 vdd.n24887 0.469
R54978 vdd.n4000 vdd.n3735 0.468
R54979 vdd.n2656 vdd.n2580 0.468
R54980 vdd.n25253 vdd.n24882 0.465
R54981 vdd.n24816 vdd.n24815 0.448
R54982 vdd.n25097 vdd.n25096 0.448
R54983 vdd.n36030 vdd.n36029 0.447
R54984 vdd.n36044 vdd.n36043 0.447
R54985 vdd.n36261 vdd.n36260 0.447
R54986 vdd.n36275 vdd.n36274 0.447
R54987 vdd.n36492 vdd.n36491 0.447
R54988 vdd.n36506 vdd.n36505 0.447
R54989 vdd.n36723 vdd.n36722 0.447
R54990 vdd.n36737 vdd.n36736 0.447
R54991 vdd.n36954 vdd.n36953 0.447
R54992 vdd.n36968 vdd.n36967 0.447
R54993 vdd.n33146 vdd.n33145 0.447
R54994 vdd.n35640 vdd.n35639 0.447
R54995 vdd.n37322 vdd.n37321 0.447
R54996 vdd.n37352 vdd.n37351 0.447
R54997 vdd.n35667 vdd.n35666 0.447
R54998 vdd.n32829 vdd.n32828 0.447
R54999 vdd.n38023 vdd.n38022 0.447
R55000 vdd.n38009 vdd.n38008 0.447
R55001 vdd.n37792 vdd.n37791 0.447
R55002 vdd.n37778 vdd.n37777 0.447
R55003 vdd.n28220 vdd.n28219 0.447
R55004 vdd.n28234 vdd.n28233 0.447
R55005 vdd.n28451 vdd.n28450 0.447
R55006 vdd.n28465 vdd.n28464 0.447
R55007 vdd.n28682 vdd.n28681 0.447
R55008 vdd.n28696 vdd.n28695 0.447
R55009 vdd.n26701 vdd.n26697 0.447
R55010 vdd.n26310 vdd.n26306 0.447
R55011 vdd.n27984 vdd.n27983 0.447
R55012 vdd.n27881 vdd.n27880 0.447
R55013 vdd.n31460 vdd.n31456 0.447
R55014 vdd.n32403 vdd.n32399 0.447
R55015 vdd.n31158 vdd.n31150 0.446
R55016 vdd.n3695 vdd.n2696 0.437
R55017 vdd.n3729 vdd.n3724 0.437
R55018 vdd.n2253 vdd.n2187 0.437
R55019 vdd.n2268 vdd.n2147 0.437
R55020 vdd.n2128 vdd.n2127 0.437
R55021 vdd.n2611 vdd.n2592 0.437
R55022 vdd.n1861 vdd.n1859 0.437
R55023 vdd.n1805 vdd.n1804 0.437
R55024 vdd.n27237 vdd.n27233 0.435
R55025 vdd.n24949 vdd.n24948 0.428
R55026 vdd.n1237 vdd.n1236 0.426
R55027 vdd.n1869 vdd.n1868 0.426
R55028 vdd.n1221 vdd.n1220 0.426
R55029 vdd.n2421 vdd.n2420 0.426
R55030 vdd.n3854 vdd.n3850 0.426
R55031 vdd.n3785 vdd.n3784 0.426
R55032 vdd.n10249 vdd.n10133 0.425
R55033 vdd.n27307 vdd.n27306 0.424
R55034 vdd.n25759 vdd.n25758 0.424
R55035 vdd.n3821 vdd.n3815 0.408
R55036 vdd.n2528 vdd.n2526 0.408
R55037 vdd.n1242 vdd.n1241 0.408
R55038 vdd.n2691 vdd.n2686 0.406
R55039 vdd.n2260 vdd.n2168 0.406
R55040 vdd.n2162 vdd.n2149 0.406
R55041 vdd.n1882 vdd.n1880 0.406
R55042 vdd.n2322 vdd.n2116 0.405
R55043 vdd.n12600 vdd.n10084 0.405
R55044 vdd.n33370 vdd.n33369 0.376
R55045 vdd.n33883 vdd.n33882 0.376
R55046 vdd.n33955 vdd.n33954 0.376
R55047 vdd.n35108 vdd.n35107 0.376
R55048 vdd.n35041 vdd.n35040 0.376
R55049 vdd.n34521 vdd.n34520 0.376
R55050 vdd.n34457 vdd.n34456 0.376
R55051 vdd.n592 vdd.n591 0.376
R55052 vdd.n261 vdd.n260 0.376
R55053 vdd.n270 vdd.n269 0.376
R55054 vdd.n23 vdd.n22 0.376
R55055 vdd.n35 vdd.n34 0.376
R55056 vdd.n580 vdd.n579 0.376
R55057 vdd.n6157 vdd.n6156 0.376
R55058 vdd.n6239 vdd.n6238 0.376
R55059 vdd.n5268 vdd.n5267 0.376
R55060 vdd.n5204 vdd.n5203 0.376
R55061 vdd.n5045 vdd.n5044 0.376
R55062 vdd.n4966 vdd.n4965 0.376
R55063 vdd.n4842 vdd.n4841 0.376
R55064 vdd.n4832 vdd.n4831 0.376
R55065 vdd.n4098 vdd.n4097 0.376
R55066 vdd.n4034 vdd.n4033 0.376
R55067 vdd.n30246 vdd.n30244 0.376
R55068 vdd.n31541 vdd.n31540 0.376
R55069 vdd.n31550 vdd.n31549 0.376
R55070 vdd.n31921 vdd.n31920 0.376
R55071 vdd.n31029 vdd.n31028 0.376
R55072 vdd.n31283 vdd.n31282 0.376
R55073 vdd.n30292 vdd.n30291 0.376
R55074 vdd.n35906 vdd.n35905 0.376
R55075 vdd.n35926 vdd.n35925 0.376
R55076 vdd.n36137 vdd.n36136 0.376
R55077 vdd.n36157 vdd.n36156 0.376
R55078 vdd.n36368 vdd.n36367 0.376
R55079 vdd.n36388 vdd.n36387 0.376
R55080 vdd.n36599 vdd.n36598 0.376
R55081 vdd.n36619 vdd.n36618 0.376
R55082 vdd.n36830 vdd.n36829 0.376
R55083 vdd.n36850 vdd.n36849 0.376
R55084 vdd.n33261 vdd.n33260 0.376
R55085 vdd.n33242 vdd.n33241 0.376
R55086 vdd.n33067 vdd.n33066 0.376
R55087 vdd.n37252 vdd.n37251 0.376
R55088 vdd.n37438 vdd.n37437 0.376
R55089 vdd.n32907 vdd.n32906 0.376
R55090 vdd.n38118 vdd.n38117 0.376
R55091 vdd.n38128 vdd.n38127 0.376
R55092 vdd.n37905 vdd.n37904 0.376
R55093 vdd.n37885 vdd.n37884 0.376
R55094 vdd.n37674 vdd.n37673 0.376
R55095 vdd.n37654 vdd.n37653 0.376
R55096 vdd.n28327 vdd.n28326 0.376
R55097 vdd.n28347 vdd.n28346 0.376
R55098 vdd.n28558 vdd.n28557 0.376
R55099 vdd.n28578 vdd.n28577 0.376
R55100 vdd.n28789 vdd.n28788 0.376
R55101 vdd.n28145 vdd.n28144 0.376
R55102 vdd.n28181 vdd.n28179 0.376
R55103 vdd.n27752 vdd.n27750 0.376
R55104 vdd.n27760 vdd.n27759 0.376
R55105 vdd.n29019 vdd.n29018 0.376
R55106 vdd.n29860 vdd.n29858 0.376
R55107 vdd.n29851 vdd.n29850 0.376
R55108 vdd.n29686 vdd.n29685 0.376
R55109 vdd.n27646 vdd.n27645 0.376
R55110 vdd.n27566 vdd.n27565 0.376
R55111 vdd.n27578 vdd.n27577 0.376
R55112 vdd.n26068 vdd.n26067 0.376
R55113 vdd.n25702 vdd.n25701 0.376
R55114 vdd.n25691 vdd.n25690 0.376
R55115 vdd.n25511 vdd.n25510 0.376
R55116 vdd.n25596 vdd.n25595 0.376
R55117 vdd.n25413 vdd.n25412 0.376
R55118 vdd.n27211 vdd.n27210 0.376
R55119 vdd.n1735 vdd.n1734 0.376
R55120 vdd.n1742 vdd.n1741 0.376
R55121 vdd.n1568 vdd.n1567 0.376
R55122 vdd.n1551 vdd.n1550 0.376
R55123 vdd.n1387 vdd.n1386 0.376
R55124 vdd.n1370 vdd.n1369 0.376
R55125 vdd.n26836 vdd.n26835 0.376
R55126 vdd.n26853 vdd.n26852 0.376
R55127 vdd.n27017 vdd.n27016 0.376
R55128 vdd.n27034 vdd.n27033 0.376
R55129 vdd.n27198 vdd.n27197 0.376
R55130 vdd.n26741 vdd.n26740 0.376
R55131 vdd.n1879 vdd.n1878 0.376
R55132 vdd.n1871 vdd.n1870 0.376
R55133 vdd.n1179 vdd.n1176 0.376
R55134 vdd.n2065 vdd.n2064 0.376
R55135 vdd.n1975 vdd.n1974 0.376
R55136 vdd.n2445 vdd.n2444 0.376
R55137 vdd.n2532 vdd.n2531 0.376
R55138 vdd.n2405 vdd.n2404 0.376
R55139 vdd.n2397 vdd.n2396 0.376
R55140 vdd.n2383 vdd.n2382 0.376
R55141 vdd.n2406 vdd.n2405 0.376
R55142 vdd.n2385 vdd.n2384 0.376
R55143 vdd.n2123 vdd.n2122 0.376
R55144 vdd.n2115 vdd.n2111 0.376
R55145 vdd.n2140 vdd.n2139 0.376
R55146 vdd.n2161 vdd.n2159 0.376
R55147 vdd.n2138 vdd.n2137 0.376
R55148 vdd.n2183 vdd.n2180 0.376
R55149 vdd.n2200 vdd.n2197 0.376
R55150 vdd.n3828 vdd.n3827 0.376
R55151 vdd.n3759 vdd.n3755 0.376
R55152 vdd.n3726 vdd.n3725 0.376
R55153 vdd.n2688 vdd.n2687 0.376
R55154 vdd.n2789 vdd.n2788 0.376
R55155 vdd.n2806 vdd.n2805 0.376
R55156 vdd.n2970 vdd.n2969 0.376
R55157 vdd.n2987 vdd.n2986 0.376
R55158 vdd.n3151 vdd.n3150 0.376
R55159 vdd.n3168 vdd.n3167 0.376
R55160 vdd.n3332 vdd.n3331 0.376
R55161 vdd.n3349 vdd.n3348 0.376
R55162 vdd.n3513 vdd.n3512 0.376
R55163 vdd.n3530 vdd.n3529 0.376
R55164 vdd.n31757 vdd.n31747 0.376
R55165 vdd.n31737 vdd.n31736 0.376
R55166 vdd.n31681 vdd.n31680 0.376
R55167 vdd.n31883 vdd.n31882 0.376
R55168 vdd.n13214 vdd.n9204 0.376
R55169 vdd.n13248 vdd.n9175 0.376
R55170 vdd.n13507 vdd.n8983 0.376
R55171 vdd.n13540 vdd.n8955 0.376
R55172 vdd.n13789 vdd.n13788 0.376
R55173 vdd.n13825 vdd.n8736 0.376
R55174 vdd.n14116 vdd.n8515 0.376
R55175 vdd.n8521 vdd.n8507 0.376
R55176 vdd.n14398 vdd.n8301 0.376
R55177 vdd.n14428 vdd.n14427 0.376
R55178 vdd.n14785 vdd.n8076 0.376
R55179 vdd.n8078 vdd.n8077 0.376
R55180 vdd.n13143 vdd.n13142 0.376
R55181 vdd.n13381 vdd.n9060 0.376
R55182 vdd.n13436 vdd.n13435 0.376
R55183 vdd.n13673 vdd.n8840 0.376
R55184 vdd.n13728 vdd.n13727 0.376
R55185 vdd.n13953 vdd.n13952 0.376
R55186 vdd.n13996 vdd.n13995 0.376
R55187 vdd.n14243 vdd.n14242 0.376
R55188 vdd.n14287 vdd.n14286 0.376
R55189 vdd.n14541 vdd.n8179 0.376
R55190 vdd.n14612 vdd.n14611 0.376
R55191 vdd.n11626 vdd.n11579 0.376
R55192 vdd.n22152 vdd.n22144 0.376
R55193 vdd.n22163 vdd.n22156 0.376
R55194 vdd.n24201 vdd.n24194 0.376
R55195 vdd.n23979 vdd.n23972 0.376
R55196 vdd.n23969 vdd.n23962 0.376
R55197 vdd.n23747 vdd.n23740 0.376
R55198 vdd.n23737 vdd.n23730 0.376
R55199 vdd.n23059 vdd.n23052 0.376
R55200 vdd.n23281 vdd.n23274 0.376
R55201 vdd.n23291 vdd.n23284 0.376
R55202 vdd.n23513 vdd.n23506 0.376
R55203 vdd.n23523 vdd.n23516 0.376
R55204 vdd.n22480 vdd.n22473 0.376
R55205 vdd.n22702 vdd.n22695 0.376
R55206 vdd.n22712 vdd.n22705 0.376
R55207 vdd.n22934 vdd.n22927 0.376
R55208 vdd.n22944 vdd.n22937 0.376
R55209 vdd.n22184 vdd.n22177 0.376
R55210 vdd.n22267 vdd.n22259 0.376
R55211 vdd.n22278 vdd.n22271 0.376
R55212 vdd.n19408 vdd.n19407 0.376
R55213 vdd.n19425 vdd.n19424 0.376
R55214 vdd.n19611 vdd.n19610 0.376
R55215 vdd.n19628 vdd.n19627 0.376
R55216 vdd.n19813 vdd.n19812 0.376
R55217 vdd.n19163 vdd.n19162 0.376
R55218 vdd.n20833 vdd.n20832 0.376
R55219 vdd.n20819 vdd.n20818 0.376
R55220 vdd.n20631 vdd.n20630 0.376
R55221 vdd.n20617 vdd.n20616 0.376
R55222 vdd.n21655 vdd.n21654 0.376
R55223 vdd.n21388 vdd.n21387 0.376
R55224 vdd.n21374 vdd.n21373 0.376
R55225 vdd.n21129 vdd.n21128 0.376
R55226 vdd.n21115 vdd.n21114 0.376
R55227 vdd.n19022 vdd.n19021 0.376
R55228 vdd.n19008 vdd.n19007 0.376
R55229 vdd.n18763 vdd.n18762 0.376
R55230 vdd.n18749 vdd.n18748 0.376
R55231 vdd.n18504 vdd.n18503 0.376
R55232 vdd.n18463 vdd.n18462 0.376
R55233 vdd.n21632 vdd.n21631 0.376
R55234 vdd.n20000 vdd.n19991 0.376
R55235 vdd.n20012 vdd.n20003 0.376
R55236 vdd.n24514 vdd.n24410 0.376
R55237 vdd.n24983 vdd.n24978 0.376
R55238 vdd.n2260 vdd.n2169 0.375
R55239 vdd.n2631 vdd.n2589 0.375
R55240 vdd.n2660 vdd.n2578 0.375
R55241 vdd.n1786 vdd.n1785 0.375
R55242 vdd.n1236 vdd.n1234 0.375
R55243 vdd.n10094 vdd.n10083 0.375
R55244 vdd.n1950 vdd.n1934 0.374
R55245 vdd.n33576 vdd.n33575 0.373
R55246 vdd.n1052 vdd.n1051 0.373
R55247 vdd.n1181 vdd.n1180 0.373
R55248 vdd.n2025 vdd.n2024 0.373
R55249 vdd.n1835 vdd.n1833 0.373
R55250 vdd.n25256 vdd.n24408 0.371
R55251 vdd.n34241 vdd.n34240 0.362
R55252 vdd.n35468 vdd.n35467 0.362
R55253 vdd.n34883 vdd.n34882 0.362
R55254 vdd.n5926 vdd.n5925 0.362
R55255 vdd.n5630 vdd.n5629 0.362
R55256 vdd.n4457 vdd.n4456 0.362
R55257 vdd.n33149 vdd.n33148 0.362
R55258 vdd.n35643 vdd.n35642 0.362
R55259 vdd.n37325 vdd.n37324 0.362
R55260 vdd.n37355 vdd.n37354 0.362
R55261 vdd.n35670 vdd.n35669 0.362
R55262 vdd.n32832 vdd.n32831 0.362
R55263 vdd.n8444 vdd.n8402 0.362
R55264 vdd.n8667 vdd.n8624 0.362
R55265 vdd.n13648 vdd.n8845 0.362
R55266 vdd.n13356 vdd.n9065 0.362
R55267 vdd.n13401 vdd.n13400 0.362
R55268 vdd.n13694 vdd.n13693 0.362
R55269 vdd.n8613 vdd.n8609 0.362
R55270 vdd.n8391 vdd.n8387 0.362
R55271 vdd.n19270 vdd.n19269 0.362
R55272 vdd.n19258 vdd.n19257 0.362
R55273 vdd.n19214 vdd.n19213 0.362
R55274 vdd.n19202 vdd.n19201 0.362
R55275 vdd.n19856 vdd.n19855 0.362
R55276 vdd.n19868 vdd.n19867 0.362
R55277 vdd.n19924 vdd.n19923 0.362
R55278 vdd.n19936 vdd.n19935 0.362
R55279 vdd.n4619 vdd.n4618 0.362
R55280 vdd.n27287 vdd.n27286 0.362
R55281 vdd.n25733 vdd.n25732 0.362
R55282 vdd.n23060 vdd.n23050 0.354
R55283 vdd.n23628 vdd.n23626 0.353
R55284 vdd.n33291 vdd.n33290 0.351
R55285 vdd.n601 vdd.n600 0.351
R55286 vdd.n509 vdd.n508 0.351
R55287 vdd.n3901 vdd.n3900 0.349
R55288 vdd.n24523 vdd.n24522 0.348
R55289 vdd.n2046 vdd.n2045 0.347
R55290 vdd.n3695 vdd.n2694 0.343
R55291 vdd.n3982 vdd.n3760 0.343
R55292 vdd.n2253 vdd.n2186 0.343
R55293 vdd.n2611 vdd.n2591 0.343
R55294 vdd.n2660 vdd.n2576 0.343
R55295 vdd.n1805 vdd.n1803 0.343
R55296 vdd.n10246 vdd.n10072 0.343
R55297 vdd.n33855 vdd.n33854 0.34
R55298 vdd.n955 vdd.n954 0.34
R55299 vdd.n386 vdd.n385 0.327
R55300 vdd.n32241 vdd.n32240 0.325
R55301 vdd.n3807 vdd.n3805 0.323
R55302 vdd.n10388 vdd.n10387 0.32
R55303 vdd.n10380 vdd.n10379 0.32
R55304 vdd.n13059 vdd.t212 0.32
R55305 vdd.n9440 vdd.n9439 0.32
R55306 vdd.n12987 vdd.n9415 0.32
R55307 vdd.n12889 vdd.n12888 0.32
R55308 vdd.n12881 vdd.n12880 0.32
R55309 vdd.n9799 vdd.n9798 0.32
R55310 vdd.n12779 vdd.n9776 0.32
R55311 vdd.n9813 vdd.t387 0.32
R55312 vdd.n12681 vdd.n12680 0.32
R55313 vdd.n12673 vdd.n12672 0.32
R55314 vdd.n10242 vdd.n10241 0.32
R55315 vdd.n10484 vdd.n10119 0.32
R55316 vdd.n10665 vdd.n10656 0.32
R55317 vdd.n10690 vdd.n10689 0.32
R55318 vdd.n10845 vdd.n10844 0.32
R55319 vdd.n10861 vdd.n10860 0.32
R55320 vdd.n12241 vdd.n12240 0.32
R55321 vdd.n12234 vdd.n11012 0.32
R55322 vdd.n12134 vdd.n12133 0.32
R55323 vdd.n12121 vdd.n11185 0.32
R55324 vdd.n12072 vdd.t302 0.32
R55325 vdd.n11354 vdd.n11353 0.32
R55326 vdd.n11370 vdd.n11369 0.32
R55327 vdd.n15252 vdd.n15251 0.32
R55328 vdd.n15241 vdd.n15240 0.32
R55329 vdd.n15495 vdd.t181 0.32
R55330 vdd.n15230 vdd.n15229 0.32
R55331 vdd.n15216 vdd.n15215 0.32
R55332 vdd.n15202 vdd.n15201 0.32
R55333 vdd.n15195 vdd.n15194 0.32
R55334 vdd.n15174 vdd.n15173 0.32
R55335 vdd.n15160 vdd.n15159 0.32
R55336 vdd.n16192 vdd.t2 0.32
R55337 vdd.n15146 vdd.n15145 0.32
R55338 vdd.n15132 vdd.n15131 0.32
R55339 vdd.n16664 vdd.n16663 0.32
R55340 vdd.n16657 vdd.n16656 0.32
R55341 vdd.n17102 vdd.n17099 0.32
R55342 vdd.n17122 vdd.n17119 0.32
R55343 vdd.n17374 vdd.n17371 0.32
R55344 vdd.n17394 vdd.n17391 0.32
R55345 vdd.n17632 vdd.n17629 0.32
R55346 vdd.n17652 vdd.n17649 0.32
R55347 vdd.n17903 vdd.n17900 0.32
R55348 vdd.n17923 vdd.n17920 0.32
R55349 vdd.t264 vdd.n18060 0.32
R55350 vdd.n18175 vdd.n18172 0.32
R55351 vdd.n18195 vdd.n18192 0.32
R55352 vdd.n11628 vdd.n11567 0.319
R55353 vdd.n13145 vdd.n9245 0.319
R55354 vdd.t324 vdd.n9213 0.319
R55355 vdd.n13204 vdd.t320 0.319
R55356 vdd.n13216 vdd.n9191 0.319
R55357 vdd.n25629 vdd.n25628 0.318
R55358 vdd.n1923 vdd.n1204 0.312
R55359 vdd.n31120 vdd.n31033 0.312
R55360 vdd.n32232 vdd.n31554 0.312
R55361 vdd.n32259 vdd.n31543 0.312
R55362 vdd.n3680 vdd.n2727 0.312
R55363 vdd.n4000 vdd.n3738 0.312
R55364 vdd.n2128 vdd.n2126 0.312
R55365 vdd.n2645 vdd.n2583 0.312
R55366 vdd.n3820 vdd.n3818 0.312
R55367 vdd.n10142 vdd.n10084 0.312
R55368 vdd.n16705 vdd.n16704 0.312
R55369 vdd.n13257 vdd.n9170 0.305
R55370 vdd.n13246 vdd.n9178 0.305
R55371 vdd.t289 vdd.n9179 0.305
R55372 vdd.n13378 vdd.n9045 0.305
R55373 vdd.n13389 vdd.n9055 0.305
R55374 vdd.n13438 vdd.n9021 0.305
R55375 vdd.n13509 vdd.n8981 0.305
R55376 vdd.n13548 vdd.n8950 0.305
R55377 vdd.n13538 vdd.n8957 0.305
R55378 vdd.n13670 vdd.n8824 0.305
R55379 vdd.n13681 vdd.n8835 0.305
R55380 vdd.n13730 vdd.n8801 0.305
R55381 vdd.n13745 vdd.t288 0.305
R55382 vdd.n13791 vdd.n8766 0.305
R55383 vdd.n13833 vdd.n8731 0.305
R55384 vdd.n13823 vdd.n13821 0.305
R55385 vdd.n8632 vdd.n8614 0.305
R55386 vdd.n14004 vdd.n8593 0.305
R55387 vdd.n13993 vdd.n13992 0.305
R55388 vdd.n14118 vdd.n8512 0.305
R55389 vdd.n8536 vdd.n8524 0.305
R55390 vdd.n14127 vdd.n14125 0.305
R55391 vdd.t132 vdd.n8497 0.305
R55392 vdd.n8410 vdd.n8392 0.305
R55393 vdd.n14295 vdd.n8371 0.305
R55394 vdd.n14284 vdd.n14283 0.305
R55395 vdd.n14396 vdd.n8303 0.305
R55396 vdd.n14407 vdd.n14406 0.305
R55397 vdd.n14430 vdd.n8274 0.305
R55398 vdd.n14439 vdd.t318 0.305
R55399 vdd.n14452 vdd.t318 0.305
R55400 vdd.n14566 vdd.n8183 0.305
R55401 vdd.n14614 vdd.n8174 0.305
R55402 vdd.n12600 vdd.n10074 0.303
R55403 vdd.n31187 vdd.n31025 0.3
R55404 vdd.n10261 vdd.n10123 0.297
R55405 vdd.n1188 vdd.n1187 0.293
R55406 vdd.n2032 vdd.n2031 0.293
R55407 vdd.n2020 vdd.n2019 0.293
R55408 vdd.n11767 vdd.n11766 0.29
R55409 vdd.n32245 vdd.n31546 0.287
R55410 vdd.n25449 vdd.n25448 0.283
R55411 vdd.n11666 vdd.n11664 0.282
R55412 vdd.n11872 vdd.n11806 0.282
R55413 vdd.n21963 vdd.n21897 0.282
R55414 vdd.n3683 vdd.n2710 0.281
R55415 vdd.n2248 vdd.n2205 0.281
R55416 vdd.n2268 vdd.n2145 0.281
R55417 vdd.n2141 vdd.n2136 0.281
R55418 vdd.n2467 vdd.n2464 0.281
R55419 vdd.n1882 vdd.n1876 0.281
R55420 vdd.n1827 vdd.n1254 0.281
R55421 vdd.n3997 vdd.n3745 0.28
R55422 vdd.n2061 vdd.n2060 0.279
R55423 vdd.n24828 vdd.n24827 0.274
R55424 vdd.n12600 vdd.n10083 0.265
R55425 vdd.n16743 vdd.n16718 0.265
R55426 vdd.n31187 vdd.n31022 0.262
R55427 vdd.n11763 vdd.n11679 0.262
R55428 vdd.n4829 vdd.n4828 0.261
R55429 vdd.n25494 vdd.n25493 0.261
R55430 vdd.n11791 vdd.n11789 0.261
R55431 vdd.n21882 vdd.n21880 0.261
R55432 vdd.n31775 vdd.n31770 0.26
R55433 vdd.n31775 vdd.n31774 0.26
R55434 vdd.n25259 vdd.n25258 0.256
R55435 vdd.n11768 vdd.n11668 0.251
R55436 vdd.n32210 vdd.n32207 0.25
R55437 vdd.n3985 vdd.n3753 0.25
R55438 vdd.n1870 vdd.n1869 0.25
R55439 vdd.n33740 vdd.n33739 0.25
R55440 vdd.n920 vdd.n919 0.25
R55441 vdd.n1912 vdd.n1911 0.249
R55442 vdd.n3692 vdd.n2704 0.249
R55443 vdd.n2250 vdd.n2201 0.249
R55444 vdd.n2387 vdd.n2386 0.249
R55445 vdd.n28118 vdd.n28115 0.247
R55446 vdd.n27841 vdd.n27839 0.247
R55447 vdd.n29822 vdd.n29819 0.247
R55448 vdd.n22153 vdd.n22152 0.247
R55449 vdd.n22164 vdd.n22163 0.247
R55450 vdd.n22185 vdd.n22184 0.247
R55451 vdd.n22268 vdd.n22267 0.247
R55452 vdd.n22279 vdd.n22278 0.247
R55453 vdd.n25255 vdd.n25254 0.247
R55454 vdd.n10246 vdd.n10122 0.237
R55455 vdd.n10385 vdd.n10341 0.237
R55456 vdd.n10377 vdd.n10342 0.237
R55457 vdd.n9437 vdd.n9436 0.237
R55458 vdd.n12990 vdd.n12989 0.237
R55459 vdd.n12891 vdd.n9605 0.237
R55460 vdd.n12883 vdd.n9612 0.237
R55461 vdd.n9796 vdd.n9795 0.237
R55462 vdd.n12782 vdd.n12781 0.237
R55463 vdd.n12683 vdd.n9965 0.237
R55464 vdd.n12675 vdd.n9972 0.237
R55465 vdd.n10600 vdd.n10590 0.237
R55466 vdd.n12479 vdd.n10588 0.237
R55467 vdd.n10661 vdd.n10660 0.237
R55468 vdd.n10692 vdd.n10678 0.237
R55469 vdd.n12378 vdd.n10751 0.237
R55470 vdd.n12374 vdd.n10754 0.237
R55471 vdd.n10847 vdd.n10831 0.237
R55472 vdd.n10858 vdd.n10853 0.237
R55473 vdd.n10943 vdd.n10919 0.237
R55474 vdd.n10947 vdd.n10920 0.237
R55475 vdd.n11021 vdd.n11019 0.237
R55476 vdd.n12232 vdd.n12231 0.237
R55477 vdd.n12182 vdd.n12181 0.237
R55478 vdd.n11122 vdd.n11121 0.237
R55479 vdd.n12136 vdd.n11176 0.237
R55480 vdd.n11202 vdd.n11182 0.237
R55481 vdd.n12076 vdd.n11245 0.237
R55482 vdd.n12068 vdd.n11271 0.237
R55483 vdd.n11356 vdd.n11340 0.237
R55484 vdd.n11367 vdd.n11362 0.237
R55485 vdd.n16669 vdd.n16647 0.237
R55486 vdd.n15254 vdd.n15247 0.237
R55487 vdd.n15243 vdd.n15236 0.237
R55488 vdd.n15232 vdd.n15222 0.237
R55489 vdd.n15218 vdd.n15208 0.237
R55490 vdd.n15204 vdd.n15182 0.237
R55491 vdd.n15192 vdd.n15191 0.237
R55492 vdd.n15176 vdd.n15166 0.237
R55493 vdd.n15162 vdd.n15152 0.237
R55494 vdd.n15148 vdd.n15138 0.237
R55495 vdd.n15134 vdd.n15124 0.237
R55496 vdd.n16979 vdd.n16978 0.237
R55497 vdd.n16995 vdd.n16993 0.237
R55498 vdd.n17096 vdd.n17095 0.237
R55499 vdd.n17112 vdd.n17111 0.237
R55500 vdd.n17251 vdd.n17250 0.237
R55501 vdd.n17267 vdd.n17265 0.237
R55502 vdd.n17368 vdd.n17367 0.237
R55503 vdd.n17384 vdd.n17383 0.237
R55504 vdd.n17523 vdd.n17522 0.237
R55505 vdd.n17539 vdd.n17537 0.237
R55506 vdd.n17626 vdd.n17625 0.237
R55507 vdd.n17642 vdd.n17641 0.237
R55508 vdd.n17781 vdd.n17780 0.237
R55509 vdd.n17797 vdd.n17795 0.237
R55510 vdd.n17897 vdd.n17896 0.237
R55511 vdd.n17913 vdd.n17912 0.237
R55512 vdd.n18052 vdd.n18051 0.237
R55513 vdd.n18068 vdd.n18066 0.237
R55514 vdd.n18169 vdd.n18168 0.237
R55515 vdd.n18185 vdd.n18184 0.237
R55516 vdd.n12600 vdd.n10073 0.236
R55517 vdd.n2623 vdd.n2617 0.233
R55518 vdd.n2623 vdd.n2619 0.233
R55519 vdd.n2240 vdd.n2234 0.233
R55520 vdd.n2240 vdd.n2236 0.233
R55521 vdd.n3954 vdd.n3949 0.233
R55522 vdd.n3954 vdd.n3950 0.233
R55523 vdd.n11871 vdd.n11870 0.233
R55524 vdd.n21962 vdd.n21961 0.233
R55525 vdd.n11818 vdd.n11808 0.233
R55526 vdd.n21909 vdd.n21899 0.233
R55527 vdd.n11758 vdd.n11757 0.23
R55528 vdd.n21838 vdd.n21837 0.23
R55529 vdd.n31075 vdd.n31074 0.225
R55530 vdd.n35910 vdd.n35909 0.223
R55531 vdd.n35931 vdd.n35930 0.223
R55532 vdd.n36141 vdd.n36140 0.223
R55533 vdd.n36162 vdd.n36161 0.223
R55534 vdd.n36372 vdd.n36371 0.223
R55535 vdd.n36393 vdd.n36392 0.223
R55536 vdd.n36603 vdd.n36602 0.223
R55537 vdd.n36624 vdd.n36623 0.223
R55538 vdd.n36834 vdd.n36833 0.223
R55539 vdd.n36855 vdd.n36854 0.223
R55540 vdd.n33265 vdd.n33264 0.223
R55541 vdd.n33247 vdd.n33246 0.223
R55542 vdd.n33071 vdd.n33070 0.223
R55543 vdd.n37257 vdd.n37256 0.223
R55544 vdd.n37442 vdd.n37441 0.223
R55545 vdd.n32911 vdd.n32910 0.223
R55546 vdd.n38122 vdd.n38121 0.223
R55547 vdd.n38133 vdd.n38132 0.223
R55548 vdd.n37909 vdd.n37908 0.223
R55549 vdd.n37889 vdd.n37888 0.223
R55550 vdd.n37678 vdd.n37677 0.223
R55551 vdd.n37658 vdd.n37657 0.223
R55552 vdd.n28331 vdd.n28330 0.223
R55553 vdd.n28352 vdd.n28351 0.223
R55554 vdd.n28562 vdd.n28561 0.223
R55555 vdd.n28583 vdd.n28582 0.223
R55556 vdd.n28793 vdd.n28792 0.223
R55557 vdd.n28150 vdd.n28149 0.223
R55558 vdd.n27764 vdd.n27763 0.223
R55559 vdd.n31887 vdd.n31886 0.223
R55560 vdd.n32225 vdd.n32224 0.223
R55561 vdd.n29691 vdd.n29690 0.223
R55562 vdd.n30296 vdd.n30295 0.223
R55563 vdd.n30565 vdd.n30564 0.223
R55564 vdd.n6363 vdd 0.219
R55565 vdd.n1923 vdd.n1189 0.218
R55566 vdd.n2228 vdd.n2209 0.218
R55567 vdd.n2484 vdd.n2453 0.218
R55568 vdd.n24970 vdd.n24957 0.215
R55569 vdd.n32004 vdd.n31618 0.212
R55570 vdd.n32331 vdd.n31491 0.212
R55571 vdd.n26178 vdd.n26165 0.212
R55572 vdd.n3902 vdd.n3901 0.209
R55573 vdd.n3902 vdd.n3898 0.209
R55574 vdd.n11891 vdd.n11798 0.206
R55575 vdd.n21982 vdd.n21889 0.206
R55576 vdd.n25397 vdd.n25396 0.206
R55577 vdd.n11727 vdd.n11722 0.204
R55578 vdd.n11896 vdd.n11795 0.202
R55579 vdd.n21987 vdd.n21886 0.202
R55580 vdd.n31104 vdd.n31100 0.2
R55581 vdd.n24557 vdd.n24534 0.195
R55582 vdd.n27224 vdd.n27223 0.193
R55583 vdd.n27219 vdd.n27218 0.193
R55584 vdd.n2802 vdd.n2798 0.19
R55585 vdd.n2891 vdd.n2888 0.19
R55586 vdd.n2898 vdd.n2891 0.19
R55587 vdd.n2983 vdd.n2979 0.19
R55588 vdd.n3072 vdd.n3069 0.19
R55589 vdd.n3079 vdd.n3072 0.19
R55590 vdd.n3164 vdd.n3160 0.19
R55591 vdd.n3253 vdd.n3250 0.19
R55592 vdd.n3260 vdd.n3253 0.19
R55593 vdd.n3345 vdd.n3341 0.19
R55594 vdd.n3434 vdd.n3431 0.19
R55595 vdd.n3441 vdd.n3434 0.19
R55596 vdd.n3526 vdd.n3522 0.19
R55597 vdd.n3615 vdd.n3612 0.19
R55598 vdd.n3622 vdd.n3615 0.19
R55599 vdd.n35922 vdd.n35918 0.19
R55600 vdd.n36037 vdd.n36033 0.19
R55601 vdd.n36047 vdd.n36037 0.19
R55602 vdd.n36153 vdd.n36149 0.19
R55603 vdd.n36268 vdd.n36264 0.19
R55604 vdd.n36278 vdd.n36268 0.19
R55605 vdd.n36384 vdd.n36380 0.19
R55606 vdd.n36499 vdd.n36495 0.19
R55607 vdd.n36509 vdd.n36499 0.19
R55608 vdd.n36615 vdd.n36611 0.19
R55609 vdd.n36730 vdd.n36726 0.19
R55610 vdd.n36740 vdd.n36730 0.19
R55611 vdd.n36846 vdd.n36842 0.19
R55612 vdd.n36961 vdd.n36957 0.19
R55613 vdd.n36971 vdd.n36961 0.19
R55614 vdd.n38026 vdd.n38016 0.19
R55615 vdd.n38016 vdd.n38012 0.19
R55616 vdd.n37901 vdd.n37897 0.19
R55617 vdd.n37795 vdd.n37785 0.19
R55618 vdd.n37785 vdd.n37781 0.19
R55619 vdd.n37670 vdd.n37666 0.19
R55620 vdd.n28227 vdd.n28223 0.19
R55621 vdd.n28237 vdd.n28227 0.19
R55622 vdd.n28343 vdd.n28339 0.19
R55623 vdd.n28458 vdd.n28454 0.19
R55624 vdd.n28468 vdd.n28458 0.19
R55625 vdd.n28574 vdd.n28570 0.19
R55626 vdd.n28689 vdd.n28685 0.19
R55627 vdd.n28699 vdd.n28689 0.19
R55628 vdd.n1660 vdd.n1653 0.19
R55629 vdd.n1653 vdd.n1650 0.19
R55630 vdd.n1564 vdd.n1560 0.19
R55631 vdd.n1479 vdd.n1472 0.19
R55632 vdd.n1472 vdd.n1469 0.19
R55633 vdd.n1383 vdd.n1379 0.19
R55634 vdd.n1298 vdd.n1291 0.19
R55635 vdd.n26849 vdd.n26845 0.19
R55636 vdd.n26938 vdd.n26935 0.19
R55637 vdd.n26945 vdd.n26938 0.19
R55638 vdd.n27030 vdd.n27026 0.19
R55639 vdd.n27119 vdd.n27116 0.19
R55640 vdd.n27126 vdd.n27119 0.19
R55641 vdd.n11751 vdd.n11720 0.19
R55642 vdd.n25028 vdd.n25026 0.19
R55643 vdd.n25026 vdd.n25022 0.19
R55644 vdd.n24603 vdd.n24600 0.19
R55645 vdd.n24600 vdd.n24597 0.19
R55646 vdd.n3946 vdd.n3945 0.189
R55647 vdd.n3928 vdd.n3927 0.189
R55648 vdd.n2391 vdd.n2390 0.189
R55649 vdd.n2552 vdd.n2551 0.189
R55650 vdd.n1895 vdd.n1894 0.189
R55651 vdd.n1228 vdd.n1227 0.189
R55652 vdd.n3793 vdd.n3792 0.189
R55653 vdd.n2412 vdd.n2411 0.189
R55654 vdd.n1875 vdd.n1874 0.189
R55655 vdd.n33793 vdd.n33792 0.189
R55656 vdd.n34223 vdd.n34222 0.189
R55657 vdd.n35344 vdd.n35343 0.189
R55658 vdd.n34760 vdd.n34759 0.189
R55659 vdd.n308 vdd.n307 0.189
R55660 vdd.n200 vdd.n199 0.189
R55661 vdd.n5850 vdd.n5849 0.189
R55662 vdd.n5507 vdd.n5506 0.189
R55663 vdd.n4938 vdd.n4937 0.189
R55664 vdd.n4334 vdd.n4333 0.189
R55665 vdd.n37123 vdd.n37122 0.189
R55666 vdd.n33179 vdd.n33178 0.189
R55667 vdd.n33016 vdd.n33015 0.189
R55668 vdd.n37300 vdd.n37299 0.189
R55669 vdd.n37512 vdd.n37511 0.189
R55670 vdd.n32853 vdd.n32852 0.189
R55671 vdd.n37125 vdd.n37124 0.189
R55672 vdd.n33183 vdd.n33182 0.189
R55673 vdd.n33018 vdd.n33017 0.189
R55674 vdd.n37302 vdd.n37301 0.189
R55675 vdd.n37514 vdd.n37513 0.189
R55676 vdd.n32855 vdd.n32854 0.189
R55677 vdd.n26401 vdd.n26400 0.189
R55678 vdd.n31766 vdd.n31765 0.189
R55679 vdd.n32083 vdd.n32082 0.189
R55680 vdd.n32115 vdd.n32114 0.189
R55681 vdd.n32494 vdd.n32493 0.189
R55682 vdd.n32470 vdd.n32469 0.189
R55683 vdd.n31764 vdd.n31763 0.189
R55684 vdd.n32113 vdd.n32112 0.189
R55685 vdd.n32424 vdd.n32423 0.189
R55686 vdd.n28923 vdd.n28922 0.189
R55687 vdd.n28932 vdd.n28931 0.189
R55688 vdd.n27946 vdd.n27945 0.189
R55689 vdd.n27923 vdd.n27922 0.189
R55690 vdd.n30633 vdd.n30632 0.189
R55691 vdd.n30623 vdd.n30622 0.189
R55692 vdd.n28930 vdd.n28929 0.189
R55693 vdd.n27920 vdd.n27919 0.189
R55694 vdd.n30226 vdd.n30225 0.189
R55695 vdd.n25395 vdd.n25394 0.189
R55696 vdd.n25421 vdd.n25420 0.189
R55697 vdd.n28921 vdd.n28920 0.188
R55698 vdd.n27900 vdd.n27899 0.188
R55699 vdd.n30211 vdd.n30210 0.188
R55700 vdd.n27654 vdd.n27653 0.188
R55701 vdd.n26076 vdd.n26075 0.188
R55702 vdd.n25393 vdd.n25392 0.188
R55703 vdd.n3777 vdd.n3776 0.188
R55704 vdd.n2389 vdd.n2388 0.188
R55705 vdd.n1212 vdd.n1211 0.188
R55706 vdd.n26399 vdd.n26398 0.188
R55707 vdd.n32081 vdd.n32080 0.188
R55708 vdd.n32415 vdd.n32414 0.188
R55709 vdd.n31988 vdd.n31634 0.187
R55710 vdd.n32043 vdd.n32041 0.187
R55711 vdd.n32340 vdd.n32338 0.187
R55712 vdd.n3730 vdd.n3729 0.187
R55713 vdd.n3873 vdd.n3868 0.187
R55714 vdd.n2257 vdd.n2184 0.187
R55715 vdd.n2315 vdd.n2121 0.187
R55716 vdd.n2558 vdd.n2407 0.187
R55717 vdd.n2514 vdd.n2436 0.187
R55718 vdd.n2501 vdd.n2442 0.187
R55719 vdd.n1854 vdd.n1852 0.187
R55720 vdd.n1839 vdd.n1838 0.187
R55721 vdd.n26349 vdd.n26338 0.187
R55722 vdd.n24988 vdd.n24987 0.187
R55723 vdd.n33288 vdd.n33286 0.185
R55724 vdd.n34102 vdd.n34100 0.185
R55725 vdd.n35481 vdd.n35479 0.185
R55726 vdd.n34960 vdd.n34958 0.185
R55727 vdd.n598 vdd.n596 0.185
R55728 vdd.n506 vdd.n504 0.185
R55729 vdd.n5810 vdd.n5808 0.185
R55730 vdd.n5707 vdd.n5705 0.185
R55731 vdd.n4534 vdd.n4532 0.185
R55732 vdd.n31129 vdd.n31128 0.185
R55733 vdd.n27383 vdd.n27381 0.185
R55734 vdd.n25826 vdd.n25824 0.185
R55735 vdd.n25566 vdd.n25564 0.185
R55736 vdd.n28143 vdd.n28140 0.185
R55737 vdd.n29033 vdd.n29030 0.185
R55738 vdd.n27795 vdd.n27794 0.185
R55739 vdd.n29695 vdd.n29694 0.185
R55740 vdd.n8076 vdd.n8067 0.185
R55741 vdd.n8077 vdd.n8066 0.185
R55742 vdd.n20001 vdd.n20000 0.185
R55743 vdd.n20013 vdd.n20012 0.185
R55744 vdd.n24515 vdd.n24514 0.185
R55745 vdd.n24984 vdd.n24983 0.185
R55746 vdd.n3664 vdd.n3663 0.184
R55747 vdd.n3670 vdd.n3669 0.184
R55748 vdd.n11716 vdd.n11687 0.183
R55749 vdd.n11708 vdd.n11692 0.183
R55750 vdd.n11861 vdd.n11860 0.183
R55751 vdd.n11843 vdd.n11841 0.183
R55752 vdd.n21795 vdd.n21794 0.183
R55753 vdd.n21780 vdd.n21779 0.183
R55754 vdd.n21952 vdd.n21951 0.183
R55755 vdd.n21934 vdd.n21932 0.183
R55756 vdd.n3965 vdd.n3964 0.178
R55757 vdd.n3908 vdd.n3907 0.178
R55758 vdd.n2360 vdd.n2359 0.178
R55759 vdd.n2538 vdd.n2537 0.178
R55760 vdd.n1921 vdd.n1920 0.178
R55761 vdd.n1850 vdd.n1849 0.178
R55762 vdd.n3799 vdd.n3798 0.178
R55763 vdd.n2430 vdd.n2429 0.178
R55764 vdd.n1232 vdd.n1231 0.178
R55765 vdd.n33688 vdd.n33687 0.178
R55766 vdd.n1154 vdd.n1153 0.178
R55767 vdd.n188 vdd.n187 0.178
R55768 vdd.n5180 vdd.n5179 0.178
R55769 vdd.n37106 vdd.n37105 0.178
R55770 vdd.n37139 vdd.n37138 0.178
R55771 vdd.n37291 vdd.n37290 0.178
R55772 vdd.n33000 vdd.n32999 0.178
R55773 vdd.n32873 vdd.n32872 0.178
R55774 vdd.n37534 vdd.n37533 0.178
R55775 vdd.n26329 vdd.n26328 0.178
R55776 vdd.n31798 vdd.n31797 0.178
R55777 vdd.n31589 vdd.n31588 0.178
R55778 vdd.n32148 vdd.n32147 0.178
R55779 vdd.n32522 vdd.n32521 0.178
R55780 vdd.n32456 vdd.n32455 0.178
R55781 vdd.n31796 vdd.n31795 0.178
R55782 vdd.n32146 vdd.n32145 0.178
R55783 vdd.n32437 vdd.n32436 0.178
R55784 vdd.n28909 vdd.n28908 0.178
R55785 vdd.n28945 vdd.n28944 0.178
R55786 vdd.n27955 vdd.n27954 0.178
R55787 vdd.n29902 vdd.n29901 0.178
R55788 vdd.n30642 vdd.n30641 0.178
R55789 vdd.n30614 vdd.n30613 0.178
R55790 vdd.n28943 vdd.n28942 0.178
R55791 vdd.n29900 vdd.n29899 0.178
R55792 vdd.n30258 vdd.n30257 0.178
R55793 vdd.n27596 vdd.n27595 0.178
R55794 vdd.n26012 vdd.n26011 0.178
R55795 vdd.n25384 vdd.n25383 0.178
R55796 vdd.n34065 vdd.n34064 0.177
R55797 vdd.n35226 vdd.n35225 0.177
R55798 vdd.n34639 vdd.n34638 0.177
R55799 vdd.n6349 vdd.n6348 0.177
R55800 vdd.n5386 vdd.n5385 0.177
R55801 vdd.n4216 vdd.n4215 0.177
R55802 vdd.n37104 vdd.n37103 0.177
R55803 vdd.n37135 vdd.n37134 0.177
R55804 vdd.n37289 vdd.n37288 0.177
R55805 vdd.n32998 vdd.n32997 0.177
R55806 vdd.n32871 vdd.n32870 0.177
R55807 vdd.n37532 vdd.n37531 0.177
R55808 vdd.n28907 vdd.n28906 0.177
R55809 vdd.n27896 vdd.n27895 0.177
R55810 vdd.n30180 vdd.n30179 0.177
R55811 vdd.n3770 vdd.n3769 0.177
R55812 vdd.n2358 vdd.n2357 0.177
R55813 vdd.n1206 vdd.n1205 0.177
R55814 vdd.n26327 vdd.n26326 0.177
R55815 vdd.n31591 vdd.n31590 0.177
R55816 vdd.n32410 vdd.n32409 0.177
R55817 vdd.n1748 vdd.n1731 0.177
R55818 vdd.n12600 vdd.n10088 0.177
R55819 vdd.n11466 vdd.n11429 0.176
R55820 vdd.n11469 vdd.n11428 0.176
R55821 vdd.n15038 vdd.n15036 0.176
R55822 vdd.n16818 vdd.n16817 0.176
R55823 vdd.n28825 vdd.n28824 0.175
R55824 vdd.n11746 vdd.n11722 0.175
R55825 vdd.n32277 vdd.n31538 0.175
R55826 vdd.n28831 vdd.n28830 0.175
R55827 vdd.n1782 vdd.n1776 0.175
R55828 vdd.n1782 vdd.n1778 0.175
R55829 vdd.n2601 vdd.n2595 0.175
R55830 vdd.n2601 vdd.n2597 0.175
R55831 vdd.n2218 vdd.n2212 0.175
R55832 vdd.n2218 vdd.n2214 0.175
R55833 vdd.n10230 vdd.n10229 0.171
R55834 vdd.n16645 vdd.n16644 0.171
R55835 vdd.n38139 vdd.n38138 0.17
R55836 vdd.n3976 vdd.n3975 0.166
R55837 vdd.n3884 vdd.n3883 0.166
R55838 vdd.n2345 vdd.n2344 0.166
R55839 vdd.n2513 vdd.n2512 0.166
R55840 vdd.n1948 vdd.n1947 0.166
R55841 vdd.n1248 vdd.n1247 0.166
R55842 vdd.n3882 vdd.n3881 0.166
R55843 vdd.n2438 vdd.n2437 0.166
R55844 vdd.n1246 vdd.n1245 0.166
R55845 vdd.n470 vdd.n469 0.166
R55846 vdd.n33205 vdd.n33204 0.166
R55847 vdd.n33154 vdd.n33153 0.166
R55848 vdd.n37267 vdd.n37266 0.166
R55849 vdd.n37332 vdd.n37331 0.166
R55850 vdd.n37485 vdd.n37484 0.166
R55851 vdd.n37540 vdd.n37539 0.166
R55852 vdd.n33210 vdd.n33209 0.166
R55853 vdd.n33156 vdd.n33155 0.166
R55854 vdd.n37269 vdd.n37268 0.166
R55855 vdd.n37334 vdd.n37333 0.166
R55856 vdd.n37487 vdd.n37486 0.166
R55857 vdd.n37542 vdd.n37541 0.166
R55858 vdd.n26290 vdd.n26289 0.166
R55859 vdd.n31818 vdd.n31817 0.166
R55860 vdd.n31602 vdd.n31601 0.166
R55861 vdd.n32176 vdd.n32175 0.166
R55862 vdd.n31445 vdd.n31444 0.166
R55863 vdd.n31062 vdd.n31061 0.166
R55864 vdd.n31816 vdd.n31815 0.166
R55865 vdd.n32174 vdd.n32173 0.166
R55866 vdd.n31060 vdd.n31059 0.166
R55867 vdd.n28896 vdd.n28895 0.166
R55868 vdd.n28957 vdd.n28956 0.166
R55869 vdd.n27963 vdd.n27962 0.166
R55870 vdd.n29915 vdd.n29914 0.166
R55871 vdd.n30651 vdd.n30650 0.166
R55872 vdd.n30605 vdd.n30604 0.166
R55873 vdd.n28955 vdd.n28954 0.166
R55874 vdd.n29913 vdd.n29912 0.166
R55875 vdd.n30262 vdd.n30261 0.166
R55876 vdd.n25388 vdd.n25387 0.166
R55877 vdd.n10248 vdd.n10225 0.166
R55878 vdd.n10232 vdd.n10069 0.166
R55879 vdd.n33456 vdd.n33455 0.166
R55880 vdd.n775 vdd.n774 0.166
R55881 vdd.n28894 vdd.n28893 0.166
R55882 vdd.n27870 vdd.n27869 0.166
R55883 vdd.n30176 vdd.n30175 0.166
R55884 vdd.n25457 vdd.n25456 0.166
R55885 vdd.n3764 vdd.n3763 0.166
R55886 vdd.n2343 vdd.n2342 0.166
R55887 vdd.n1940 vdd.n1939 0.166
R55888 vdd.n26288 vdd.n26287 0.166
R55889 vdd.n31604 vdd.n31603 0.166
R55890 vdd.n31443 vdd.n31442 0.166
R55891 vdd.n32071 vdd.n32070 0.166
R55892 vdd.n11753 vdd.n11752 0.164
R55893 vdd.n21833 vdd.n21832 0.164
R55894 vdd.n12600 vdd.n10067 0.163
R55895 vdd.n11803 vdd.n11802 0.163
R55896 vdd.n21894 vdd.n21893 0.163
R55897 vdd.n24911 vdd.n24892 0.163
R55898 vdd.n31939 vdd.n31670 0.162
R55899 vdd.n31973 vdd.n31643 0.162
R55900 vdd.n32047 vdd.n31587 0.162
R55901 vdd.n32306 vdd.n31519 0.162
R55902 vdd.n31761 vdd.n31739 0.162
R55903 vdd.n27241 vdd.n27214 0.162
R55904 vdd.n26609 vdd.n26604 0.162
R55905 vdd.n26402 vdd.n26396 0.162
R55906 vdd.n26302 vdd.n26300 0.162
R55907 vdd.n25252 vdd.n24976 0.161
R55908 vdd.n25140 vdd.n25054 0.161
R55909 vdd.n24722 vdd.n24635 0.161
R55910 vdd.n4658 vdd.n4657 0.158
R55911 vdd.n2692 vdd.n2691 0.156
R55912 vdd.n3841 vdd.n3838 0.156
R55913 vdd.n9995 vdd.n9972 0.156
R55914 vdd.n12684 vdd.n12683 0.156
R55915 vdd.n12781 vdd.n9780 0.156
R55916 vdd.n9795 vdd.n9785 0.156
R55917 vdd.n9635 vdd.n9612 0.156
R55918 vdd.n12892 vdd.n12891 0.156
R55919 vdd.n12989 vdd.n9419 0.156
R55920 vdd.n9436 vdd.n9425 0.156
R55921 vdd.n10377 vdd.n10376 0.156
R55922 vdd.n10346 vdd.n10341 0.156
R55923 vdd.n15136 vdd.n15134 0.156
R55924 vdd.n15150 vdd.n15148 0.156
R55925 vdd.n15164 vdd.n15162 0.156
R55926 vdd.n15178 vdd.n15176 0.156
R55927 vdd.n15192 vdd.n15180 0.156
R55928 vdd.n15206 vdd.n15204 0.156
R55929 vdd.n15220 vdd.n15218 0.156
R55930 vdd.n15234 vdd.n15232 0.156
R55931 vdd.n15245 vdd.n15243 0.156
R55932 vdd.n15256 vdd.n15254 0.156
R55933 vdd.n34012 vdd.n34011 0.156
R55934 vdd.n35175 vdd.n35174 0.156
R55935 vdd.n34600 vdd.n34599 0.156
R55936 vdd.n6312 vdd.n6311 0.156
R55937 vdd.n5347 vdd.n5346 0.156
R55938 vdd.n4178 vdd.n4177 0.156
R55939 vdd.n4876 vdd.n4875 0.155
R55940 vdd.n3991 vdd.n3990 0.155
R55941 vdd.n3872 vdd.n3871 0.155
R55942 vdd.n2326 vdd.n2325 0.155
R55943 vdd.n2499 vdd.n2498 0.155
R55944 vdd.n2079 vdd.n2078 0.155
R55945 vdd.n1824 vdd.n1823 0.155
R55946 vdd.n3870 vdd.n3869 0.155
R55947 vdd.n2448 vdd.n2447 0.155
R55948 vdd.n1822 vdd.n1821 0.155
R55949 vdd.n37087 vdd.n37086 0.155
R55950 vdd.n37163 vdd.n37162 0.155
R55951 vdd.n33049 vdd.n33048 0.155
R55952 vdd.n37344 vdd.n37343 0.155
R55953 vdd.n32882 vdd.n32881 0.155
R55954 vdd.n32821 vdd.n32820 0.155
R55955 vdd.n26685 vdd.n26684 0.155
R55956 vdd.n31837 vdd.n31836 0.155
R55957 vdd.n31608 vdd.n31607 0.155
R55958 vdd.n32198 vdd.n32197 0.155
R55959 vdd.n32371 vdd.n32370 0.155
R55960 vdd.n31085 vdd.n31084 0.155
R55961 vdd.n31835 vdd.n31834 0.155
R55962 vdd.n32196 vdd.n32195 0.155
R55963 vdd.n31083 vdd.n31082 0.155
R55964 vdd.n28881 vdd.n28880 0.155
R55965 vdd.n29002 vdd.n29001 0.155
R55966 vdd.n27972 vdd.n27971 0.155
R55967 vdd.n29928 vdd.n29927 0.155
R55968 vdd.n30669 vdd.n30668 0.155
R55969 vdd.n30596 vdd.n30595 0.155
R55970 vdd.n29000 vdd.n28999 0.155
R55971 vdd.n29926 vdd.n29925 0.155
R55972 vdd.n30281 vdd.n30280 0.155
R55973 vdd.n37079 vdd.n37078 0.155
R55974 vdd.n37161 vdd.n37160 0.155
R55975 vdd.n33044 vdd.n33043 0.155
R55976 vdd.n37342 vdd.n37341 0.155
R55977 vdd.n32880 vdd.n32879 0.155
R55978 vdd.n32819 vdd.n32818 0.155
R55979 vdd.n28879 vdd.n28878 0.155
R55980 vdd.n27865 vdd.n27864 0.155
R55981 vdd.n30667 vdd.n30666 0.155
R55982 vdd.n3749 vdd.n3748 0.155
R55983 vdd.n2324 vdd.n2323 0.155
R55984 vdd.n2074 vdd.n2073 0.155
R55985 vdd.n26675 vdd.n26674 0.155
R55986 vdd.n31606 vdd.n31605 0.155
R55987 vdd.n32373 vdd.n32372 0.155
R55988 vdd.n24942 vdd.n24941 0.155
R55989 vdd.n32408 vdd.n32406 0.154
R55990 vdd.n1771 vdd.n1770 0.154
R55991 vdd.n13086 vdd.n13085 0.153
R55992 vdd.n19299 vdd.n14976 0.153
R55993 vdd.n11727 vdd.n11720 0.151
R55994 vdd.n21800 vdd.n21799 0.151
R55995 vdd.n31286 vdd.n31281 0.15
R55996 vdd.n31936 vdd.n31675 0.15
R55997 vdd.n31936 vdd.n31924 0.15
R55998 vdd.n31537 vdd.n31532 0.15
R55999 vdd.n32296 vdd.n31529 0.15
R56000 vdd.n32306 vdd.n32305 0.15
R56001 vdd.n31761 vdd.n31740 0.15
R56002 vdd.n27238 vdd.n27230 0.15
R56003 vdd.n26155 vdd.n26154 0.15
R56004 vdd.n26609 vdd.n26605 0.15
R56005 vdd.n31071 vdd.n31069 0.149
R56006 vdd.n32185 vdd.n32183 0.149
R56007 vdd.n31824 vdd.n31716 0.149
R56008 vdd.n24974 vdd.n24883 0.149
R56009 vdd.n11845 vdd.n11844 0.146
R56010 vdd.n21936 vdd.n21935 0.146
R56011 ldomc_0.pmosm_0.vdd vdd.n38216 0.145
R56012 vdd.n35214 vdd.n35213 0.144
R56013 vdd.n6338 vdd.n6337 0.144
R56014 vdd.n11918 vdd.n11662 0.144
R56015 vdd.n4006 vdd.n4005 0.144
R56016 vdd.n3857 vdd.n3856 0.144
R56017 vdd.n2307 vdd.n2306 0.144
R56018 vdd.n2482 vdd.n2481 0.144
R56019 vdd.n2088 vdd.n2087 0.144
R56020 vdd.n1801 vdd.n1800 0.144
R56021 vdd.n3831 vdd.n3830 0.144
R56022 vdd.n2456 vdd.n2455 0.144
R56023 vdd.n1259 vdd.n1258 0.144
R56024 vdd.n36983 vdd.n36982 0.144
R56025 vdd.n33231 vdd.n33230 0.144
R56026 vdd.n35624 vdd.n35623 0.144
R56027 vdd.n37244 vdd.n37243 0.144
R56028 vdd.n32965 vdd.n32964 0.144
R56029 vdd.n32899 vdd.n32898 0.144
R56030 vdd.n37559 vdd.n37558 0.144
R56031 vdd.n36985 vdd.n36984 0.144
R56032 vdd.n33239 vdd.n33238 0.144
R56033 vdd.n35626 vdd.n35625 0.144
R56034 vdd.n37249 vdd.n37248 0.144
R56035 vdd.n32967 vdd.n32966 0.144
R56036 vdd.n32904 vdd.n32903 0.144
R56037 vdd.n37561 vdd.n37560 0.144
R56038 vdd.n26611 vdd.n26610 0.144
R56039 vdd.n31862 vdd.n31861 0.144
R56040 vdd.n32000 vdd.n31999 0.144
R56041 vdd.n32220 vdd.n32219 0.144
R56042 vdd.n31467 vdd.n31466 0.144
R56043 vdd.n31114 vdd.n31113 0.144
R56044 vdd.n31860 vdd.n31859 0.144
R56045 vdd.n32218 vdd.n32217 0.144
R56046 vdd.n31112 vdd.n31111 0.144
R56047 vdd.n28869 vdd.n28868 0.144
R56048 vdd.n29015 vdd.n29014 0.144
R56049 vdd.n27994 vdd.n27993 0.144
R56050 vdd.n29936 vdd.n29935 0.144
R56051 vdd.n30657 vdd.n30656 0.144
R56052 vdd.n30586 vdd.n30585 0.144
R56053 vdd.n29013 vdd.n29012 0.144
R56054 vdd.n29933 vdd.n29932 0.144
R56055 vdd.n30290 vdd.n30289 0.144
R56056 vdd.n25000 vdd.n24999 0.144
R56057 vdd.n24576 vdd.n24575 0.144
R56058 vdd.n2761 vdd.n2754 0.144
R56059 vdd.n2772 vdd.n2765 0.144
R56060 vdd.n2783 vdd.n2776 0.144
R56061 vdd.n2794 vdd.n2787 0.144
R56062 vdd.n2813 vdd.n2811 0.144
R56063 vdd.n2824 vdd.n2822 0.144
R56064 vdd.n2835 vdd.n2833 0.144
R56065 vdd.n2846 vdd.n2844 0.144
R56066 vdd.n2857 vdd.n2855 0.144
R56067 vdd.n2868 vdd.n2866 0.144
R56068 vdd.n2879 vdd.n2877 0.144
R56069 vdd.n2909 vdd.n2902 0.144
R56070 vdd.n2920 vdd.n2913 0.144
R56071 vdd.n2931 vdd.n2924 0.144
R56072 vdd.n2942 vdd.n2935 0.144
R56073 vdd.n2953 vdd.n2946 0.144
R56074 vdd.n2964 vdd.n2957 0.144
R56075 vdd.n2975 vdd.n2968 0.144
R56076 vdd.n2994 vdd.n2992 0.144
R56077 vdd.n3005 vdd.n3003 0.144
R56078 vdd.n3016 vdd.n3014 0.144
R56079 vdd.n3027 vdd.n3025 0.144
R56080 vdd.n3038 vdd.n3036 0.144
R56081 vdd.n3049 vdd.n3047 0.144
R56082 vdd.n3060 vdd.n3058 0.144
R56083 vdd.n3090 vdd.n3083 0.144
R56084 vdd.n3101 vdd.n3094 0.144
R56085 vdd.n3112 vdd.n3105 0.144
R56086 vdd.n3123 vdd.n3116 0.144
R56087 vdd.n3134 vdd.n3127 0.144
R56088 vdd.n3145 vdd.n3138 0.144
R56089 vdd.n3156 vdd.n3149 0.144
R56090 vdd.n3175 vdd.n3173 0.144
R56091 vdd.n3186 vdd.n3184 0.144
R56092 vdd.n3197 vdd.n3195 0.144
R56093 vdd.n3208 vdd.n3206 0.144
R56094 vdd.n3219 vdd.n3217 0.144
R56095 vdd.n3230 vdd.n3228 0.144
R56096 vdd.n3241 vdd.n3239 0.144
R56097 vdd.n3271 vdd.n3264 0.144
R56098 vdd.n3282 vdd.n3275 0.144
R56099 vdd.n3293 vdd.n3286 0.144
R56100 vdd.n3304 vdd.n3297 0.144
R56101 vdd.n3315 vdd.n3308 0.144
R56102 vdd.n3326 vdd.n3319 0.144
R56103 vdd.n3337 vdd.n3330 0.144
R56104 vdd.n3356 vdd.n3354 0.144
R56105 vdd.n3367 vdd.n3365 0.144
R56106 vdd.n3378 vdd.n3376 0.144
R56107 vdd.n3389 vdd.n3387 0.144
R56108 vdd.n3400 vdd.n3398 0.144
R56109 vdd.n3411 vdd.n3409 0.144
R56110 vdd.n3422 vdd.n3420 0.144
R56111 vdd.n3452 vdd.n3445 0.144
R56112 vdd.n3463 vdd.n3456 0.144
R56113 vdd.n3474 vdd.n3467 0.144
R56114 vdd.n3485 vdd.n3478 0.144
R56115 vdd.n3496 vdd.n3489 0.144
R56116 vdd.n3507 vdd.n3500 0.144
R56117 vdd.n3518 vdd.n3511 0.144
R56118 vdd.n3537 vdd.n3535 0.144
R56119 vdd.n3548 vdd.n3546 0.144
R56120 vdd.n3559 vdd.n3557 0.144
R56121 vdd.n3570 vdd.n3568 0.144
R56122 vdd.n3581 vdd.n3579 0.144
R56123 vdd.n3592 vdd.n3590 0.144
R56124 vdd.n3603 vdd.n3601 0.144
R56125 vdd.n1761 vdd.n1759 0.144
R56126 vdd.n35872 vdd.n35862 0.144
R56127 vdd.n35886 vdd.n35876 0.144
R56128 vdd.n35900 vdd.n35890 0.144
R56129 vdd.n35914 vdd.n35904 0.144
R56130 vdd.n35937 vdd.n35935 0.144
R56131 vdd.n35951 vdd.n35949 0.144
R56132 vdd.n35965 vdd.n35963 0.144
R56133 vdd.n35979 vdd.n35977 0.144
R56134 vdd.n35993 vdd.n35991 0.144
R56135 vdd.n36007 vdd.n36005 0.144
R56136 vdd.n36021 vdd.n36019 0.144
R56137 vdd.n36061 vdd.n36051 0.144
R56138 vdd.n36075 vdd.n36065 0.144
R56139 vdd.n36089 vdd.n36079 0.144
R56140 vdd.n36103 vdd.n36093 0.144
R56141 vdd.n36117 vdd.n36107 0.144
R56142 vdd.n36131 vdd.n36121 0.144
R56143 vdd.n36145 vdd.n36135 0.144
R56144 vdd.n36168 vdd.n36166 0.144
R56145 vdd.n36182 vdd.n36180 0.144
R56146 vdd.n36196 vdd.n36194 0.144
R56147 vdd.n36210 vdd.n36208 0.144
R56148 vdd.n36224 vdd.n36222 0.144
R56149 vdd.n36238 vdd.n36236 0.144
R56150 vdd.n36252 vdd.n36250 0.144
R56151 vdd.n36292 vdd.n36282 0.144
R56152 vdd.n36306 vdd.n36296 0.144
R56153 vdd.n36320 vdd.n36310 0.144
R56154 vdd.n36334 vdd.n36324 0.144
R56155 vdd.n36348 vdd.n36338 0.144
R56156 vdd.n36362 vdd.n36352 0.144
R56157 vdd.n36376 vdd.n36366 0.144
R56158 vdd.n36399 vdd.n36397 0.144
R56159 vdd.n36413 vdd.n36411 0.144
R56160 vdd.n36427 vdd.n36425 0.144
R56161 vdd.n36441 vdd.n36439 0.144
R56162 vdd.n36455 vdd.n36453 0.144
R56163 vdd.n36469 vdd.n36467 0.144
R56164 vdd.n36483 vdd.n36481 0.144
R56165 vdd.n36523 vdd.n36513 0.144
R56166 vdd.n36537 vdd.n36527 0.144
R56167 vdd.n36551 vdd.n36541 0.144
R56168 vdd.n36565 vdd.n36555 0.144
R56169 vdd.n36579 vdd.n36569 0.144
R56170 vdd.n36593 vdd.n36583 0.144
R56171 vdd.n36607 vdd.n36597 0.144
R56172 vdd.n36630 vdd.n36628 0.144
R56173 vdd.n36644 vdd.n36642 0.144
R56174 vdd.n36658 vdd.n36656 0.144
R56175 vdd.n36672 vdd.n36670 0.144
R56176 vdd.n36686 vdd.n36684 0.144
R56177 vdd.n36700 vdd.n36698 0.144
R56178 vdd.n36714 vdd.n36712 0.144
R56179 vdd.n36754 vdd.n36744 0.144
R56180 vdd.n36768 vdd.n36758 0.144
R56181 vdd.n36782 vdd.n36772 0.144
R56182 vdd.n36796 vdd.n36786 0.144
R56183 vdd.n36810 vdd.n36800 0.144
R56184 vdd.n36824 vdd.n36814 0.144
R56185 vdd.n36838 vdd.n36828 0.144
R56186 vdd.n36861 vdd.n36859 0.144
R56187 vdd.n36875 vdd.n36873 0.144
R56188 vdd.n36889 vdd.n36887 0.144
R56189 vdd.n36903 vdd.n36901 0.144
R56190 vdd.n36917 vdd.n36915 0.144
R56191 vdd.n36931 vdd.n36929 0.144
R56192 vdd.n36945 vdd.n36943 0.144
R56193 vdd.n38110 vdd.n38100 0.144
R56194 vdd.n38096 vdd.n38086 0.144
R56195 vdd.n38082 vdd.n38072 0.144
R56196 vdd.n38068 vdd.n38058 0.144
R56197 vdd.n38054 vdd.n38044 0.144
R56198 vdd.n38040 vdd.n38030 0.144
R56199 vdd.n38000 vdd.n37998 0.144
R56200 vdd.n37986 vdd.n37984 0.144
R56201 vdd.n37972 vdd.n37970 0.144
R56202 vdd.n37958 vdd.n37956 0.144
R56203 vdd.n37944 vdd.n37942 0.144
R56204 vdd.n37930 vdd.n37928 0.144
R56205 vdd.n37916 vdd.n37914 0.144
R56206 vdd.n37893 vdd.n37883 0.144
R56207 vdd.n37879 vdd.n37869 0.144
R56208 vdd.n37865 vdd.n37855 0.144
R56209 vdd.n37851 vdd.n37841 0.144
R56210 vdd.n37837 vdd.n37827 0.144
R56211 vdd.n37823 vdd.n37813 0.144
R56212 vdd.n37809 vdd.n37799 0.144
R56213 vdd.n37769 vdd.n37767 0.144
R56214 vdd.n37755 vdd.n37753 0.144
R56215 vdd.n37741 vdd.n37739 0.144
R56216 vdd.n37727 vdd.n37725 0.144
R56217 vdd.n37713 vdd.n37711 0.144
R56218 vdd.n37699 vdd.n37697 0.144
R56219 vdd.n37685 vdd.n37683 0.144
R56220 vdd.n37662 vdd.n37652 0.144
R56221 vdd.n37648 vdd.n37638 0.144
R56222 vdd.n37634 vdd.n37624 0.144
R56223 vdd.n37620 vdd.n37610 0.144
R56224 vdd.n28197 vdd.n28195 0.144
R56225 vdd.n28211 vdd.n28209 0.144
R56226 vdd.n28251 vdd.n28241 0.144
R56227 vdd.n28265 vdd.n28255 0.144
R56228 vdd.n28279 vdd.n28269 0.144
R56229 vdd.n28293 vdd.n28283 0.144
R56230 vdd.n28307 vdd.n28297 0.144
R56231 vdd.n28321 vdd.n28311 0.144
R56232 vdd.n28335 vdd.n28325 0.144
R56233 vdd.n28358 vdd.n28356 0.144
R56234 vdd.n28372 vdd.n28370 0.144
R56235 vdd.n28386 vdd.n28384 0.144
R56236 vdd.n28400 vdd.n28398 0.144
R56237 vdd.n28414 vdd.n28412 0.144
R56238 vdd.n28428 vdd.n28426 0.144
R56239 vdd.n28442 vdd.n28440 0.144
R56240 vdd.n28482 vdd.n28472 0.144
R56241 vdd.n28496 vdd.n28486 0.144
R56242 vdd.n28510 vdd.n28500 0.144
R56243 vdd.n28524 vdd.n28514 0.144
R56244 vdd.n28538 vdd.n28528 0.144
R56245 vdd.n28552 vdd.n28542 0.144
R56246 vdd.n28566 vdd.n28556 0.144
R56247 vdd.n28589 vdd.n28587 0.144
R56248 vdd.n28603 vdd.n28601 0.144
R56249 vdd.n28617 vdd.n28615 0.144
R56250 vdd.n28631 vdd.n28629 0.144
R56251 vdd.n28645 vdd.n28643 0.144
R56252 vdd.n28659 vdd.n28657 0.144
R56253 vdd.n28673 vdd.n28671 0.144
R56254 vdd.n28713 vdd.n28703 0.144
R56255 vdd.n28727 vdd.n28717 0.144
R56256 vdd.n28741 vdd.n28731 0.144
R56257 vdd.n28755 vdd.n28745 0.144
R56258 vdd.n28769 vdd.n28759 0.144
R56259 vdd.n28783 vdd.n28773 0.144
R56260 vdd.n28797 vdd.n28787 0.144
R56261 vdd.n1726 vdd.n1719 0.144
R56262 vdd.n1715 vdd.n1708 0.144
R56263 vdd.n1704 vdd.n1697 0.144
R56264 vdd.n1693 vdd.n1686 0.144
R56265 vdd.n1682 vdd.n1675 0.144
R56266 vdd.n1671 vdd.n1664 0.144
R56267 vdd.n1641 vdd.n1639 0.144
R56268 vdd.n1630 vdd.n1628 0.144
R56269 vdd.n1619 vdd.n1617 0.144
R56270 vdd.n1608 vdd.n1606 0.144
R56271 vdd.n1597 vdd.n1595 0.144
R56272 vdd.n1586 vdd.n1584 0.144
R56273 vdd.n1575 vdd.n1573 0.144
R56274 vdd.n1556 vdd.n1549 0.144
R56275 vdd.n1545 vdd.n1538 0.144
R56276 vdd.n1534 vdd.n1527 0.144
R56277 vdd.n1523 vdd.n1516 0.144
R56278 vdd.n1512 vdd.n1505 0.144
R56279 vdd.n1501 vdd.n1494 0.144
R56280 vdd.n1490 vdd.n1483 0.144
R56281 vdd.n1460 vdd.n1458 0.144
R56282 vdd.n1449 vdd.n1447 0.144
R56283 vdd.n1438 vdd.n1436 0.144
R56284 vdd.n1427 vdd.n1425 0.144
R56285 vdd.n1416 vdd.n1414 0.144
R56286 vdd.n1405 vdd.n1403 0.144
R56287 vdd.n1394 vdd.n1392 0.144
R56288 vdd.n1375 vdd.n1368 0.144
R56289 vdd.n1364 vdd.n1357 0.144
R56290 vdd.n1353 vdd.n1346 0.144
R56291 vdd.n1342 vdd.n1335 0.144
R56292 vdd.n1331 vdd.n1324 0.144
R56293 vdd.n1320 vdd.n1313 0.144
R56294 vdd.n1309 vdd.n1302 0.144
R56295 vdd.n26775 vdd.n26768 0.144
R56296 vdd.n26786 vdd.n26779 0.144
R56297 vdd.n26797 vdd.n26790 0.144
R56298 vdd.n26808 vdd.n26801 0.144
R56299 vdd.n26819 vdd.n26812 0.144
R56300 vdd.n26830 vdd.n26823 0.144
R56301 vdd.n26841 vdd.n26834 0.144
R56302 vdd.n26860 vdd.n26858 0.144
R56303 vdd.n26871 vdd.n26869 0.144
R56304 vdd.n26882 vdd.n26880 0.144
R56305 vdd.n26893 vdd.n26891 0.144
R56306 vdd.n26904 vdd.n26902 0.144
R56307 vdd.n26915 vdd.n26913 0.144
R56308 vdd.n26926 vdd.n26924 0.144
R56309 vdd.n26956 vdd.n26949 0.144
R56310 vdd.n26967 vdd.n26960 0.144
R56311 vdd.n26978 vdd.n26971 0.144
R56312 vdd.n26989 vdd.n26982 0.144
R56313 vdd.n27000 vdd.n26993 0.144
R56314 vdd.n27011 vdd.n27004 0.144
R56315 vdd.n27022 vdd.n27015 0.144
R56316 vdd.n27041 vdd.n27039 0.144
R56317 vdd.n27052 vdd.n27050 0.144
R56318 vdd.n27063 vdd.n27061 0.144
R56319 vdd.n27074 vdd.n27072 0.144
R56320 vdd.n27085 vdd.n27083 0.144
R56321 vdd.n27096 vdd.n27094 0.144
R56322 vdd.n27107 vdd.n27105 0.144
R56323 vdd.n27137 vdd.n27130 0.144
R56324 vdd.n27148 vdd.n27141 0.144
R56325 vdd.n27159 vdd.n27152 0.144
R56326 vdd.n27170 vdd.n27163 0.144
R56327 vdd.n27181 vdd.n27174 0.144
R56328 vdd.n27192 vdd.n27185 0.144
R56329 vdd.n27203 vdd.n27196 0.144
R56330 vdd.n11702 vdd.n11701 0.144
R56331 vdd.n21774 vdd.n21772 0.144
R56332 vdd.n25042 vdd.n25039 0.144
R56333 vdd.n25035 vdd.n25032 0.144
R56334 vdd.n25017 vdd.n25015 0.144
R56335 vdd.n25010 vdd.n25008 0.144
R56336 vdd.n25003 vdd.n25001 0.144
R56337 vdd.n24617 vdd.n24614 0.144
R56338 vdd.n24610 vdd.n24607 0.144
R56339 vdd.n24593 vdd.n24591 0.144
R56340 vdd.n24586 vdd.n24584 0.144
R56341 vdd.n24579 vdd.n24577 0.144
R56342 vdd.n34053 vdd.n34052 0.144
R56343 vdd.n34627 vdd.n34626 0.144
R56344 vdd.n5374 vdd.n5373 0.144
R56345 vdd.n5168 vdd.n5167 0.144
R56346 vdd.n4204 vdd.n4203 0.144
R56347 vdd.n27605 vdd.n27604 0.144
R56348 vdd.n26021 vdd.n26020 0.144
R56349 vdd.n28867 vdd.n28866 0.144
R56350 vdd.n27860 vdd.n27859 0.144
R56351 vdd.n30655 vdd.n30654 0.144
R56352 vdd.n3732 vdd.n3731 0.144
R56353 vdd.n2305 vdd.n2304 0.144
R56354 vdd.n2086 vdd.n2085 0.144
R56355 vdd.n26603 vdd.n26602 0.144
R56356 vdd.n31998 vdd.n31997 0.144
R56357 vdd.n31465 vdd.n31464 0.144
R56358 vdd.n10249 vdd.n10130 0.141
R56359 vdd.n31451 vdd.n31450 0.137
R56360 vdd.n31562 vdd.n31561 0.137
R56361 vdd.n31554 vdd.n31553 0.137
R56362 vdd.n31745 vdd.n31741 0.137
R56363 vdd.n27241 vdd.n27209 0.137
R56364 vdd.n26595 vdd.n26592 0.137
R56365 vdd.n31707 vdd.n31705 0.137
R56366 vdd.n31161 vdd.n31160 0.135
R56367 vdd.n24567 vdd.n24533 0.134
R56368 vdd.n11784 vdd.n11777 0.134
R56369 vdd.n21876 vdd.n21869 0.134
R56370 vdd.n35384 vdd.n35383 0.133
R56371 vdd.n6077 vdd.n6076 0.133
R56372 vdd.n3716 vdd.n3715 0.133
R56373 vdd.n3836 vdd.n3835 0.133
R56374 vdd.n2289 vdd.n2288 0.133
R56375 vdd.n2462 vdd.n2461 0.133
R56376 vdd.n1997 vdd.n1996 0.133
R56377 vdd.n3834 vdd.n3833 0.133
R56378 vdd.n2460 vdd.n2459 0.133
R56379 vdd.n36999 vdd.n36998 0.133
R56380 vdd.n37074 vdd.n37073 0.133
R56381 vdd.n33120 vdd.n33119 0.133
R56382 vdd.n33086 vdd.n33085 0.133
R56383 vdd.n37374 vdd.n37373 0.133
R56384 vdd.n37455 vdd.n37454 0.133
R56385 vdd.n37586 vdd.n37585 0.133
R56386 vdd.n26590 vdd.n26589 0.133
R56387 vdd.n31879 vdd.n31878 0.133
R56388 vdd.n31985 vdd.n31984 0.133
R56389 vdd.n32252 vdd.n32251 0.133
R56390 vdd.n32344 vdd.n32343 0.133
R56391 vdd.n31183 vdd.n31182 0.133
R56392 vdd.n31877 vdd.n31876 0.133
R56393 vdd.n32250 vdd.n32249 0.133
R56394 vdd.n31127 vdd.n31126 0.133
R56395 vdd.n28857 vdd.n28856 0.133
R56396 vdd.n28043 vdd.n28042 0.133
R56397 vdd.n28003 vdd.n28002 0.133
R56398 vdd.n29797 vdd.n29796 0.133
R56399 vdd.n29731 vdd.n29730 0.133
R56400 vdd.n30307 vdd.n30306 0.133
R56401 vdd.n27773 vdd.n27772 0.133
R56402 vdd.n29795 vdd.n29794 0.133
R56403 vdd.n30309 vdd.n30308 0.133
R56404 vdd.n24616 vdd.n24615 0.133
R56405 vdd.n24583 vdd.n24582 0.133
R56406 vdd.n34426 vdd.n34425 0.132
R56407 vdd.n34856 vdd.n34855 0.132
R56408 vdd.n5603 vdd.n5602 0.132
R56409 vdd.n4718 vdd.n4717 0.132
R56410 vdd.n4430 vdd.n4429 0.132
R56411 vdd.n27647 vdd.n27646 0.132
R56412 vdd.n26069 vdd.n26068 0.132
R56413 vdd.n36997 vdd.n36996 0.132
R56414 vdd.n37066 vdd.n37065 0.132
R56415 vdd.n33118 vdd.n33117 0.132
R56416 vdd.n33078 vdd.n33077 0.132
R56417 vdd.n37372 vdd.n37371 0.132
R56418 vdd.n37450 vdd.n37449 0.132
R56419 vdd.n37584 vdd.n37583 0.132
R56420 vdd.n28855 vdd.n28854 0.132
R56421 vdd.n27855 vdd.n27854 0.132
R56422 vdd.n29707 vdd.n29706 0.132
R56423 vdd.n25528 vdd.n25527 0.132
R56424 vdd.n3714 vdd.n3713 0.132
R56425 vdd.n2287 vdd.n2286 0.132
R56426 vdd.n1982 vdd.n1981 0.132
R56427 vdd.n26588 vdd.n26587 0.132
R56428 vdd.n31983 vdd.n31982 0.132
R56429 vdd.n32342 vdd.n32341 0.132
R56430 vdd.n25007 vdd.n25006 0.132
R56431 vdd.n25041 vdd.n25040 0.132
R56432 vdd.n12600 vdd.n10078 0.132
R56433 vdd.n38155 vdd.n38153 0.127
R56434 vdd.n27482 vdd.n27480 0.127
R56435 vdd.n25918 vdd.n25718 0.127
R56436 vdd.n24994 vdd.n24992 0.126
R56437 vdd.n24570 vdd.n24568 0.126
R56438 vdd.n31950 vdd.n31669 0.125
R56439 vdd.n31950 vdd.n31948 0.125
R56440 vdd.n31988 vdd.n31987 0.125
R56441 vdd.n32277 vdd.n32274 0.125
R56442 vdd.n32315 vdd.n32314 0.125
R56443 vdd.n3711 vdd.n2692 0.125
R56444 vdd.n4012 vdd.n3730 0.125
R56445 vdd.n3959 vdd.n3774 0.125
R56446 vdd.n3914 vdd.n3910 0.125
R56447 vdd.n3859 vdd.n3825 0.125
R56448 vdd.n2284 vdd.n2142 0.125
R56449 vdd.n2303 vdd.n2128 0.125
R56450 vdd.n26683 vdd.n26676 0.125
R56451 vdd.n12600 vdd.n10093 0.125
R56452 vdd.n11802 vdd.n11798 0.125
R56453 vdd.n21893 vdd.n21889 0.125
R56454 vdd.n32454 vdd.n32452 0.124
R56455 vdd.n32162 vdd.n32161 0.124
R56456 vdd.n2265 vdd.n2162 0.124
R56457 vdd.n2549 vdd.n2424 0.124
R56458 vdd.n34330 vdd.n34329 0.122
R56459 vdd.n35008 vdd.n35007 0.122
R56460 vdd.n5755 vdd.n5754 0.122
R56461 vdd.n4695 vdd.n4694 0.122
R56462 vdd.n4585 vdd.n4584 0.122
R56463 vdd.n27649 vdd.n27648 0.122
R56464 vdd.n26071 vdd.n26070 0.122
R56465 vdd.n3699 vdd.n3698 0.121
R56466 vdd.n2232 vdd.n2231 0.121
R56467 vdd.n2272 vdd.n2271 0.121
R56468 vdd.n2615 vdd.n2614 0.121
R56469 vdd.n1966 vdd.n1965 0.121
R56470 vdd.n2230 vdd.n2229 0.121
R56471 vdd.n2613 vdd.n2612 0.121
R56472 vdd.n26189 vdd.n26188 0.121
R56473 vdd.n31904 vdd.n31903 0.121
R56474 vdd.n31971 vdd.n31970 0.121
R56475 vdd.n32269 vdd.n32268 0.121
R56476 vdd.n32327 vdd.n32326 0.121
R56477 vdd.n31902 vdd.n31901 0.121
R56478 vdd.n32267 vdd.n32266 0.121
R56479 vdd.n27777 vdd.n27776 0.121
R56480 vdd.n29807 vdd.n29806 0.121
R56481 vdd.n25595 vdd.n25594 0.121
R56482 vdd.n25401 vdd.n25400 0.121
R56483 vdd.n28842 vdd.n28841 0.121
R56484 vdd.n28034 vdd.n28033 0.121
R56485 vdd.n28012 vdd.n28011 0.121
R56486 vdd.n29809 vdd.n29808 0.121
R56487 vdd.n29740 vdd.n29739 0.121
R56488 vdd.n25034 vdd.n25033 0.121
R56489 vdd.n25014 vdd.n25013 0.121
R56490 vdd.n24609 vdd.n24608 0.121
R56491 vdd.n24590 vdd.n24589 0.121
R56492 vdd.n35596 vdd.n35595 0.121
R56493 vdd.n6031 vdd.n6030 0.121
R56494 vdd.n24859 vdd.n24853 0.121
R56495 vdd.n28840 vdd.n28839 0.121
R56496 vdd.n27828 vdd.n27827 0.121
R56497 vdd.n29703 vdd.n29702 0.121
R56498 vdd.n25521 vdd.n25520 0.121
R56499 vdd.n25611 vdd.n25610 0.121
R56500 vdd.n3697 vdd.n3696 0.121
R56501 vdd.n2270 vdd.n2269 0.121
R56502 vdd.n1964 vdd.n1963 0.121
R56503 vdd.n26187 vdd.n26186 0.121
R56504 vdd.n31969 vdd.n31968 0.121
R56505 vdd.n32325 vdd.n32324 0.121
R56506 vdd.n29853 vdd.n29852 0.12
R56507 vdd.n29021 vdd.n29020 0.12
R56508 vdd.n24565 vdd.n24564 0.119
R56509 vdd.n24624 vdd.n24622 0.119
R56510 vdd.n24902 vdd.n24901 0.118
R56511 vdd.n24930 vdd.n24920 0.118
R56512 vdd.n11545 vdd.n11449 0.118
R56513 vdd.n15026 vdd.n15025 0.118
R56514 vdd.n24933 vdd.n24932 0.117
R56515 vdd.n1798 vdd.n1792 0.117
R56516 vdd.n1798 vdd.n1794 0.117
R56517 vdd.n2479 vdd.n2473 0.117
R56518 vdd.n2479 vdd.n2475 0.117
R56519 vdd.n31150 vdd.n31149 0.116
R56520 vdd.n12577 vdd.n12576 0.115
R56521 vdd.n11897 vdd.n11896 0.115
R56522 vdd.n21988 vdd.n21987 0.115
R56523 vdd.n31104 vdd.n31035 0.112
R56524 vdd.n31594 vdd.n31593 0.112
R56525 vdd.n31562 vdd.n31555 0.112
R56526 vdd.n26193 vdd.n26185 0.112
R56527 vdd.n26341 vdd.n26340 0.112
R56528 vdd.n33949 vdd.n33948 0.11
R56529 vdd.n34451 vdd.n34450 0.11
R56530 vdd.n5198 vdd.n5197 0.11
R56531 vdd.n5039 vdd.n5038 0.11
R56532 vdd.n4028 vdd.n4027 0.11
R56533 vdd.n31174 vdd.n31172 0.11
R56534 vdd.n31166 vdd.n31165 0.11
R56535 vdd.n24602 vdd.n24601 0.11
R56536 vdd.n35035 vdd.n35034 0.11
R56537 vdd.n6233 vdd.n6232 0.11
R56538 vdd.n25021 vdd.n25020 0.109
R56539 vdd.n25052 vdd.n24988 0.109
R56540 vdd.n24938 vdd.n24937 0.109
R56541 vdd.n22481 bandgapmd_0.pnp_groupm_0.vdd 0.108
R56542 vdd.n24203 vdd.n24202 0.107
R56543 vdd.n31304 vdd.n31015 0.105
R56544 vdd.n31097 vdd.n31043 0.104
R56545 vdd.n32204 vdd.n31562 0.104
R56546 vdd.n32284 vdd.n31537 0.104
R56547 vdd.n31849 vdd.n31707 0.104
R56548 vdd.n24092 vdd.n24090 0.104
R56549 vdd.n24090 vdd.n24082 0.104
R56550 vdd.n23980 vdd.n23970 0.104
R56551 vdd.n23860 vdd.n23858 0.104
R56552 vdd.n23858 vdd.n23850 0.104
R56553 vdd.n23748 vdd.n23738 0.104
R56554 vdd.n23170 vdd.n23162 0.104
R56555 vdd.n23172 vdd.n23170 0.104
R56556 vdd.n23292 vdd.n23282 0.104
R56557 vdd.n23402 vdd.n23394 0.104
R56558 vdd.n23404 vdd.n23402 0.104
R56559 vdd.n23524 vdd.n23514 0.104
R56560 vdd.n22591 vdd.n22583 0.104
R56561 vdd.n22593 vdd.n22591 0.104
R56562 vdd.n22713 vdd.n22703 0.104
R56563 vdd.n22823 vdd.n22815 0.104
R56564 vdd.n22825 vdd.n22823 0.104
R56565 vdd.n22945 vdd.n22935 0.104
R56566 vdd.n24537 vdd.n24536 0.103
R56567 vdd.n586 vdd.n585 0.102
R56568 vdd.n34072 vdd.n33965 0.102
R56569 vdd.n35234 vdd.n35126 0.102
R56570 vdd.n34647 vdd.n34539 0.102
R56571 vdd.n6357 vdd.n6250 0.102
R56572 vdd.n5394 vdd.n5286 0.102
R56573 vdd.n4224 vdd.n4116 0.102
R56574 vdd.n12582 vdd.n10125 0.101
R56575 vdd.n24864 vdd.n24861 0.101
R56576 vdd.n33474 vdd.n33473 0.101
R56577 vdd.n787 vdd.n786 0.101
R56578 vdd.n31022 vdd.n31018 0.1
R56579 vdd.n32004 vdd.n32003 0.1
R56580 vdd.n32047 vdd.n32046 0.1
R56581 vdd.n32133 vdd.n32132 0.1
R56582 vdd.n31543 vdd.n31539 0.1
R56583 vdd.n32296 vdd.n32293 0.1
R56584 vdd.n32331 vdd.n32330 0.1
R56585 vdd.n26402 vdd.n26392 0.1
R56586 vdd.n32162 vdd.n31576 0.099
R56587 vdd.n25257 bandgapmd_0.vdd 0.099
R56588 vdd.n24875 vdd.n24872 0.099
R56589 vdd.n32129 vdd.n32128 0.099
R56590 vdd.n27486 vdd.n27485 0.098
R56591 vdd.n4800 vdd.n4799 0.098
R56592 vdd.n27376 vdd.n27374 0.098
R56593 vdd.n25819 vdd.n25742 0.098
R56594 vdd.n25707 vdd.n25706 0.098
R56595 vdd.n31500 vdd.n31494 0.098
R56596 vdd.n31500 vdd.n31496 0.098
R56597 vdd.n31660 vdd.n31649 0.098
R56598 vdd.n31660 vdd.n31650 0.098
R56599 vdd.n32432 vdd.n32427 0.098
R56600 vdd.n32432 vdd.n32428 0.098
R56601 vdd.n26177 vdd.n26172 0.098
R56602 vdd.n26177 vdd.n26173 0.098
R56603 vdd.n25996 vdd.n25694 0.098
R56604 vdd.n12582 vdd.n10126 0.095
R56605 vdd.n11903 vdd.n11791 0.095
R56606 vdd.n11763 vdd.n11762 0.095
R56607 vdd.n11752 vdd.n11719 0.095
R56608 vdd.n11878 vdd.n11877 0.095
R56609 vdd.n21994 vdd.n21882 0.095
R56610 vdd.n21843 vdd.n21842 0.095
R56611 vdd.n21832 vdd.n21831 0.095
R56612 vdd.n21969 vdd.n21968 0.095
R56613 vdd.n24853 vdd.n24838 0.095
R56614 vdd.n27486 vdd.n27482 0.094
R56615 vdd.n24513 vdd.n24512 0.094
R56616 vdd.n24911 vdd.n24910 0.093
R56617 vdd.n24572 vdd.n24570 0.092
R56618 vdd.n27569 vdd.n27558 0.091
R56619 vdd.n943 vdd.n940 0.091
R56620 vdd.n11766 vdd.n11676 0.091
R56621 vdd.n11774 vdd.n11664 0.091
R56622 vdd.n11873 vdd.n11872 0.091
R56623 vdd.n21862 vdd.n21861 0.091
R56624 vdd.n21964 vdd.n21963 0.091
R56625 vdd.n25480 vdd.n25478 0.09
R56626 vdd.n11770 vdd.n11769 0.09
R56627 vdd.n21858 vdd.n21857 0.09
R56628 vdd.n25914 vdd.n25913 0.089
R56629 vdd.n25812 vdd.n25811 0.089
R56630 vdd.n26007 vdd.n25999 0.089
R56631 vdd.n10126 vdd.n10124 0.089
R56632 vdd.n11672 vdd.n11668 0.089
R56633 vdd.n21757 vdd.n21756 0.089
R56634 vdd.n10223 vdd.n10132 0.089
R56635 vdd.n16679 vdd.n16599 0.089
R56636 vdd.n24996 vdd.n24994 0.088
R56637 vdd.n11759 vdd.n11758 0.088
R56638 vdd.n21839 vdd.n21838 0.088
R56639 vdd.n458 vdd.n457 0.088
R56640 vdd.n3850 vdd.n3849 0.088
R56641 vdd.n33444 vdd.n33443 0.087
R56642 vdd.n763 vdd.n762 0.087
R56643 vdd.n11754 vdd.n11753 0.087
R56644 vdd.n21834 vdd.n21833 0.087
R56645 vdd.n31033 vdd.n31032 0.087
R56646 vdd.n31043 vdd.n31042 0.087
R56647 vdd.n31948 vdd.n31943 0.087
R56648 vdd.n32293 vdd.n32289 0.087
R56649 vdd.n32310 vdd.n31518 0.087
R56650 vdd.n24621 vdd.n24620 0.087
R56651 vdd.n24898 vdd.n24897 0.086
R56652 vdd.n24930 vdd.n24928 0.086
R56653 vdd.n24918 vdd.n24917 0.086
R56654 vdd.n31517 vdd.n31514 0.085
R56655 vdd.n10257 vdd.n10255 0.085
R56656 vdd.n11870 vdd.n11807 0.085
R56657 vdd.n21961 vdd.n21898 0.085
R56658 vdd.n11786 vdd.n11785 0.084
R56659 vdd.n25828 vdd.n25819 0.084
R56660 vdd.n960 vdd.n958 0.084
R56661 vdd.n11892 vdd.n11891 0.084
R56662 vdd.n21983 vdd.n21982 0.084
R56663 vdd.n27468 vdd.n27467 0.084
R56664 vdd.n27360 vdd.n27359 0.084
R56665 vdd.n27591 vdd.n27583 0.083
R56666 vdd.n25797 vdd.n25786 0.083
R56667 vdd.n26032 vdd.n26023 0.083
R56668 vdd.n25929 vdd.n25920 0.083
R56669 vdd.n25837 vdd.n25830 0.083
R56670 vdd.n25815 vdd.n25814 0.083
R56671 vdd.n11811 vdd.n11808 0.082
R56672 vdd.n21902 vdd.n21899 0.082
R56673 vdd.n10134 vdd.n10068 0.082
R56674 vdd.n25902 vdd.n25892 0.081
R56675 vdd.n25994 vdd.n25984 0.081
R56676 vdd.n1750 vdd.n1748 0.081
R56677 vdd.n1748 vdd.n1730 0.081
R56678 vdd.n11712 vdd.n11699 0.081
R56679 vdd.n11712 vdd.n11711 0.081
R56680 vdd.n11857 vdd.n11856 0.081
R56681 vdd.n11856 vdd.n11839 0.081
R56682 vdd.n21791 vdd.n21789 0.081
R56683 vdd.n21789 vdd.n21785 0.081
R56684 vdd.n21948 vdd.n21947 0.081
R56685 vdd.n21947 vdd.n21930 0.081
R56686 vdd.n25646 vdd.n25405 0.081
R56687 vdd.n25785 vdd.n25775 0.08
R56688 vdd.n35423 vdd.n35418 0.08
R56689 vdd.n34827 vdd.n34822 0.08
R56690 vdd.n5574 vdd.n5569 0.08
R56691 vdd.n4400 vdd.n4395 0.08
R56692 vdd.n24557 vdd.n24556 0.08
R56693 vdd.n34051 vdd.n34050 0.08
R56694 vdd.n35487 vdd.n35486 0.08
R56695 vdd.n34962 vdd.n34961 0.08
R56696 vdd.n34625 vdd.n34624 0.08
R56697 vdd.n5709 vdd.n5708 0.08
R56698 vdd.n5372 vdd.n5371 0.08
R56699 vdd.n5166 vdd.n5068 0.08
R56700 vdd.n4927 vdd.n4877 0.08
R56701 vdd.n4536 vdd.n4535 0.08
R56702 vdd.n25663 vdd.n25662 0.079
R56703 vdd.n30508 vdd.n30507 0.079
R56704 vdd.n24881 vdd.n24859 0.079
R56705 vdd.n27345 vdd.n27334 0.079
R56706 vdd.n27385 vdd.n27376 0.079
R56707 vdd.n27363 vdd.n27362 0.078
R56708 vdd.n10265 vdd.n10123 0.078
R56709 vdd.n15053 vdd.n15052 0.078
R56710 vdd.n35858 vdd.n35848 0.078
R56711 vdd.n26429 vdd.n26420 0.078
R56712 vdd.n31805 vdd.n31729 0.078
R56713 vdd.n12478 vdd.n10601 0.078
R56714 vdd.n10684 vdd.n10683 0.078
R56715 vdd.n12376 vdd.n12375 0.078
R56716 vdd.n12331 vdd.n10851 0.078
R56717 vdd.n10946 vdd.n10945 0.078
R56718 vdd.n11032 vdd.n11017 0.078
R56719 vdd.n11113 vdd.n11091 0.078
R56720 vdd.n12127 vdd.n12126 0.078
R56721 vdd.n12077 vdd.n11267 0.078
R56722 vdd.n12025 vdd.n11360 0.078
R56723 vdd.n11764 vdd.n11678 0.078
R56724 vdd.n24190 vdd.n24188 0.078
R56725 vdd.n24176 vdd.n24174 0.078
R56726 vdd.n24162 vdd.n24160 0.078
R56727 vdd.n24148 vdd.n24146 0.078
R56728 vdd.n24134 vdd.n24132 0.078
R56729 vdd.n24120 vdd.n24118 0.078
R56730 vdd.n24106 vdd.n24104 0.078
R56731 vdd.n24078 vdd.n24068 0.078
R56732 vdd.n24064 vdd.n24054 0.078
R56733 vdd.n24050 vdd.n24040 0.078
R56734 vdd.n24036 vdd.n24026 0.078
R56735 vdd.n24022 vdd.n24012 0.078
R56736 vdd.n24008 vdd.n23998 0.078
R56737 vdd.n23994 vdd.n23984 0.078
R56738 vdd.n23958 vdd.n23956 0.078
R56739 vdd.n23944 vdd.n23942 0.078
R56740 vdd.n23930 vdd.n23928 0.078
R56741 vdd.n23916 vdd.n23914 0.078
R56742 vdd.n23902 vdd.n23900 0.078
R56743 vdd.n23888 vdd.n23886 0.078
R56744 vdd.n23874 vdd.n23872 0.078
R56745 vdd.n23846 vdd.n23836 0.078
R56746 vdd.n23832 vdd.n23822 0.078
R56747 vdd.n23818 vdd.n23808 0.078
R56748 vdd.n23804 vdd.n23794 0.078
R56749 vdd.n23790 vdd.n23780 0.078
R56750 vdd.n23776 vdd.n23766 0.078
R56751 vdd.n23762 vdd.n23752 0.078
R56752 vdd.n23726 vdd.n23724 0.078
R56753 vdd.n23712 vdd.n23710 0.078
R56754 vdd.n23698 vdd.n23696 0.078
R56755 vdd.n23684 vdd.n23682 0.078
R56756 vdd.n23670 vdd.n23668 0.078
R56757 vdd.n23656 vdd.n23654 0.078
R56758 vdd.n23642 vdd.n23640 0.078
R56759 vdd.n23074 vdd.n23064 0.078
R56760 vdd.n23088 vdd.n23078 0.078
R56761 vdd.n23102 vdd.n23092 0.078
R56762 vdd.n23116 vdd.n23106 0.078
R56763 vdd.n23130 vdd.n23120 0.078
R56764 vdd.n23144 vdd.n23134 0.078
R56765 vdd.n23158 vdd.n23148 0.078
R56766 vdd.n23186 vdd.n23184 0.078
R56767 vdd.n23200 vdd.n23198 0.078
R56768 vdd.n23214 vdd.n23212 0.078
R56769 vdd.n23228 vdd.n23226 0.078
R56770 vdd.n23242 vdd.n23240 0.078
R56771 vdd.n23256 vdd.n23254 0.078
R56772 vdd.n23270 vdd.n23268 0.078
R56773 vdd.n23306 vdd.n23296 0.078
R56774 vdd.n23320 vdd.n23310 0.078
R56775 vdd.n23334 vdd.n23324 0.078
R56776 vdd.n23348 vdd.n23338 0.078
R56777 vdd.n23362 vdd.n23352 0.078
R56778 vdd.n23376 vdd.n23366 0.078
R56779 vdd.n23390 vdd.n23380 0.078
R56780 vdd.n23418 vdd.n23416 0.078
R56781 vdd.n23432 vdd.n23430 0.078
R56782 vdd.n23446 vdd.n23444 0.078
R56783 vdd.n23460 vdd.n23458 0.078
R56784 vdd.n23474 vdd.n23472 0.078
R56785 vdd.n23488 vdd.n23486 0.078
R56786 vdd.n23502 vdd.n23500 0.078
R56787 vdd.n23538 vdd.n23528 0.078
R56788 vdd.n23552 vdd.n23542 0.078
R56789 vdd.n23566 vdd.n23556 0.078
R56790 vdd.n23580 vdd.n23570 0.078
R56791 vdd.n23594 vdd.n23584 0.078
R56792 vdd.n23608 vdd.n23598 0.078
R56793 vdd.n23622 vdd.n23612 0.078
R56794 vdd.n22495 vdd.n22485 0.078
R56795 vdd.n22509 vdd.n22499 0.078
R56796 vdd.n22523 vdd.n22513 0.078
R56797 vdd.n22537 vdd.n22527 0.078
R56798 vdd.n22551 vdd.n22541 0.078
R56799 vdd.n22565 vdd.n22555 0.078
R56800 vdd.n22579 vdd.n22569 0.078
R56801 vdd.n22607 vdd.n22605 0.078
R56802 vdd.n22621 vdd.n22619 0.078
R56803 vdd.n22635 vdd.n22633 0.078
R56804 vdd.n22649 vdd.n22647 0.078
R56805 vdd.n22663 vdd.n22661 0.078
R56806 vdd.n22677 vdd.n22675 0.078
R56807 vdd.n22691 vdd.n22689 0.078
R56808 vdd.n22727 vdd.n22717 0.078
R56809 vdd.n22741 vdd.n22731 0.078
R56810 vdd.n22755 vdd.n22745 0.078
R56811 vdd.n22769 vdd.n22759 0.078
R56812 vdd.n22783 vdd.n22773 0.078
R56813 vdd.n22797 vdd.n22787 0.078
R56814 vdd.n22811 vdd.n22801 0.078
R56815 vdd.n22839 vdd.n22837 0.078
R56816 vdd.n22853 vdd.n22851 0.078
R56817 vdd.n22867 vdd.n22865 0.078
R56818 vdd.n22881 vdd.n22879 0.078
R56819 vdd.n22895 vdd.n22893 0.078
R56820 vdd.n22909 vdd.n22907 0.078
R56821 vdd.n22923 vdd.n22921 0.078
R56822 vdd.n22959 vdd.n22949 0.078
R56823 vdd.n22973 vdd.n22963 0.078
R56824 vdd.n22987 vdd.n22977 0.078
R56825 vdd.n23001 vdd.n22991 0.078
R56826 vdd.n23015 vdd.n23005 0.078
R56827 vdd.n23029 vdd.n23019 0.078
R56828 vdd.n23043 vdd.n23033 0.078
R56829 vdd.n16982 vdd.n16981 0.078
R56830 vdd.n17127 vdd.n17109 0.078
R56831 vdd.n17254 vdd.n17253 0.078
R56832 vdd.n17399 vdd.n17381 0.078
R56833 vdd.n17526 vdd.n17525 0.078
R56834 vdd.n17657 vdd.n17639 0.078
R56835 vdd.n17784 vdd.n17783 0.078
R56836 vdd.n17928 vdd.n17910 0.078
R56837 vdd.n18055 vdd.n18054 0.078
R56838 vdd.n18200 vdd.n18182 0.078
R56839 vdd.n21844 vdd.n21841 0.078
R56840 vdd.n24530 vdd.n24529 0.078
R56841 vdd.n27611 vdd.n27607 0.078
R56842 vdd.n27492 vdd.n27488 0.078
R56843 vdd.n27391 vdd.n27387 0.078
R56844 vdd.n25774 vdd.n25766 0.078
R56845 vdd.n27468 vdd.n27279 0.078
R56846 vdd.n27360 vdd.n27302 0.078
R56847 vdd.n25659 vdd.n25652 0.077
R56848 vdd.n26043 vdd.n26034 0.077
R56849 vdd.n25891 vdd.n25883 0.077
R56850 vdd.n25914 vdd.n25725 0.077
R56851 vdd.n25812 vdd.n25754 0.077
R56852 vdd.n31161 vdd.n31132 0.077
R56853 vdd.n25663 vdd.n25404 0.077
R56854 vdd.n25480 vdd.n25479 0.077
R56855 vdd.n11765 vdd.n11677 0.077
R56856 vdd.n21847 vdd.n21846 0.077
R56857 vdd.n27456 vdd.n27446 0.077
R56858 vdd.n25940 vdd.n25931 0.077
R56859 vdd.n25848 vdd.n25839 0.077
R56860 vdd.n27557 vdd.n27547 0.077
R56861 vdd.n25481 vdd.n25480 0.077
R56862 vdd.n25983 vdd.n25973 0.076
R56863 vdd.n38141 vdd.n38139 0.076
R56864 vdd.n25600 vdd.n25598 0.076
R56865 vdd.n24548 vdd.n24547 0.076
R56866 vdd.n25641 vdd.n25633 0.076
R56867 vdd.n26052 vdd.n26045 0.076
R56868 vdd.n34331 vdd.n34328 0.076
R56869 vdd.n34213 vdd.n34159 0.076
R56870 vdd.n35597 vdd.n35594 0.076
R56871 vdd.n35333 vdd.n35279 0.076
R56872 vdd.n35009 vdd.n35006 0.076
R56873 vdd.n34749 vdd.n34695 0.076
R56874 vdd.n6032 vdd.n6029 0.076
R56875 vdd.n5914 vdd.n5860 0.076
R56876 vdd.n5756 vdd.n5753 0.076
R56877 vdd.n5496 vdd.n5442 0.076
R56878 vdd.n4696 vdd.n4620 0.076
R56879 vdd.n4586 vdd.n4583 0.076
R56880 vdd.n4323 vdd.n4269 0.076
R56881 vdd.n25882 vdd.n25874 0.076
R56882 vdd.n25765 vdd.n25760 0.076
R56883 vdd.n27333 vdd.n27323 0.075
R56884 vdd.n25507 vdd.n25497 0.075
R56885 vdd.n25581 vdd.n25571 0.075
R56886 vdd.n25625 vdd.n25616 0.075
R56887 vdd.n25547 vdd.n25538 0.075
R56888 vdd.n25461 vdd.n25454 0.075
R56889 vdd.n32016 vdd.n32015 0.075
R56890 vdd.n32034 vdd.n32033 0.075
R56891 vdd.n32348 vdd.n32347 0.075
R56892 vdd.n32375 vdd.n32374 0.075
R56893 vdd.n31729 vdd.n31727 0.075
R56894 vdd.n31781 vdd.n31780 0.075
R56895 vdd.n26297 vdd.n26293 0.075
R56896 vdd.n26337 vdd.n26324 0.075
R56897 vdd.n12577 vdd.n10256 0.075
R56898 vdd.n15066 vdd.n15063 0.075
R56899 vdd.n24548 vdd.n24545 0.075
R56900 vdd.n2535 vdd.n2534 0.075
R56901 vdd.n25947 vdd.n25942 0.074
R56902 vdd.n25873 vdd.n25867 0.074
R56903 vdd.n26059 vdd.n26054 0.074
R56904 vdd.n25972 vdd.n25964 0.074
R56905 vdd.n31824 vdd.n31710 0.074
R56906 vdd.n11902 vdd.n11901 0.074
R56907 vdd.n21993 vdd.n21992 0.074
R56908 vdd.n25856 vdd.n25850 0.074
R56909 vdd.n1218 vdd.n1217 0.074
R56910 vdd.n27622 vdd.n27613 0.074
R56911 vdd.n31490 vdd.n31478 0.074
R56912 vdd.n31490 vdd.n31480 0.074
R56913 vdd.n31642 vdd.n31637 0.074
R56914 vdd.n31642 vdd.n31638 0.074
R56915 vdd.n26212 vdd.n26201 0.074
R56916 vdd.n26212 vdd.n26202 0.074
R56917 vdd.n26062 vdd.n26061 0.073
R56918 vdd.n25953 vdd.n25949 0.073
R56919 vdd.n25963 vdd.n25957 0.073
R56920 vdd.n25866 vdd.n25860 0.073
R56921 vdd.n27445 vdd.n27437 0.073
R56922 vdd.n27322 vdd.n27314 0.073
R56923 vdd.n10201 vdd.n10088 0.073
R56924 vdd.n10208 vdd.n10078 0.073
R56925 vdd.n10213 vdd.n10093 0.073
R56926 vdd.n10218 vdd.n10067 0.073
R56927 vdd.n12577 vdd.n10255 0.073
R56928 vdd.n16736 vdd.n16732 0.073
R56929 vdd.n10224 vdd.n10223 0.073
R56930 vdd.n16679 vdd.n16670 0.073
R56931 vdd.n27503 vdd.n27494 0.073
R56932 vdd.n27402 vdd.n27393 0.073
R56933 vdd.n842 vdd.n835 0.072
R56934 vdd.n27546 vdd.n27536 0.072
R56935 vdd.n30629 vdd.n30223 0.072
R56936 vdd.n31377 vdd.n31376 0.072
R56937 vdd.n11776 vdd.n11775 0.072
R56938 vdd.n11871 vdd.n11805 0.072
R56939 vdd.n11908 vdd.n11907 0.072
R56940 vdd.n21868 vdd.n21867 0.072
R56941 vdd.n21962 vdd.n21896 0.072
R56942 vdd.n25454 vdd.n25453 0.072
R56943 vdd.n27631 vdd.n27624 0.071
R56944 vdd.n27436 vdd.n27428 0.071
R56945 vdd.n27313 vdd.n27308 0.071
R56946 vdd.n33445 vdd.n33442 0.071
R56947 vdd.n764 vdd.n761 0.071
R56948 vdd.n948 vdd.n921 0.071
R56949 vdd.n459 vdd.n456 0.071
R56950 vdd.n176 vdd.n89 0.071
R56951 vdd.n371 vdd.n320 0.071
R56952 vdd.n25538 vdd.n25537 0.071
R56953 vdd.n31180 vdd.n31175 0.071
R56954 vdd.n31319 vdd.n31308 0.071
R56955 vdd.n12583 vdd.n10124 0.071
R56956 vdd.n12600 vdd.n10075 0.071
R56957 vdd.n16743 vdd.n16680 0.071
R56958 vdd.n25473 vdd.n25469 0.071
R56959 vdd.n27427 vdd.n27421 0.07
R56960 vdd.n27638 vdd.n27633 0.07
R56961 vdd.n27510 vdd.n27505 0.07
R56962 vdd.n27535 vdd.n27527 0.07
R56963 vdd.n38139 vdd.n38114 0.07
R56964 vdd.n11757 vdd.n11756 0.07
R56965 vdd.n21837 vdd.n21836 0.07
R56966 vdd.n27410 vdd.n27404 0.07
R56967 vdd.n27526 vdd.n27520 0.069
R56968 vdd.n27516 vdd.n27512 0.069
R56969 vdd.n33435 vdd.n33405 0.069
R56970 vdd.n33569 vdd.n33483 0.069
R56971 vdd.n33537 vdd.n33534 0.069
R56972 vdd.n34412 vdd.n34396 0.069
R56973 vdd.n34409 vdd.n34402 0.069
R56974 vdd.n34031 vdd.n34003 0.069
R56975 vdd.n35193 vdd.n35165 0.069
R56976 vdd.n35430 vdd.n35417 0.069
R56977 vdd.n35436 vdd.n35412 0.069
R56978 vdd.n34839 vdd.n34816 0.069
R56979 vdd.n34834 vdd.n34821 0.069
R56980 vdd.n34613 vdd.n34585 0.069
R56981 vdd.n755 vdd.n726 0.069
R56982 vdd.n1046 vdd.n968 0.069
R56983 vdd.n69 vdd.n36 0.069
R56984 vdd.n440 vdd.n437 0.069
R56985 vdd.n298 vdd.n234 0.069
R56986 vdd.n6324 vdd.n6296 0.069
R56987 vdd.n6116 vdd.n6109 0.069
R56988 vdd.n5586 vdd.n5563 0.069
R56989 vdd.n5581 vdd.n5568 0.069
R56990 vdd.n5360 vdd.n5332 0.069
R56991 vdd.n4908 vdd.n4903 0.069
R56992 vdd.n5126 vdd.n5123 0.069
R56993 vdd.n4871 vdd.n4807 0.069
R56994 vdd.n4742 vdd.n4739 0.069
R56995 vdd.n4733 vdd.n4731 0.069
R56996 vdd.n4413 vdd.n4389 0.069
R56997 vdd.n4407 vdd.n4394 0.069
R56998 vdd.n4191 vdd.n4163 0.069
R56999 vdd.n27470 vdd.n27273 0.069
R57000 vdd.n27526 vdd.n27524 0.069
R57001 vdd.n27582 vdd.n27580 0.069
R57002 vdd.n27591 vdd.n27589 0.069
R57003 vdd.n27420 vdd.n27418 0.069
R57004 vdd.n27427 vdd.n27425 0.069
R57005 vdd.n27313 vdd.n27311 0.069
R57006 vdd.n25916 vdd.n25719 0.069
R57007 vdd.n25963 vdd.n25961 0.069
R57008 vdd.n25998 vdd.n25693 0.069
R57009 vdd.n26007 vdd.n26005 0.069
R57010 vdd.n25866 vdd.n25864 0.069
R57011 vdd.n25873 vdd.n25871 0.069
R57012 vdd.n25765 vdd.n25763 0.069
R57013 vdd.n14494 ldomc_0.otaldom_0.vdd 0.069
R57014 bandgapmd_0.otam_1.vdd vdd.n19969 0.069
R57015 vdd.n25048 vdd.n24991 0.069
R57016 vdd.n31777 vdd.n31776 0.069
R57017 vdd.n27641 vdd.n27640 0.068
R57018 vdd.n27420 vdd.n27414 0.068
R57019 vdd.n31326 vdd.n31322 0.068
R57020 vdd.n31302 vdd.n31291 0.068
R57021 vdd.n11895 vdd.n11794 0.068
R57022 vdd.n21986 vdd.n21885 0.068
R57023 vdd.n25262 vdd.n25259 0.068
R57024 vdd.n33353 vdd.n33292 0.068
R57025 vdd.n33677 vdd.n33577 0.068
R57026 vdd.n33844 vdd.n33795 0.068
R57027 vdd.n671 vdd.n602 0.068
R57028 vdd.n1142 vdd.n1053 0.068
R57029 vdd.n563 vdd.n510 0.068
R57030 vdd.n33376 vdd.n33375 0.068
R57031 vdd.n690 vdd.n689 0.068
R57032 vdd.n2750 vdd.n2743 0.067
R57033 vdd.n24533 vdd.n24531 0.067
R57034 vdd.n24566 vdd.n24565 0.067
R57035 vdd.n24567 vdd.n24566 0.066
R57036 vdd.n33337 vdd.n33334 0.066
R57037 vdd.n33718 vdd.n33717 0.066
R57038 vdd.n34083 vdd.n34082 0.066
R57039 vdd.n33938 vdd.n33919 0.066
R57040 vdd.n35242 vdd.n35241 0.066
R57041 vdd.n35068 vdd.n35065 0.066
R57042 vdd.n34655 vdd.n34654 0.066
R57043 vdd.n34481 vdd.n34478 0.066
R57044 vdd.n666 vdd.n623 0.066
R57045 vdd.n912 vdd.n911 0.066
R57046 vdd.n555 vdd.n525 0.066
R57047 vdd.n60 vdd.n54 0.066
R57048 vdd.n264 vdd.n263 0.066
R57049 vdd.n5785 vdd.n5784 0.066
R57050 vdd.n6222 vdd.n6193 0.066
R57051 vdd.n5402 vdd.n5401 0.066
R57052 vdd.n5228 vdd.n5225 0.066
R57053 vdd.n5022 vdd.n4996 0.066
R57054 vdd.n4232 vdd.n4231 0.066
R57055 vdd.n4058 vdd.n4055 0.066
R57056 vdd.n27535 vdd.n27533 0.066
R57057 vdd.n25972 vdd.n25970 0.066
R57058 vdd.n24968 vdd.n24966 0.066
R57059 vdd.n33506 vdd.n33505 0.065
R57060 vdd.n1030 vdd.n1029 0.065
R57061 vdd.n33552 vdd.n33514 0.065
R57062 vdd.n35098 vdd.n35045 0.065
R57063 vdd.n69 vdd.n38 0.065
R57064 vdd.n6244 vdd.n6243 0.065
R57065 vdd.n24939 vdd.n24938 0.065
R57066 vdd.n24865 vdd.n24864 0.065
R57067 vdd.n10132 vdd.n10131 0.065
R57068 vdd.n16599 vdd.n16598 0.065
R57069 vdd.n27387 vdd.n27386 0.064
R57070 vdd.n35452 vdd.n35391 0.064
R57071 vdd.n6128 vdd.n6126 0.064
R57072 vdd.n4088 vdd.n4025 0.064
R57073 vdd.n27569 vdd.n27568 0.064
R57074 vdd.n27482 vdd.n27481 0.064
R57075 vdd.n10262 vdd.n10124 0.064
R57076 vdd.n15058 vdd.n15057 0.064
R57077 vdd.n25633 vdd.n25632 0.064
R57078 vdd.n34436 vdd.n34368 0.064
R57079 vdd.n35458 vdd.n35455 0.064
R57080 vdd.n34869 vdd.n34866 0.064
R57081 vdd.n488 vdd.n487 0.064
R57082 vdd.n6131 vdd.n6074 0.064
R57083 vdd.n5616 vdd.n5613 0.064
R57084 vdd.n4787 vdd.n4712 0.064
R57085 vdd.n4443 vdd.n4440 0.064
R57086 vdd.n35499 vdd.n35498 0.063
R57087 vdd.n34947 vdd.n34946 0.063
R57088 vdd.n6000 vdd.n5999 0.063
R57089 vdd.n5694 vdd.n5693 0.063
R57090 vdd.n4521 vdd.n4520 0.063
R57091 vdd.n11879 vdd.n11803 0.063
R57092 vdd.n21970 vdd.n21894 0.063
R57093 vdd.n24559 vdd.n24558 0.063
R57094 vdd.n12600 vdd.n10068 0.063
R57095 vdd.n16743 vdd.n16583 0.063
R57096 vdd.n33429 vdd.n33412 0.062
R57097 vdd.n33543 vdd.n33530 0.062
R57098 vdd.n34150 vdd.n34090 0.062
R57099 vdd.n33959 vdd.n33956 0.062
R57100 vdd.n34036 vdd.n33998 0.062
R57101 vdd.n35198 vdd.n35160 0.062
R57102 vdd.n35272 vdd.n35251 0.062
R57103 vdd.n34688 vdd.n34664 0.062
R57104 vdd.n34511 vdd.n34458 0.062
R57105 vdd.n34616 vdd.n34578 0.062
R57106 vdd.n752 vdd.n736 0.062
R57107 vdd.n1019 vdd.n1013 0.062
R57108 vdd.n1037 vdd.n1027 0.062
R57109 vdd.n86 vdd.n6 0.062
R57110 vdd.n430 vdd.n427 0.062
R57111 vdd.n227 vdd.n226 0.062
R57112 vdd.n160 vdd.n157 0.062
R57113 vdd.n6327 vdd.n6289 0.062
R57114 vdd.n5836 vdd.n5792 0.062
R57115 vdd.n5435 vdd.n5411 0.062
R57116 vdd.n5258 vdd.n5205 0.062
R57117 vdd.n5363 vdd.n5325 0.062
R57118 vdd.n5137 vdd.n5134 0.062
R57119 vdd.n5048 vdd.n4971 0.062
R57120 vdd.n4262 vdd.n4241 0.062
R57121 vdd.n4088 vdd.n4035 0.062
R57122 vdd.n4437 vdd.n4367 0.062
R57123 vdd.n4194 vdd.n4156 0.062
R57124 vdd.n1915 vdd.n1209 0.062
R57125 vdd.n31052 vdd.n31049 0.062
R57126 vdd.n32300 vdd.n31528 0.062
R57127 vdd.n27569 vdd.n27567 0.062
R57128 vdd.n25996 vdd.n25703 0.062
R57129 vdd.n30707 vdd.n30706 0.062
R57130 vdd.n26483 vdd.n26482 0.062
R57131 vdd.n26548 vdd.n26544 0.062
R57132 vdd.n3943 vdd.n3783 0.062
R57133 vdd.n3930 vdd.n3791 0.062
R57134 vdd.n2540 vdd.n2427 0.062
R57135 vdd.n31707 vdd.n31706 0.062
R57136 vdd.n13948 vdd.n8598 0.062
R57137 vdd.n14150 vdd.n8495 0.062
R57138 vdd.n14150 vdd.n14149 0.062
R57139 vdd.n14238 vdd.n8376 0.062
R57140 vdd.n14416 vdd.n14412 0.062
R57141 vdd.n14416 vdd.n14415 0.062
R57142 vdd.n14608 vdd.n14607 0.062
R57143 vdd.n9183 vdd.n9154 0.062
R57144 vdd.n13280 vdd.n9154 0.062
R57145 vdd.n13385 vdd.n13384 0.062
R57146 vdd.n8962 vdd.n8933 0.062
R57147 vdd.n13572 vdd.n8933 0.062
R57148 vdd.n13677 vdd.n13676 0.062
R57149 vdd.n10448 vdd.n10447 0.062
R57150 vdd.n10447 vdd.n10293 0.062
R57151 vdd.n10350 vdd.n10349 0.062
R57152 vdd.n9350 vdd.n9349 0.062
R57153 vdd.n13038 vdd.n9350 0.062
R57154 vdd.n9448 vdd.n9447 0.062
R57155 vdd.n12940 vdd.n9515 0.062
R57156 vdd.n9533 vdd.n9515 0.062
R57157 vdd.n9634 vdd.n9603 0.062
R57158 vdd.n9710 vdd.n9709 0.062
R57159 vdd.n12830 vdd.n9710 0.062
R57160 vdd.n9807 vdd.n9806 0.062
R57161 vdd.n12732 vdd.n9875 0.062
R57162 vdd.n9894 vdd.n9875 0.062
R57163 vdd.n9994 vdd.n9963 0.062
R57164 vdd.n19020 vdd.n19019 0.062
R57165 vdd.n18906 vdd.n18894 0.062
R57166 vdd.n18894 vdd.n18888 0.062
R57167 vdd.n18761 vdd.n18760 0.062
R57168 vdd.n18647 vdd.n18635 0.062
R57169 vdd.n18635 vdd.n18629 0.062
R57170 vdd.n18502 vdd.n18501 0.062
R57171 vdd.n21531 vdd.n21519 0.062
R57172 vdd.n21519 vdd.n21513 0.062
R57173 vdd.n21386 vdd.n21385 0.062
R57174 vdd.n21272 vdd.n21260 0.062
R57175 vdd.n21260 vdd.n21254 0.062
R57176 vdd.n21127 vdd.n21126 0.062
R57177 vdd.n15313 vdd.n15309 0.062
R57178 vdd.n15314 vdd.n15313 0.062
R57179 vdd.n15418 vdd.n15417 0.062
R57180 vdd.n15541 vdd.n15537 0.062
R57181 vdd.n15542 vdd.n15541 0.062
R57182 vdd.n15668 vdd.n15667 0.062
R57183 vdd.n15797 vdd.n15793 0.062
R57184 vdd.n15798 vdd.n15797 0.062
R57185 vdd.n15924 vdd.n15923 0.062
R57186 vdd.n16053 vdd.n16049 0.062
R57187 vdd.n16054 vdd.n16053 0.062
R57188 vdd.n16180 vdd.n16179 0.062
R57189 vdd.n16309 vdd.n16305 0.062
R57190 vdd.n16310 vdd.n16309 0.062
R57191 vdd.n16436 vdd.n16435 0.062
R57192 vdd.n24968 vdd.n24967 0.062
R57193 vdd.n24880 vdd.n24876 0.062
R57194 vdd.n24968 vdd.n24965 0.062
R57195 vdd.n11906 vdd.n11788 0.062
R57196 vdd.n21997 vdd.n21879 0.062
R57197 vdd.n27363 vdd.n27296 0.061
R57198 vdd.n1037 vdd.n1024 0.061
R57199 vdd.n69 vdd.n68 0.061
R57200 vdd.n11707 vdd.n11706 0.061
R57201 vdd.n11850 vdd.n11849 0.061
R57202 vdd.n21781 vdd.n21778 0.061
R57203 vdd.n21941 vdd.n21940 0.061
R57204 vdd.n25815 vdd.n25748 0.061
R57205 vdd.n11771 vdd.n11665 0.061
R57206 vdd.n11876 vdd.n11875 0.061
R57207 vdd.n21866 vdd.n21865 0.061
R57208 vdd.n21967 vdd.n21966 0.061
R57209 vdd.n32090 vdd.n32089 0.061
R57210 vdd.n32513 vdd.n32512 0.061
R57211 vdd.n25587 vdd.n25586 0.061
R57212 vdd.n25555 vdd.n25554 0.061
R57213 vdd.n25469 vdd.n25468 0.061
R57214 vdd.n35314 vdd.n35306 0.06
R57215 vdd.n5870 vdd.n5869 0.06
R57216 vdd.n33959 vdd.n33958 0.06
R57217 vdd.n34511 vdd.n34448 0.06
R57218 vdd.n5258 vdd.n5195 0.06
R57219 vdd.n4771 vdd.n4715 0.06
R57220 vdd.n25918 vdd.n25710 0.06
R57221 vdd.n13861 vdd.n13860 0.06
R57222 vdd.n13861 vdd.n8717 0.06
R57223 vdd.n21012 vdd.n19140 0.06
R57224 vdd.n21015 vdd.n21012 0.06
R57225 vdd.n24943 vdd.n24942 0.06
R57226 vdd.n24950 vdd.n24949 0.06
R57227 vdd.n4908 vdd.n4901 0.06
R57228 vdd.n281 vdd.n280 0.06
R57229 vdd.n31784 vdd.n31783 0.06
R57230 vdd.n11746 vdd.n11745 0.06
R57231 vdd.n21828 vdd.n21827 0.06
R57232 vdd.n25652 vdd.n25651 0.06
R57233 vdd.n81 vdd.n78 0.06
R57234 vdd.n27611 vdd.n27610 0.059
R57235 vdd.n27492 vdd.n27491 0.059
R57236 vdd.n27391 vdd.n27390 0.059
R57237 vdd.n25830 vdd.n25829 0.059
R57238 vdd.n34433 vdd.n34423 0.059
R57239 vdd.n33959 vdd.n33946 0.059
R57240 vdd.n34434 vdd.n34433 0.059
R57241 vdd.n35591 vdd.n35590 0.059
R57242 vdd.n35578 vdd.n35577 0.059
R57243 vdd.n35566 vdd.n35565 0.059
R57244 vdd.n35554 vdd.n35553 0.059
R57245 vdd.n35095 vdd.n35094 0.059
R57246 vdd.n35082 vdd.n35081 0.059
R57247 vdd.n35068 vdd.n35067 0.059
R57248 vdd.n35056 vdd.n35055 0.059
R57249 vdd.n35430 vdd.n35429 0.059
R57250 vdd.n35436 vdd.n35435 0.059
R57251 vdd.n35442 vdd.n35441 0.059
R57252 vdd.n35448 vdd.n35447 0.059
R57253 vdd.n35193 vdd.n35192 0.059
R57254 vdd.n35198 vdd.n35197 0.059
R57255 vdd.n35204 vdd.n35203 0.059
R57256 vdd.n35210 vdd.n35209 0.059
R57257 vdd.n35331 vdd.n35282 0.059
R57258 vdd.n35328 vdd.n35294 0.059
R57259 vdd.n35325 vdd.n35305 0.059
R57260 vdd.n34511 vdd.n34510 0.059
R57261 vdd.n34864 vdd.n34863 0.059
R57262 vdd.n34863 vdd.n34793 0.059
R57263 vdd.n1038 vdd.n1037 0.059
R57264 vdd.n6027 vdd.n5929 0.059
R57265 vdd.n6024 vdd.n5940 0.059
R57266 vdd.n6021 vdd.n5949 0.059
R57267 vdd.n6018 vdd.n5958 0.059
R57268 vdd.n6228 vdd.n6164 0.059
R57269 vdd.n6225 vdd.n6175 0.059
R57270 vdd.n6222 vdd.n6186 0.059
R57271 vdd.n6219 vdd.n6195 0.059
R57272 vdd.n6116 vdd.n6111 0.059
R57273 vdd.n6119 vdd.n6103 0.059
R57274 vdd.n6122 vdd.n6092 0.059
R57275 vdd.n6324 vdd.n6298 0.059
R57276 vdd.n6327 vdd.n6291 0.059
R57277 vdd.n6330 vdd.n6281 0.059
R57278 vdd.n6333 vdd.n6269 0.059
R57279 vdd.n5911 vdd.n5910 0.059
R57280 vdd.n5897 vdd.n5896 0.059
R57281 vdd.n5883 vdd.n5874 0.059
R57282 vdd.n5258 vdd.n5257 0.059
R57283 vdd.n5611 vdd.n5610 0.059
R57284 vdd.n5610 vdd.n5540 0.059
R57285 vdd.n25996 vdd.n25995 0.059
R57286 vdd.n25918 vdd.n25917 0.059
R57287 vdd.n25663 vdd.n25398 0.059
R57288 vdd.n10547 vdd.n10539 0.059
R57289 vdd.n10549 vdd.n10534 0.059
R57290 vdd.n12508 vdd.n10560 0.059
R57291 vdd.n12506 vdd.n10561 0.059
R57292 vdd.n12495 vdd.n12494 0.059
R57293 vdd.n10592 vdd.n10570 0.059
R57294 vdd.n12476 vdd.n10602 0.059
R57295 vdd.n12465 vdd.n12464 0.059
R57296 vdd.n10639 vdd.n10634 0.059
R57297 vdd.n10641 vdd.n10630 0.059
R57298 vdd.n12449 vdd.n10652 0.059
R57299 vdd.n12447 vdd.n10653 0.059
R57300 vdd.n12436 vdd.n12435 0.059
R57301 vdd.n10685 vdd.n10677 0.059
R57302 vdd.n12420 vdd.n10696 0.059
R57303 vdd.n12418 vdd.n10697 0.059
R57304 vdd.n12407 vdd.n12406 0.059
R57305 vdd.n10732 vdd.n10705 0.059
R57306 vdd.n10734 vdd.n10725 0.059
R57307 vdd.n12389 vdd.n10745 0.059
R57308 vdd.n12387 vdd.n10746 0.059
R57309 vdd.n10790 vdd.n10785 0.059
R57310 vdd.n10792 vdd.n10781 0.059
R57311 vdd.n12360 vdd.n10803 0.059
R57312 vdd.n12358 vdd.n10804 0.059
R57313 vdd.n12347 vdd.n12346 0.059
R57314 vdd.n10840 vdd.n10836 0.059
R57315 vdd.n10838 vdd.n10830 0.059
R57316 vdd.n12330 vdd.n12329 0.059
R57317 vdd.n10879 vdd.n10855 0.059
R57318 vdd.n10881 vdd.n10872 0.059
R57319 vdd.n12312 vdd.n10892 0.059
R57320 vdd.n12310 vdd.n10893 0.059
R57321 vdd.n12299 vdd.n12298 0.059
R57322 vdd.n10932 vdd.n10902 0.059
R57323 vdd.n10934 vdd.n10926 0.059
R57324 vdd.n10950 vdd.n10949 0.059
R57325 vdd.n10977 vdd.n10972 0.059
R57326 vdd.n10979 vdd.n10967 0.059
R57327 vdd.n12259 vdd.n10990 0.059
R57328 vdd.n12257 vdd.n10991 0.059
R57329 vdd.n12246 vdd.n12245 0.059
R57330 vdd.n11025 vdd.n11023 0.059
R57331 vdd.n12229 vdd.n11033 0.059
R57332 vdd.n12227 vdd.n11034 0.059
R57333 vdd.n12216 vdd.n12215 0.059
R57334 vdd.n11069 vdd.n11042 0.059
R57335 vdd.n11071 vdd.n11062 0.059
R57336 vdd.n12198 vdd.n11082 0.059
R57337 vdd.n12196 vdd.n11083 0.059
R57338 vdd.n12185 vdd.n12184 0.059
R57339 vdd.n12169 vdd.n11124 0.059
R57340 vdd.n12167 vdd.n11125 0.059
R57341 vdd.n12156 vdd.n12155 0.059
R57342 vdd.n11162 vdd.n11157 0.059
R57343 vdd.n11164 vdd.n11153 0.059
R57344 vdd.n12140 vdd.n11174 0.059
R57345 vdd.n12138 vdd.n11175 0.059
R57346 vdd.n11204 vdd.n11180 0.059
R57347 vdd.n11206 vdd.n11197 0.059
R57348 vdd.n12110 vdd.n11217 0.059
R57349 vdd.n12108 vdd.n11218 0.059
R57350 vdd.n12097 vdd.n12096 0.059
R57351 vdd.n11253 vdd.n11227 0.059
R57352 vdd.n11255 vdd.n11246 0.059
R57353 vdd.n12079 vdd.n11266 0.059
R57354 vdd.n11299 vdd.n11294 0.059
R57355 vdd.n11301 vdd.n11289 0.059
R57356 vdd.n12054 vdd.n11312 0.059
R57357 vdd.n12052 vdd.n11313 0.059
R57358 vdd.n12041 vdd.n12040 0.059
R57359 vdd.n11349 vdd.n11345 0.059
R57360 vdd.n11347 vdd.n11339 0.059
R57361 vdd.n12024 vdd.n12023 0.059
R57362 vdd.n11388 vdd.n11364 0.059
R57363 vdd.n11390 vdd.n11381 0.059
R57364 vdd.n12006 vdd.n11401 0.059
R57365 vdd.n12004 vdd.n11402 0.059
R57366 vdd.n11993 vdd.n11992 0.059
R57367 vdd.n11476 vdd.n11411 0.059
R57368 vdd.n16889 vdd.n16888 0.059
R57369 vdd.n16905 vdd.n16904 0.059
R57370 vdd.n16921 vdd.n16920 0.059
R57371 vdd.n16937 vdd.n16936 0.059
R57372 vdd.n16953 vdd.n16952 0.059
R57373 vdd.n16969 vdd.n16968 0.059
R57374 vdd.n16998 vdd.n16997 0.059
R57375 vdd.n17014 vdd.n17013 0.059
R57376 vdd.n17030 vdd.n17029 0.059
R57377 vdd.n17046 vdd.n17045 0.059
R57378 vdd.n17062 vdd.n17061 0.059
R57379 vdd.n17078 vdd.n17077 0.059
R57380 vdd.n17094 vdd.n17093 0.059
R57381 vdd.n17129 vdd.n17128 0.059
R57382 vdd.n17145 vdd.n17144 0.059
R57383 vdd.n17161 vdd.n17160 0.059
R57384 vdd.n17177 vdd.n17176 0.059
R57385 vdd.n17193 vdd.n17192 0.059
R57386 vdd.n17209 vdd.n17208 0.059
R57387 vdd.n17225 vdd.n17224 0.059
R57388 vdd.n17241 vdd.n17240 0.059
R57389 vdd.n17270 vdd.n17269 0.059
R57390 vdd.n17286 vdd.n17285 0.059
R57391 vdd.n17302 vdd.n17301 0.059
R57392 vdd.n17318 vdd.n17317 0.059
R57393 vdd.n17334 vdd.n17333 0.059
R57394 vdd.n17350 vdd.n17349 0.059
R57395 vdd.n17366 vdd.n17365 0.059
R57396 vdd.n17401 vdd.n17400 0.059
R57397 vdd.n17417 vdd.n17416 0.059
R57398 vdd.n17433 vdd.n17432 0.059
R57399 vdd.n17449 vdd.n17448 0.059
R57400 vdd.n17465 vdd.n17464 0.059
R57401 vdd.n17481 vdd.n17480 0.059
R57402 vdd.n17497 vdd.n17496 0.059
R57403 vdd.n17513 vdd.n17512 0.059
R57404 vdd.n17542 vdd.n17541 0.059
R57405 vdd.n17558 vdd.n17557 0.059
R57406 vdd.n17574 vdd.n17573 0.059
R57407 vdd.n17590 vdd.n17589 0.059
R57408 vdd.n17591 vdd.n16819 0.059
R57409 vdd.n17608 vdd.n17607 0.059
R57410 vdd.n17624 vdd.n17623 0.059
R57411 vdd.n17659 vdd.n17658 0.059
R57412 vdd.n17675 vdd.n17674 0.059
R57413 vdd.n17691 vdd.n17690 0.059
R57414 vdd.n17707 vdd.n17706 0.059
R57415 vdd.n17723 vdd.n17722 0.059
R57416 vdd.n17739 vdd.n17738 0.059
R57417 vdd.n17755 vdd.n17754 0.059
R57418 vdd.n17771 vdd.n17770 0.059
R57419 vdd.n17800 vdd.n17799 0.059
R57420 vdd.n17816 vdd.n17815 0.059
R57421 vdd.n17832 vdd.n17831 0.059
R57422 vdd.n17848 vdd.n17847 0.059
R57423 vdd.n17864 vdd.n17863 0.059
R57424 vdd.n17879 vdd.n17878 0.059
R57425 vdd.n17895 vdd.n17894 0.059
R57426 vdd.n17930 vdd.n17929 0.059
R57427 vdd.n17946 vdd.n17945 0.059
R57428 vdd.n17962 vdd.n17961 0.059
R57429 vdd.n17978 vdd.n17977 0.059
R57430 vdd.n17994 vdd.n17993 0.059
R57431 vdd.n18010 vdd.n18009 0.059
R57432 vdd.n18026 vdd.n18025 0.059
R57433 vdd.n18042 vdd.n18041 0.059
R57434 vdd.n18071 vdd.n18070 0.059
R57435 vdd.n18087 vdd.n18086 0.059
R57436 vdd.n18103 vdd.n18102 0.059
R57437 vdd.n18119 vdd.n18118 0.059
R57438 vdd.n18135 vdd.n18134 0.059
R57439 vdd.n18151 vdd.n18150 0.059
R57440 vdd.n18167 vdd.n18166 0.059
R57441 vdd.n18202 vdd.n18201 0.059
R57442 vdd.n18218 vdd.n18217 0.059
R57443 vdd.n18233 vdd.n18232 0.059
R57444 vdd.n18248 vdd.n18247 0.059
R57445 vdd.n18263 vdd.n18262 0.059
R57446 vdd.n18278 vdd.n18277 0.059
R57447 vdd.n18293 vdd.n18292 0.059
R57448 vdd.n33750 vdd.n33749 0.059
R57449 vdd.n1817 vdd.n1813 0.059
R57450 vdd.n26032 vdd.n26031 0.059
R57451 vdd.n25929 vdd.n25928 0.059
R57452 vdd.n25837 vdd.n25836 0.059
R57453 vdd.n4312 vdd.n4304 0.058
R57454 vdd.n10238 vdd.n10236 0.058
R57455 vdd.n16668 vdd.n16665 0.058
R57456 vdd.n33325 vdd.n33322 0.058
R57457 vdd.n33552 vdd.n33551 0.058
R57458 vdd.n33710 vdd.n33709 0.058
R57459 vdd.n33746 vdd.n33745 0.058
R57460 vdd.n33661 vdd.n33658 0.058
R57461 vdd.n34300 vdd.n34297 0.058
R57462 vdd.n34431 vdd.n34428 0.058
R57463 vdd.n33935 vdd.n33927 0.058
R57464 vdd.n33960 vdd.n33959 0.058
R57465 vdd.n34433 vdd.n34420 0.058
R57466 vdd.n35566 vdd.n35563 0.058
R57467 vdd.n35056 vdd.n35053 0.058
R57468 vdd.n35389 vdd.n35386 0.058
R57469 vdd.n35452 vdd.n35389 0.058
R57470 vdd.n34998 vdd.n34913 0.058
R57471 vdd.n34861 vdd.n34858 0.058
R57472 vdd.n34469 vdd.n34466 0.058
R57473 vdd.n34512 vdd.n34511 0.058
R57474 vdd.n34863 vdd.n34853 0.058
R57475 vdd.n663 vdd.n632 0.058
R57476 vdd.n915 vdd.n914 0.058
R57477 vdd.n1137 vdd.n1074 0.058
R57478 vdd.n549 vdd.n532 0.058
R57479 vdd.n6021 vdd.n5956 0.058
R57480 vdd.n6219 vdd.n6201 0.058
R57481 vdd.n6082 vdd.n6079 0.058
R57482 vdd.n6128 vdd.n6082 0.058
R57483 vdd.n5745 vdd.n5660 0.058
R57484 vdd.n5608 vdd.n5605 0.058
R57485 vdd.n5216 vdd.n5213 0.058
R57486 vdd.n5259 vdd.n5258 0.058
R57487 vdd.n5610 vdd.n5600 0.058
R57488 vdd.n4680 vdd.n4642 0.058
R57489 vdd.n4835 vdd.n4834 0.058
R57490 vdd.n4771 vdd.n4723 0.058
R57491 vdd.n4723 vdd.n4720 0.058
R57492 vdd.n5017 vdd.n5002 0.058
R57493 vdd.n4772 vdd.n4771 0.058
R57494 vdd.n5048 vdd.n5036 0.058
R57495 vdd.n4575 vdd.n4487 0.058
R57496 vdd.n4435 vdd.n4432 0.058
R57497 vdd.n4046 vdd.n4043 0.058
R57498 vdd.n27482 vdd.n27272 0.058
R57499 vdd.n27436 vdd.n27434 0.058
R57500 vdd.n25918 vdd.n25709 0.058
R57501 vdd.n25997 vdd.n25996 0.058
R57502 vdd.n25919 vdd.n25918 0.058
R57503 vdd.n25882 vdd.n25880 0.058
R57504 vdd.n10095 vdd.n10094 0.058
R57505 vdd.n11900 vdd.n11899 0.057
R57506 vdd.n21991 vdd.n21990 0.057
R57507 vdd.n33424 vdd.n33423 0.057
R57508 vdd.n33429 vdd.n33428 0.057
R57509 vdd.n33435 vdd.n33434 0.057
R57510 vdd.n33440 vdd.n33439 0.057
R57511 vdd.n33350 vdd.n33349 0.057
R57512 vdd.n33337 vdd.n33336 0.057
R57513 vdd.n33325 vdd.n33324 0.057
R57514 vdd.n33313 vdd.n33312 0.057
R57515 vdd.n33537 vdd.n33536 0.057
R57516 vdd.n33543 vdd.n33542 0.057
R57517 vdd.n33549 vdd.n33548 0.057
R57518 vdd.n33674 vdd.n33673 0.057
R57519 vdd.n33661 vdd.n33660 0.057
R57520 vdd.n33649 vdd.n33648 0.057
R57521 vdd.n33841 vdd.n33840 0.057
R57522 vdd.n33829 vdd.n33828 0.057
R57523 vdd.n33817 vdd.n33816 0.057
R57524 vdd.n35188 vdd.n35187 0.057
R57525 vdd.n6321 vdd.n6305 0.057
R57526 vdd.n4581 vdd.n4460 0.057
R57527 vdd.n4578 vdd.n4471 0.057
R57528 vdd.n4575 vdd.n4480 0.057
R57529 vdd.n4572 vdd.n4489 0.057
R57530 vdd.n4321 vdd.n4272 0.057
R57531 vdd.n4318 vdd.n4284 0.057
R57532 vdd.n4315 vdd.n4295 0.057
R57533 vdd.n4085 vdd.n4084 0.057
R57534 vdd.n4072 vdd.n4071 0.057
R57535 vdd.n4058 vdd.n4057 0.057
R57536 vdd.n4046 vdd.n4045 0.057
R57537 vdd.n4407 vdd.n4406 0.057
R57538 vdd.n4413 vdd.n4412 0.057
R57539 vdd.n4419 vdd.n4418 0.057
R57540 vdd.n4425 vdd.n4424 0.057
R57541 vdd.n4191 vdd.n4165 0.057
R57542 vdd.n4194 vdd.n4158 0.057
R57543 vdd.n4197 vdd.n4148 0.057
R57544 vdd.n4200 vdd.n4136 0.057
R57545 vdd.n27557 vdd.n27556 0.057
R57546 vdd.n27546 vdd.n27545 0.057
R57547 vdd.n27535 vdd.n27534 0.057
R57548 vdd.n27526 vdd.n27525 0.057
R57549 vdd.n27456 vdd.n27455 0.057
R57550 vdd.n27445 vdd.n27444 0.057
R57551 vdd.n27436 vdd.n27435 0.057
R57552 vdd.n27427 vdd.n27426 0.057
R57553 vdd.n27345 vdd.n27344 0.057
R57554 vdd.n27333 vdd.n27332 0.057
R57555 vdd.n27322 vdd.n27321 0.057
R57556 vdd.n27313 vdd.n27312 0.057
R57557 vdd.n10094 vdd.n10077 0.057
R57558 vdd.n11898 vdd.n11897 0.057
R57559 vdd.n21989 vdd.n21988 0.057
R57560 vdd.n33829 vdd.n33796 0.057
R57561 vdd.n812 vdd.n807 0.057
R57562 vdd.n927 vdd.n926 0.057
R57563 vdd.n33564 vdd.n33561 0.057
R57564 vdd.n34144 vdd.n34141 0.057
R57565 vdd.n35266 vdd.n35263 0.057
R57566 vdd.n34685 vdd.n34679 0.057
R57567 vdd.n1043 vdd.n982 0.057
R57568 vdd.n901 vdd.n900 0.057
R57569 vdd.n503 vdd.n488 0.057
R57570 vdd.n5833 vdd.n5807 0.057
R57571 vdd.n5432 vdd.n5426 0.057
R57572 vdd.n4259 vdd.n4256 0.057
R57573 vdd.n24635 vdd.n24632 0.056
R57574 vdd.n33553 vdd.n33552 0.056
R57575 vdd.n33637 vdd.n33636 0.056
R57576 vdd.n544 vdd.n543 0.056
R57577 vdd.n549 vdd.n548 0.056
R57578 vdd.n555 vdd.n554 0.056
R57579 vdd.n560 vdd.n559 0.056
R57580 vdd.n70 vdd.n69 0.056
R57581 vdd.n453 vdd.n452 0.056
R57582 vdd.n440 vdd.n439 0.056
R57583 vdd.n430 vdd.n429 0.056
R57584 vdd.n418 vdd.n417 0.056
R57585 vdd.n60 vdd.n59 0.056
R57586 vdd.n66 vdd.n65 0.056
R57587 vdd.n173 vdd.n172 0.056
R57588 vdd.n160 vdd.n159 0.056
R57589 vdd.n148 vdd.n147 0.056
R57590 vdd.n136 vdd.n135 0.056
R57591 vdd.n275 vdd.n274 0.056
R57592 vdd.n368 vdd.n367 0.056
R57593 vdd.n354 vdd.n353 0.056
R57594 vdd.n342 vdd.n341 0.056
R57595 vdd.n5164 vdd.n5163 0.056
R57596 vdd.n5151 vdd.n5150 0.056
R57597 vdd.n5137 vdd.n5136 0.056
R57598 vdd.n5126 vdd.n5125 0.056
R57599 vdd.n4848 vdd.n4847 0.056
R57600 vdd.n4771 vdd.n4770 0.056
R57601 vdd.n5049 vdd.n5048 0.056
R57602 vdd.n4768 vdd.n4767 0.056
R57603 vdd.n4755 vdd.n4754 0.056
R57604 vdd.n4742 vdd.n4741 0.056
R57605 vdd.n4733 vdd.n4732 0.056
R57606 vdd.n5017 vdd.n5016 0.056
R57607 vdd.n5022 vdd.n5021 0.056
R57608 vdd.n5028 vdd.n5027 0.056
R57609 vdd.n5034 vdd.n5033 0.056
R57610 vdd.n4675 vdd.n4674 0.056
R57611 vdd.n4680 vdd.n4679 0.056
R57612 vdd.n4686 vdd.n4685 0.056
R57613 vdd.n4691 vdd.n4690 0.056
R57614 vdd.n4925 vdd.n4880 0.056
R57615 vdd.n4922 vdd.n4891 0.056
R57616 vdd.n4919 vdd.n4900 0.056
R57617 vdd.n4088 vdd.n4087 0.056
R57618 vdd.n4438 vdd.n4437 0.056
R57619 vdd.n4188 vdd.n4172 0.056
R57620 vdd.n27482 vdd.n27471 0.056
R57621 vdd.n27591 vdd.n27590 0.056
R57622 vdd.n27420 vdd.n27419 0.056
R57623 vdd.n25581 vdd.n25580 0.056
R57624 vdd.n25507 vdd.n25506 0.056
R57625 vdd.n32245 vdd.n32243 0.056
R57626 vdd.n31187 vdd.n31023 0.056
R57627 vdd.n11751 vdd.n11750 0.056
R57628 vdd.n21822 vdd.n21821 0.056
R57629 vdd.n4908 vdd.n4907 0.056
R57630 vdd.n34169 vdd.n34168 0.055
R57631 vdd.n34738 vdd.n34730 0.055
R57632 vdd.n5485 vdd.n5477 0.055
R57633 vdd.n10263 vdd.n10123 0.055
R57634 vdd.n15053 vdd.n15050 0.055
R57635 vdd.n33591 vdd.n33590 0.055
R57636 vdd.n951 vdd.n950 0.055
R57637 vdd.n33424 vdd.n33417 0.055
R57638 vdd.n33763 vdd.n33727 0.055
R57639 vdd.n34439 vdd.n34352 0.055
R57640 vdd.n35463 vdd.n35370 0.055
R57641 vdd.n35098 vdd.n35097 0.055
R57642 vdd.n35453 vdd.n35452 0.055
R57643 vdd.n34874 vdd.n34780 0.055
R57644 vdd.n749 vdd.n743 0.055
R57645 vdd.n899 vdd.n891 0.055
R57646 vdd.n418 vdd.n415 0.055
R57647 vdd.n148 vdd.n145 0.055
R57648 vdd.n354 vdd.n351 0.055
R57649 vdd.n6134 vdd.n6058 0.055
R57650 vdd.n6244 vdd.n6230 0.055
R57651 vdd.n6129 vdd.n6128 0.055
R57652 vdd.n5621 vdd.n5527 0.055
R57653 vdd.n4868 vdd.n4816 0.055
R57654 vdd.n4799 vdd.n4796 0.055
R57655 vdd.n4448 vdd.n4354 0.055
R57656 vdd.n4089 vdd.n4088 0.055
R57657 vdd.n4437 vdd.n4427 0.055
R57658 vdd.n27570 vdd.n27569 0.055
R57659 vdd.n11889 vdd.n11797 0.055
R57660 vdd.n21980 vdd.n21888 0.055
R57661 vdd.n24955 vdd.n24954 0.055
R57662 vdd.n35490 vdd.n35489 0.055
R57663 vdd.n5818 vdd.n5817 0.055
R57664 vdd.n28802 vdd.n28801 0.055
R57665 vdd.n34169 vdd.n34164 0.054
R57666 vdd.n34738 vdd.n34737 0.054
R57667 vdd.n5485 vdd.n5484 0.054
R57668 vdd.n25481 vdd.n25447 0.054
R57669 vdd.n34325 vdd.n34324 0.054
R57670 vdd.n34312 vdd.n34311 0.054
R57671 vdd.n34300 vdd.n34299 0.054
R57672 vdd.n34288 vdd.n34287 0.054
R57673 vdd.n34130 vdd.n34129 0.054
R57674 vdd.n34210 vdd.n34209 0.054
R57675 vdd.n34196 vdd.n34195 0.054
R57676 vdd.n34182 vdd.n34181 0.054
R57677 vdd.n33944 vdd.n33890 0.054
R57678 vdd.n33941 vdd.n33901 0.054
R57679 vdd.n33938 vdd.n33912 0.054
R57680 vdd.n33935 vdd.n33921 0.054
R57681 vdd.n34409 vdd.n34404 0.054
R57682 vdd.n34412 vdd.n34398 0.054
R57683 vdd.n34415 vdd.n34390 0.054
R57684 vdd.n34418 vdd.n34378 0.054
R57685 vdd.n34031 vdd.n34030 0.054
R57686 vdd.n34036 vdd.n34035 0.054
R57687 vdd.n34042 vdd.n34041 0.054
R57688 vdd.n34047 vdd.n34046 0.054
R57689 vdd.n35543 vdd.n35542 0.054
R57690 vdd.n35099 vdd.n35098 0.054
R57691 vdd.n35452 vdd.n35450 0.054
R57692 vdd.n35004 vdd.n34886 0.054
R57693 vdd.n35001 vdd.n34897 0.054
R57694 vdd.n34998 vdd.n34906 0.054
R57695 vdd.n34995 vdd.n34915 0.054
R57696 vdd.n34747 vdd.n34698 0.054
R57697 vdd.n34744 vdd.n34710 0.054
R57698 vdd.n34741 vdd.n34721 0.054
R57699 vdd.n34508 vdd.n34507 0.054
R57700 vdd.n34495 vdd.n34494 0.054
R57701 vdd.n34481 vdd.n34480 0.054
R57702 vdd.n34469 vdd.n34468 0.054
R57703 vdd.n34834 vdd.n34833 0.054
R57704 vdd.n34839 vdd.n34838 0.054
R57705 vdd.n34845 vdd.n34844 0.054
R57706 vdd.n34851 vdd.n34850 0.054
R57707 vdd.n34613 vdd.n34587 0.054
R57708 vdd.n34616 vdd.n34580 0.054
R57709 vdd.n34619 vdd.n34570 0.054
R57710 vdd.n34622 vdd.n34559 0.054
R57711 vdd.n749 vdd.n745 0.054
R57712 vdd.n752 vdd.n738 0.054
R57713 vdd.n755 vdd.n728 0.054
R57714 vdd.n758 vdd.n721 0.054
R57715 vdd.n669 vdd.n605 0.054
R57716 vdd.n666 vdd.n616 0.054
R57717 vdd.n663 vdd.n625 0.054
R57718 vdd.n660 vdd.n634 0.054
R57719 vdd.n1019 vdd.n1015 0.054
R57720 vdd.n1022 vdd.n1006 0.054
R57721 vdd.n1140 vdd.n1056 0.054
R57722 vdd.n1137 vdd.n1067 0.054
R57723 vdd.n1134 vdd.n1076 0.054
R57724 vdd.n801 vdd.n796 0.054
R57725 vdd.n807 vdd.n803 0.054
R57726 vdd.n835 vdd.n814 0.054
R57727 vdd.n330 vdd.n329 0.054
R57728 vdd.n6015 vdd.n5966 0.054
R57729 vdd.n6245 vdd.n6244 0.054
R57730 vdd.n6128 vdd.n6124 0.054
R57731 vdd.n5751 vdd.n5633 0.054
R57732 vdd.n5748 vdd.n5644 0.054
R57733 vdd.n5745 vdd.n5653 0.054
R57734 vdd.n5742 vdd.n5662 0.054
R57735 vdd.n5494 vdd.n5445 0.054
R57736 vdd.n5491 vdd.n5457 0.054
R57737 vdd.n5488 vdd.n5468 0.054
R57738 vdd.n5255 vdd.n5254 0.054
R57739 vdd.n5242 vdd.n5241 0.054
R57740 vdd.n5228 vdd.n5227 0.054
R57741 vdd.n5216 vdd.n5215 0.054
R57742 vdd.n5581 vdd.n5580 0.054
R57743 vdd.n5586 vdd.n5585 0.054
R57744 vdd.n5592 vdd.n5591 0.054
R57745 vdd.n5598 vdd.n5597 0.054
R57746 vdd.n5360 vdd.n5334 0.054
R57747 vdd.n5363 vdd.n5327 0.054
R57748 vdd.n5366 vdd.n5317 0.054
R57749 vdd.n5369 vdd.n5306 0.054
R57750 vdd.n5116 vdd.n5115 0.054
R57751 vdd.n27643 vdd.n27642 0.054
R57752 vdd.n27640 vdd.n27639 0.054
R57753 vdd.n27624 vdd.n27623 0.054
R57754 vdd.n27518 vdd.n27517 0.054
R57755 vdd.n27470 vdd.n27469 0.054
R57756 vdd.n27376 vdd.n27375 0.054
R57757 vdd.n27365 vdd.n27364 0.054
R57758 vdd.n27362 vdd.n27361 0.054
R57759 vdd.n25600 vdd.n25599 0.054
R57760 vdd.n29479 vdd.n29477 0.054
R57761 vdd.n10094 vdd.n10071 0.054
R57762 vdd.n26425 vdd.n26421 0.054
R57763 vdd.n29 vdd.n28 0.054
R57764 vdd.n4527 vdd.n4526 0.053
R57765 vdd.n24548 vdd.n24543 0.053
R57766 vdd.n10249 vdd.n10132 0.053
R57767 vdd.n34325 vdd.n34314 0.053
R57768 vdd.n34312 vdd.n34302 0.053
R57769 vdd.n34300 vdd.n34290 0.053
R57770 vdd.n34288 vdd.n34279 0.053
R57771 vdd.n34251 vdd.n34250 0.053
R57772 vdd.n34130 vdd.n34126 0.053
R57773 vdd.n34210 vdd.n34198 0.053
R57774 vdd.n34196 vdd.n34184 0.053
R57775 vdd.n34182 vdd.n34171 0.053
R57776 vdd.n33932 vdd.n33928 0.053
R57777 vdd.n33944 vdd.n33943 0.053
R57778 vdd.n33941 vdd.n33940 0.053
R57779 vdd.n33938 vdd.n33937 0.053
R57780 vdd.n33935 vdd.n33934 0.053
R57781 vdd.n34409 vdd.n34408 0.053
R57782 vdd.n34412 vdd.n34411 0.053
R57783 vdd.n34415 vdd.n34414 0.053
R57784 vdd.n34418 vdd.n34417 0.053
R57785 vdd.n34031 vdd.n34028 0.053
R57786 vdd.n34036 vdd.n34033 0.053
R57787 vdd.n34042 vdd.n34038 0.053
R57788 vdd.n34047 vdd.n34044 0.053
R57789 vdd.n34026 vdd.n34025 0.053
R57790 vdd.n35004 vdd.n35003 0.053
R57791 vdd.n35001 vdd.n35000 0.053
R57792 vdd.n34998 vdd.n34997 0.053
R57793 vdd.n34995 vdd.n34994 0.053
R57794 vdd.n34984 vdd.n34983 0.053
R57795 vdd.n34970 vdd.n34969 0.053
R57796 vdd.n34967 vdd.n34966 0.053
R57797 vdd.n34747 vdd.n34746 0.053
R57798 vdd.n34744 vdd.n34743 0.053
R57799 vdd.n34741 vdd.n34740 0.053
R57800 vdd.n34508 vdd.n34497 0.053
R57801 vdd.n34495 vdd.n34483 0.053
R57802 vdd.n34481 vdd.n34471 0.053
R57803 vdd.n34469 vdd.n34462 0.053
R57804 vdd.n34834 vdd.n34831 0.053
R57805 vdd.n34839 vdd.n34836 0.053
R57806 vdd.n34845 vdd.n34841 0.053
R57807 vdd.n34851 vdd.n34847 0.053
R57808 vdd.n34610 vdd.n34594 0.053
R57809 vdd.n34613 vdd.n34612 0.053
R57810 vdd.n34616 vdd.n34615 0.053
R57811 vdd.n34619 vdd.n34618 0.053
R57812 vdd.n34622 vdd.n34621 0.053
R57813 vdd.n749 vdd.n748 0.053
R57814 vdd.n752 vdd.n751 0.053
R57815 vdd.n755 vdd.n754 0.053
R57816 vdd.n758 vdd.n757 0.053
R57817 vdd.n669 vdd.n668 0.053
R57818 vdd.n666 vdd.n665 0.053
R57819 vdd.n663 vdd.n662 0.053
R57820 vdd.n660 vdd.n659 0.053
R57821 vdd.n651 vdd.n650 0.053
R57822 vdd.n1019 vdd.n1018 0.053
R57823 vdd.n1022 vdd.n1021 0.053
R57824 vdd.n1131 vdd.n1085 0.053
R57825 vdd.n1140 vdd.n1139 0.053
R57826 vdd.n1137 vdd.n1136 0.053
R57827 vdd.n1134 vdd.n1133 0.053
R57828 vdd.n1123 vdd.n1122 0.053
R57829 vdd.n1120 vdd.n1119 0.053
R57830 vdd.n801 vdd.n800 0.053
R57831 vdd.n807 vdd.n806 0.053
R57832 vdd.n835 vdd.n834 0.053
R57833 vdd.n5751 vdd.n5750 0.053
R57834 vdd.n5748 vdd.n5747 0.053
R57835 vdd.n5745 vdd.n5744 0.053
R57836 vdd.n5742 vdd.n5741 0.053
R57837 vdd.n5731 vdd.n5730 0.053
R57838 vdd.n5717 vdd.n5716 0.053
R57839 vdd.n5714 vdd.n5713 0.053
R57840 vdd.n5494 vdd.n5493 0.053
R57841 vdd.n5491 vdd.n5490 0.053
R57842 vdd.n5488 vdd.n5487 0.053
R57843 vdd.n5255 vdd.n5244 0.053
R57844 vdd.n5242 vdd.n5230 0.053
R57845 vdd.n5228 vdd.n5218 0.053
R57846 vdd.n5216 vdd.n5209 0.053
R57847 vdd.n5581 vdd.n5578 0.053
R57848 vdd.n5586 vdd.n5583 0.053
R57849 vdd.n5592 vdd.n5588 0.053
R57850 vdd.n5598 vdd.n5594 0.053
R57851 vdd.n5357 vdd.n5341 0.053
R57852 vdd.n5360 vdd.n5359 0.053
R57853 vdd.n5363 vdd.n5362 0.053
R57854 vdd.n5366 vdd.n5365 0.053
R57855 vdd.n5369 vdd.n5368 0.053
R57856 vdd.n27633 vdd.n27632 0.053
R57857 vdd.n27512 vdd.n27511 0.053
R57858 vdd.n26007 vdd.n26006 0.053
R57859 vdd.n25994 vdd.n25993 0.053
R57860 vdd.n25983 vdd.n25982 0.053
R57861 vdd.n25972 vdd.n25971 0.053
R57862 vdd.n25963 vdd.n25962 0.053
R57863 vdd.n25902 vdd.n25901 0.053
R57864 vdd.n25891 vdd.n25890 0.053
R57865 vdd.n25882 vdd.n25881 0.053
R57866 vdd.n25873 vdd.n25872 0.053
R57867 vdd.n25866 vdd.n25865 0.053
R57868 vdd.n25797 vdd.n25796 0.053
R57869 vdd.n25785 vdd.n25784 0.053
R57870 vdd.n25774 vdd.n25773 0.053
R57871 vdd.n25765 vdd.n25764 0.053
R57872 vdd.n4016 vdd.n2679 0.053
R57873 vdd.n10094 vdd.n10089 0.053
R57874 vdd.n10221 vdd.n10220 0.053
R57875 vdd.n10221 vdd.n10128 0.053
R57876 vdd.n11886 vdd.n11880 0.053
R57877 vdd.n16788 vdd.n16787 0.053
R57878 vdd.n16789 vdd.n16788 0.053
R57879 vdd.n21977 vdd.n21971 0.053
R57880 vdd.n33391 vdd.n33376 0.053
R57881 vdd.n705 vdd.n690 0.053
R57882 vdd.n294 vdd.n291 0.053
R57883 vdd.n4868 vdd.n4865 0.053
R57884 vdd.n4312 vdd.n4311 0.052
R57885 vdd.n33805 vdd.n33804 0.052
R57886 vdd.n33932 vdd.n33931 0.052
R57887 vdd.n34026 vdd.n34023 0.052
R57888 vdd.n34825 vdd.n34824 0.052
R57889 vdd.n34610 vdd.n34609 0.052
R57890 vdd.n1131 vdd.n1130 0.052
R57891 vdd.n544 vdd.n541 0.052
R57892 vdd.n549 vdd.n546 0.052
R57893 vdd.n555 vdd.n551 0.052
R57894 vdd.n560 vdd.n557 0.052
R57895 vdd.n453 vdd.n442 0.052
R57896 vdd.n440 vdd.n432 0.052
R57897 vdd.n430 vdd.n420 0.052
R57898 vdd.n418 vdd.n409 0.052
R57899 vdd.n391 vdd.n390 0.052
R57900 vdd.n60 vdd.n56 0.052
R57901 vdd.n66 vdd.n62 0.052
R57902 vdd.n173 vdd.n162 0.052
R57903 vdd.n160 vdd.n150 0.052
R57904 vdd.n148 vdd.n138 0.052
R57905 vdd.n136 vdd.n127 0.052
R57906 vdd.n106 vdd.n105 0.052
R57907 vdd.n94 vdd.n93 0.052
R57908 vdd.n275 vdd.n272 0.052
R57909 vdd.n368 vdd.n356 0.052
R57910 vdd.n354 vdd.n344 0.052
R57911 vdd.n342 vdd.n332 0.052
R57912 vdd.n5572 vdd.n5571 0.052
R57913 vdd.n5357 vdd.n5356 0.052
R57914 vdd.n5164 vdd.n5153 0.052
R57915 vdd.n5151 vdd.n5139 0.052
R57916 vdd.n5137 vdd.n5128 0.052
R57917 vdd.n5126 vdd.n5118 0.052
R57918 vdd.n5089 vdd.n5088 0.052
R57919 vdd.n5075 vdd.n5074 0.052
R57920 vdd.n4848 vdd.n4845 0.052
R57921 vdd.n4768 vdd.n4757 0.052
R57922 vdd.n4755 vdd.n4744 0.052
R57923 vdd.n4742 vdd.n4735 0.052
R57924 vdd.n4733 vdd.n4728 0.052
R57925 vdd.n5017 vdd.n5014 0.052
R57926 vdd.n5022 vdd.n5019 0.052
R57927 vdd.n5028 vdd.n5024 0.052
R57928 vdd.n5034 vdd.n5030 0.052
R57929 vdd.n4675 vdd.n4672 0.052
R57930 vdd.n4680 vdd.n4677 0.052
R57931 vdd.n4686 vdd.n4682 0.052
R57932 vdd.n4691 vdd.n4688 0.052
R57933 vdd.n4925 vdd.n4924 0.052
R57934 vdd.n4922 vdd.n4921 0.052
R57935 vdd.n4919 vdd.n4910 0.052
R57936 vdd.n4569 vdd.n4497 0.052
R57937 vdd.n25646 vdd.n25645 0.052
R57938 vdd.n4018 vdd.n4017 0.052
R57939 vdd.n11728 vdd.n11723 0.052
R57940 vdd.n21804 vdd.n21802 0.052
R57941 vdd.n24940 vdd.n24939 0.052
R57942 ldomc_0.vdd vdd.n6363 0.052
R57943 vdd.n35314 vdd.n35313 0.051
R57944 vdd.n5870 vdd.n5865 0.051
R57945 vdd.n4855 vdd.n4854 0.051
R57946 vdd.n22341 vdd.n22340 0.051
R57947 vdd.n24304 vdd.n24303 0.051
R57948 vdd.n278 vdd.n277 0.051
R57949 vdd.n33424 vdd.n33421 0.051
R57950 vdd.n33429 vdd.n33426 0.051
R57951 vdd.n33435 vdd.n33431 0.051
R57952 vdd.n33440 vdd.n33437 0.051
R57953 vdd.n33511 vdd.n33508 0.051
R57954 vdd.n33313 vdd.n33310 0.051
R57955 vdd.n33350 vdd.n33339 0.051
R57956 vdd.n33337 vdd.n33327 0.051
R57957 vdd.n33325 vdd.n33315 0.051
R57958 vdd.n33313 vdd.n33305 0.051
R57959 vdd.n33537 vdd.n33535 0.051
R57960 vdd.n33543 vdd.n33539 0.051
R57961 vdd.n33549 vdd.n33545 0.051
R57962 vdd.n33649 vdd.n33646 0.051
R57963 vdd.n33674 vdd.n33663 0.051
R57964 vdd.n33661 vdd.n33651 0.051
R57965 vdd.n33649 vdd.n33639 0.051
R57966 vdd.n33607 vdd.n33606 0.051
R57967 vdd.n33595 vdd.n33594 0.051
R57968 vdd.n33587 vdd.n33586 0.051
R57969 vdd.n33829 vdd.n33826 0.051
R57970 vdd.n33841 vdd.n33831 0.051
R57971 vdd.n33829 vdd.n33819 0.051
R57972 vdd.n33817 vdd.n33807 0.051
R57973 vdd.n34108 vdd.n34107 0.051
R57974 vdd.n34288 vdd.n34285 0.051
R57975 vdd.n33932 vdd.n33929 0.051
R57976 vdd.n33953 vdd.n33952 0.051
R57977 vdd.n35554 vdd.n35551 0.051
R57978 vdd.n35039 vdd.n35038 0.051
R57979 vdd.n34995 vdd.n34921 0.051
R57980 vdd.n34455 vdd.n34454 0.051
R57981 vdd.n1035 vdd.n1032 0.051
R57982 vdd.n660 vdd.n639 0.051
R57983 vdd.n1134 vdd.n1083 0.051
R57984 vdd.n943 vdd.n942 0.051
R57985 vdd.n544 vdd.n537 0.051
R57986 vdd.n26 vdd.n25 0.051
R57987 vdd.n407 vdd.n406 0.051
R57988 vdd.n6018 vdd.n5964 0.051
R57989 vdd.n5816 vdd.n5815 0.051
R57990 vdd.n6237 vdd.n6236 0.051
R57991 vdd.n6216 vdd.n6202 0.051
R57992 vdd.n5742 vdd.n5668 0.051
R57993 vdd.n5202 vdd.n5201 0.051
R57994 vdd.n4675 vdd.n4648 0.051
R57995 vdd.n5012 vdd.n5003 0.051
R57996 vdd.n5043 vdd.n5042 0.051
R57997 vdd.n4670 vdd.n4669 0.051
R57998 vdd.n4572 vdd.n4495 0.051
R57999 vdd.n4581 vdd.n4580 0.051
R58000 vdd.n4578 vdd.n4577 0.051
R58001 vdd.n4575 vdd.n4574 0.051
R58002 vdd.n4572 vdd.n4571 0.051
R58003 vdd.n4561 vdd.n4560 0.051
R58004 vdd.n4547 vdd.n4546 0.051
R58005 vdd.n4544 vdd.n4543 0.051
R58006 vdd.n4321 vdd.n4320 0.051
R58007 vdd.n4318 vdd.n4317 0.051
R58008 vdd.n4315 vdd.n4314 0.051
R58009 vdd.n4032 vdd.n4031 0.051
R58010 vdd.n4085 vdd.n4074 0.051
R58011 vdd.n4072 vdd.n4060 0.051
R58012 vdd.n4058 vdd.n4048 0.051
R58013 vdd.n4046 vdd.n4039 0.051
R58014 vdd.n4407 vdd.n4404 0.051
R58015 vdd.n4413 vdd.n4409 0.051
R58016 vdd.n4419 vdd.n4415 0.051
R58017 vdd.n4425 vdd.n4421 0.051
R58018 vdd.n4191 vdd.n4190 0.051
R58019 vdd.n4194 vdd.n4193 0.051
R58020 vdd.n4197 vdd.n4196 0.051
R58021 vdd.n4200 vdd.n4199 0.051
R58022 vdd.n27564 vdd.n27563 0.051
R58023 vdd.n27582 vdd.n27581 0.051
R58024 vdd.n27505 vdd.n27504 0.051
R58025 vdd.n27488 vdd.n27487 0.051
R58026 vdd.n27404 vdd.n27403 0.051
R58027 vdd.n27322 vdd.n27320 0.051
R58028 vdd.n25700 vdd.n25699 0.051
R58029 vdd.n25819 vdd.n25734 0.051
R58030 vdd.n25774 vdd.n25772 0.051
R58031 vdd.n30807 vdd.n30806 0.051
R58032 vdd.n11774 vdd.n11773 0.051
R58033 vdd.n11874 vdd.n11873 0.051
R58034 vdd.n21863 vdd.n21862 0.051
R58035 vdd.n21965 vdd.n21964 0.051
R58036 vdd.n35489 vdd.n35488 0.051
R58037 vdd.n5819 vdd.n5818 0.051
R58038 vdd.n354 vdd.n321 0.051
R58039 vdd.n24976 vdd.n24974 0.05
R58040 vdd.n34136 vdd.n34135 0.05
R58041 vdd.n34953 vdd.n34952 0.05
R58042 vdd.n5700 vdd.n5699 0.05
R58043 vdd.n34267 vdd.n34266 0.05
R58044 vdd.n34139 vdd.n34138 0.05
R58045 vdd.n34145 vdd.n34144 0.05
R58046 vdd.n34151 vdd.n34150 0.05
R58047 vdd.n34277 vdd.n34276 0.05
R58048 vdd.n33963 vdd.n33962 0.05
R58049 vdd.n34437 vdd.n34436 0.05
R58050 vdd.n34022 vdd.n34021 0.05
R58051 vdd.n35591 vdd.n35580 0.05
R58052 vdd.n35578 vdd.n35568 0.05
R58053 vdd.n35566 vdd.n35556 0.05
R58054 vdd.n35554 vdd.n35545 0.05
R58055 vdd.n35517 vdd.n35516 0.05
R58056 vdd.n35503 vdd.n35502 0.05
R58057 vdd.n35492 vdd.n35491 0.05
R58058 vdd.n35095 vdd.n35084 0.05
R58059 vdd.n35082 vdd.n35070 0.05
R58060 vdd.n35068 vdd.n35058 0.05
R58061 vdd.n35056 vdd.n35049 0.05
R58062 vdd.n35430 vdd.n35427 0.05
R58063 vdd.n35436 vdd.n35432 0.05
R58064 vdd.n35442 vdd.n35438 0.05
R58065 vdd.n35448 vdd.n35444 0.05
R58066 vdd.n35193 vdd.n35190 0.05
R58067 vdd.n35198 vdd.n35195 0.05
R58068 vdd.n35204 vdd.n35200 0.05
R58069 vdd.n35210 vdd.n35206 0.05
R58070 vdd.n35331 vdd.n35330 0.05
R58071 vdd.n35328 vdd.n35327 0.05
R58072 vdd.n35325 vdd.n35316 0.05
R58073 vdd.n34992 vdd.n34923 0.05
R58074 vdd.n34990 vdd.n34989 0.05
R58075 vdd.n34683 vdd.n34682 0.05
R58076 vdd.n34686 vdd.n34685 0.05
R58077 vdd.n34689 vdd.n34688 0.05
R58078 vdd.n34528 vdd.n34527 0.05
R58079 vdd.n34870 vdd.n34869 0.05
R58080 vdd.n34608 vdd.n34607 0.05
R58081 vdd.n1041 vdd.n1040 0.05
R58082 vdd.n1044 vdd.n1043 0.05
R58083 vdd.n1129 vdd.n1128 0.05
R58084 vdd.n1126 vdd.n1125 0.05
R58085 vdd.n943 vdd.n930 0.05
R58086 vdd.n897 vdd.n896 0.05
R58087 vdd.n832 vdd.n824 0.05
R58088 vdd.n330 vdd.n325 0.05
R58089 vdd.n6027 vdd.n6026 0.05
R58090 vdd.n6024 vdd.n6023 0.05
R58091 vdd.n6021 vdd.n6020 0.05
R58092 vdd.n6018 vdd.n6017 0.05
R58093 vdd.n6007 vdd.n6006 0.05
R58094 vdd.n6004 vdd.n6003 0.05
R58095 vdd.n6228 vdd.n6227 0.05
R58096 vdd.n6225 vdd.n6224 0.05
R58097 vdd.n6222 vdd.n6221 0.05
R58098 vdd.n6219 vdd.n6218 0.05
R58099 vdd.n6116 vdd.n6115 0.05
R58100 vdd.n6119 vdd.n6118 0.05
R58101 vdd.n6122 vdd.n6121 0.05
R58102 vdd.n6324 vdd.n6323 0.05
R58103 vdd.n6327 vdd.n6326 0.05
R58104 vdd.n6330 vdd.n6329 0.05
R58105 vdd.n6333 vdd.n6332 0.05
R58106 vdd.n5911 vdd.n5899 0.05
R58107 vdd.n5897 vdd.n5885 0.05
R58108 vdd.n5883 vdd.n5872 0.05
R58109 vdd.n5739 vdd.n5670 0.05
R58110 vdd.n5737 vdd.n5736 0.05
R58111 vdd.n5430 vdd.n5429 0.05
R58112 vdd.n5433 vdd.n5432 0.05
R58113 vdd.n5436 vdd.n5435 0.05
R58114 vdd.n5275 vdd.n5274 0.05
R58115 vdd.n5617 vdd.n5616 0.05
R58116 vdd.n5355 vdd.n5354 0.05
R58117 vdd.n5116 vdd.n5107 0.05
R58118 vdd.n5012 vdd.n5011 0.05
R58119 vdd.n31288 vdd.n31286 0.05
R58120 vdd.n32087 vdd.n32085 0.05
R58121 vdd.n32359 vdd.n32358 0.05
R58122 vdd.n27613 vdd.n27612 0.05
R58123 vdd.n27494 vdd.n27493 0.05
R58124 vdd.n27412 vdd.n27411 0.05
R58125 vdd.n27393 vdd.n27392 0.05
R58126 vdd.n26064 vdd.n26063 0.05
R58127 vdd.n26061 vdd.n26060 0.05
R58128 vdd.n26054 vdd.n26053 0.05
R58129 vdd.n26045 vdd.n26044 0.05
R58130 vdd.n25955 vdd.n25954 0.05
R58131 vdd.n25949 vdd.n25948 0.05
R58132 vdd.n25916 vdd.n25915 0.05
R58133 vdd.n25819 vdd.n25818 0.05
R58134 vdd.n25817 vdd.n25816 0.05
R58135 vdd.n25814 vdd.n25813 0.05
R58136 vdd.n25600 vdd.n25588 0.05
R58137 vdd.n25475 vdd.n25474 0.05
R58138 vdd.n10094 vdd.n10085 0.05
R58139 vdd.n11904 vdd.n11903 0.05
R58140 vdd.n11893 vdd.n11892 0.05
R58141 vdd.n21995 vdd.n21994 0.05
R58142 vdd.n21984 vdd.n21983 0.05
R58143 vdd.n33661 vdd.n33578 0.05
R58144 vdd.n1137 vdd.n1065 0.05
R58145 vdd.n32076 vdd.n32075 0.049
R58146 vdd.n31782 vdd.n31781 0.049
R58147 vdd.n4526 vdd.n4525 0.049
R58148 vdd.n31475 vdd.n31469 0.049
R58149 vdd.n31475 vdd.n31471 0.049
R58150 vdd.n31631 vdd.n31620 0.049
R58151 vdd.n31631 vdd.n31621 0.049
R58152 vdd.n26619 vdd.n26614 0.049
R58153 vdd.n26619 vdd.n26615 0.049
R58154 vdd.n34132 vdd.n34131 0.049
R58155 vdd.n34965 vdd.n34964 0.049
R58156 vdd.n5712 vdd.n5711 0.049
R58157 vdd.n34261 vdd.n34258 0.049
R58158 vdd.n35527 vdd.n35524 0.049
R58159 vdd.n34986 vdd.n34939 0.049
R58160 vdd.n6009 vdd.n5982 0.049
R58161 vdd.n5733 vdd.n5686 0.049
R58162 vdd.n4563 vdd.n4513 0.049
R58163 vdd.n33303 vdd.n33302 0.049
R58164 vdd.n33637 vdd.n33628 0.049
R58165 vdd.n34277 vdd.n34268 0.049
R58166 vdd.n34992 vdd.n34991 0.049
R58167 vdd.n658 vdd.n657 0.049
R58168 vdd.n832 vdd.n831 0.049
R58169 vdd.n76 vdd.n75 0.049
R58170 vdd.n82 vdd.n81 0.049
R58171 vdd.n115 vdd.n114 0.049
R58172 vdd.n283 vdd.n282 0.049
R58173 vdd.n289 vdd.n288 0.049
R58174 vdd.n295 vdd.n294 0.049
R58175 vdd.n299 vdd.n298 0.049
R58176 vdd.n5739 vdd.n5738 0.049
R58177 vdd.n5106 vdd.n5105 0.049
R58178 vdd.n4857 vdd.n4856 0.049
R58179 vdd.n4863 vdd.n4862 0.049
R58180 vdd.n4869 vdd.n4868 0.049
R58181 vdd.n4788 vdd.n4787 0.049
R58182 vdd.n5055 vdd.n5054 0.049
R58183 vdd.n4666 vdd.n4665 0.049
R58184 vdd.n4398 vdd.n4397 0.049
R58185 vdd.n4188 vdd.n4187 0.049
R58186 vdd.n10201 vdd.n10200 0.049
R58187 vdd.n10223 vdd.n10133 0.049
R58188 vdd.n11749 vdd.n11721 0.049
R58189 vdd.n16694 vdd.n16693 0.049
R58190 vdd.n16679 vdd.n16678 0.049
R58191 vdd.n21824 vdd.n21823 0.049
R58192 vdd.n812 vdd.n811 0.049
R58193 vdd.n212 vdd.n211 0.049
R58194 vdd.n33763 vdd.n33760 0.049
R58195 vdd.n34150 vdd.n34147 0.049
R58196 vdd.n35272 vdd.n35269 0.049
R58197 vdd.n34688 vdd.n34667 0.049
R58198 vdd.n900 vdd.n899 0.049
R58199 vdd.n5836 vdd.n5795 0.049
R58200 vdd.n5435 vdd.n5414 0.049
R58201 vdd.n4262 vdd.n4244 0.049
R58202 vdd.n945 vdd.n944 0.048
R58203 vdd.n24902 vdd.n24899 0.048
R58204 vdd.n4854 vdd.n4853 0.048
R58205 vdd.n4851 vdd.n4850 0.048
R58206 vdd.n33559 vdd.n33558 0.048
R58207 vdd.n33565 vdd.n33564 0.048
R58208 vdd.n33627 vdd.n33626 0.048
R58209 vdd.n33616 vdd.n33615 0.048
R58210 vdd.n33752 vdd.n33751 0.048
R58211 vdd.n33758 vdd.n33757 0.048
R58212 vdd.n33764 vdd.n33763 0.048
R58213 vdd.n33769 vdd.n33768 0.048
R58214 vdd.n35421 vdd.n35420 0.048
R58215 vdd.n35188 vdd.n35185 0.048
R58216 vdd.n125 vdd.n124 0.048
R58217 vdd.n6216 vdd.n6215 0.048
R58218 vdd.n6321 vdd.n6320 0.048
R58219 vdd.n4567 vdd.n4566 0.048
R58220 vdd.n4260 vdd.n4259 0.048
R58221 vdd.n4263 vdd.n4262 0.048
R58222 vdd.n4105 vdd.n4104 0.048
R58223 vdd.n4444 vdd.n4443 0.048
R58224 vdd.n4186 vdd.n4185 0.048
R58225 vdd.n27376 vdd.n27366 0.048
R58226 vdd.n25998 vdd.n25683 0.048
R58227 vdd.n25917 vdd.n25916 0.048
R58228 vdd.n25818 vdd.n25817 0.048
R58229 vdd.n24547 vdd.n24546 0.048
R58230 vdd.n24970 vdd.n24958 0.048
R58231 vdd.n105 vdd.n102 0.047
R58232 vdd.n34137 vdd.n34136 0.047
R58233 vdd.n34952 vdd.n34951 0.047
R58234 vdd.n5699 vdd.n5698 0.047
R58235 vdd.n928 vdd.n927 0.047
R58236 vdd.n33748 vdd.n33747 0.047
R58237 vdd.n31314 vdd.n31313 0.047
R58238 vdd.n33440 vdd.n33400 0.047
R58239 vdd.n33419 vdd.n33418 0.047
R58240 vdd.n33564 vdd.n33492 0.047
R58241 vdd.n33549 vdd.n33523 0.047
R58242 vdd.n33350 vdd.n33347 0.047
R58243 vdd.n33586 vdd.n33582 0.047
R58244 vdd.n34130 vdd.n34116 0.047
R58245 vdd.n34124 vdd.n34122 0.047
R58246 vdd.n34325 vdd.n34322 0.047
R58247 vdd.n34418 vdd.n34376 0.047
R58248 vdd.n34415 vdd.n34388 0.047
R58249 vdd.n33941 vdd.n33910 0.047
R58250 vdd.n33944 vdd.n33898 0.047
R58251 vdd.n33965 vdd.n33872 0.047
R58252 vdd.n34047 vdd.n33982 0.047
R58253 vdd.n34042 vdd.n33991 0.047
R58254 vdd.n34026 vdd.n34008 0.047
R58255 vdd.n35188 vdd.n35170 0.047
R58256 vdd.n35204 vdd.n35153 0.047
R58257 vdd.n35591 vdd.n35588 0.047
R58258 vdd.n35491 vdd.n35472 0.047
R58259 vdd.n35533 vdd.n35532 0.047
R58260 vdd.n35267 vdd.n35266 0.047
R58261 vdd.n35273 vdd.n35272 0.047
R58262 vdd.n35126 vdd.n35123 0.047
R58263 vdd.n35095 vdd.n35092 0.047
R58264 vdd.n35082 vdd.n35079 0.047
R58265 vdd.n35442 vdd.n35407 0.047
R58266 vdd.n35448 vdd.n35399 0.047
R58267 vdd.n35115 vdd.n35114 0.047
R58268 vdd.n35459 vdd.n35458 0.047
R58269 vdd.n35210 vdd.n35144 0.047
R58270 vdd.n35184 vdd.n35183 0.047
R58271 vdd.n35183 vdd.n35182 0.047
R58272 vdd.n34966 vdd.n34950 0.047
R58273 vdd.n35004 vdd.n34894 0.047
R58274 vdd.n34851 vdd.n34802 0.047
R58275 vdd.n34845 vdd.n34811 0.047
R58276 vdd.n34495 vdd.n34492 0.047
R58277 vdd.n34508 vdd.n34505 0.047
R58278 vdd.n34539 vdd.n34536 0.047
R58279 vdd.n34622 vdd.n34557 0.047
R58280 vdd.n34619 vdd.n34568 0.047
R58281 vdd.n34610 vdd.n34592 0.047
R58282 vdd.n758 vdd.n719 0.047
R58283 vdd.n1043 vdd.n979 0.047
R58284 vdd.n1022 vdd.n1004 0.047
R58285 vdd.n669 vdd.n613 0.047
R58286 vdd.n657 vdd.n640 0.047
R58287 vdd.n947 vdd.n925 0.047
R58288 vdd.n560 vdd.n518 0.047
R58289 vdd.n540 vdd.n539 0.047
R58290 vdd.n66 vdd.n47 0.047
R58291 vdd.n407 vdd.n405 0.047
R58292 vdd.n453 vdd.n450 0.047
R58293 vdd.n407 vdd.n404 0.047
R58294 vdd.n294 vdd.n245 0.047
R58295 vdd.n275 vdd.n271 0.047
R58296 vdd.n136 vdd.n133 0.047
R58297 vdd.n173 vdd.n170 0.047
R58298 vdd.n126 vdd.n125 0.047
R58299 vdd.n342 vdd.n339 0.047
R58300 vdd.n6321 vdd.n6303 0.047
R58301 vdd.n6330 vdd.n6279 0.047
R58302 vdd.n6027 vdd.n5937 0.047
R58303 vdd.n5826 vdd.n5824 0.047
R58304 vdd.n6013 vdd.n6012 0.047
R58305 vdd.n5831 vdd.n5830 0.047
R58306 vdd.n5834 vdd.n5833 0.047
R58307 vdd.n5837 vdd.n5836 0.047
R58308 vdd.n6250 vdd.n6146 0.047
R58309 vdd.n6228 vdd.n6172 0.047
R58310 vdd.n6225 vdd.n6184 0.047
R58311 vdd.n6119 vdd.n6101 0.047
R58312 vdd.n6122 vdd.n6090 0.047
R58313 vdd.n6248 vdd.n6247 0.047
R58314 vdd.n6132 vdd.n6131 0.047
R58315 vdd.n6333 vdd.n6267 0.047
R58316 vdd.n6318 vdd.n6307 0.047
R58317 vdd.n6319 vdd.n6318 0.047
R58318 vdd.n5713 vdd.n5697 0.047
R58319 vdd.n5751 vdd.n5641 0.047
R58320 vdd.n5598 vdd.n5549 0.047
R58321 vdd.n5592 vdd.n5558 0.047
R58322 vdd.n5242 vdd.n5239 0.047
R58323 vdd.n5255 vdd.n5252 0.047
R58324 vdd.n5286 vdd.n5283 0.047
R58325 vdd.n5369 vdd.n5304 0.047
R58326 vdd.n5366 vdd.n5315 0.047
R58327 vdd.n5357 vdd.n5339 0.047
R58328 vdd.n4912 vdd.n4911 0.047
R58329 vdd.n5164 vdd.n5161 0.047
R58330 vdd.n5151 vdd.n5148 0.047
R58331 vdd.n5116 vdd.n5113 0.047
R58332 vdd.n4848 vdd.n4843 0.047
R58333 vdd.n4768 vdd.n4765 0.047
R58334 vdd.n4755 vdd.n4752 0.047
R58335 vdd.n5028 vdd.n4989 0.047
R58336 vdd.n5034 vdd.n4980 0.047
R58337 vdd.n5059 vdd.n4958 0.047
R58338 vdd.n4691 vdd.n4628 0.047
R58339 vdd.n4670 vdd.n4667 0.047
R58340 vdd.n4925 vdd.n4888 0.047
R58341 vdd.n4543 vdd.n4524 0.047
R58342 vdd.n4581 vdd.n4468 0.047
R58343 vdd.n4425 vdd.n4376 0.047
R58344 vdd.n4419 vdd.n4384 0.047
R58345 vdd.n4072 vdd.n4069 0.047
R58346 vdd.n4085 vdd.n4082 0.047
R58347 vdd.n4116 vdd.n4113 0.047
R58348 vdd.n4200 vdd.n4134 0.047
R58349 vdd.n4197 vdd.n4146 0.047
R58350 vdd.n4188 vdd.n4170 0.047
R58351 vdd.n27607 vdd.n27260 0.047
R58352 vdd.n27488 vdd.n27270 0.047
R58353 vdd.n27546 vdd.n27544 0.047
R58354 vdd.n27557 vdd.n27555 0.047
R58355 vdd.n27387 vdd.n27290 0.047
R58356 vdd.n27456 vdd.n27454 0.047
R58357 vdd.n26034 vdd.n26033 0.047
R58358 vdd.n25983 vdd.n25981 0.047
R58359 vdd.n25994 vdd.n25992 0.047
R58360 vdd.n25998 vdd.n25997 0.047
R58361 vdd.n25942 vdd.n25941 0.047
R58362 vdd.n25931 vdd.n25930 0.047
R58363 vdd.n25920 vdd.n25919 0.047
R58364 vdd.n25902 vdd.n25900 0.047
R58365 vdd.n25858 vdd.n25857 0.047
R58366 vdd.n25850 vdd.n25849 0.047
R58367 vdd.n25839 vdd.n25838 0.047
R58368 vdd.n25507 vdd.n25505 0.047
R58369 vdd.n25646 vdd.n25414 0.047
R58370 vdd.n25581 vdd.n25579 0.047
R58371 vdd.n25518 vdd.n25441 0.047
R58372 vdd.n30163 vdd.n30161 0.047
R58373 vdd.n27668 vdd.n27667 0.047
R58374 vdd.n10217 vdd.n10073 0.047
R58375 vdd.n10222 vdd.n10074 0.047
R58376 vdd.n13876 vdd.n13875 0.047
R58377 vdd.n13885 vdd.n13883 0.047
R58378 vdd.n13923 vdd.n8651 0.047
R58379 vdd.n13921 vdd.n8652 0.047
R58380 vdd.n13940 vdd.n13939 0.047
R58381 vdd.n13957 vdd.n13947 0.047
R58382 vdd.n13955 vdd.n13949 0.047
R58383 vdd.n13999 vdd.n13998 0.047
R58384 vdd.n14017 vdd.n14015 0.047
R58385 vdd.n14027 vdd.n8580 0.047
R58386 vdd.n14035 vdd.n14034 0.047
R58387 vdd.n14085 vdd.n8546 0.047
R58388 vdd.n14083 vdd.n8547 0.047
R58389 vdd.n14101 vdd.n14100 0.047
R58390 vdd.n14165 vdd.n14164 0.047
R58391 vdd.n14174 vdd.n14172 0.047
R58392 vdd.n14213 vdd.n8431 0.047
R58393 vdd.n14211 vdd.n8432 0.047
R58394 vdd.n14230 vdd.n14229 0.047
R58395 vdd.n14247 vdd.n14237 0.047
R58396 vdd.n14245 vdd.n14239 0.047
R58397 vdd.n14290 vdd.n14289 0.047
R58398 vdd.n14306 vdd.n14305 0.047
R58399 vdd.n14315 vdd.n14313 0.047
R58400 vdd.n14367 vdd.n8323 0.047
R58401 vdd.n14365 vdd.n8324 0.047
R58402 vdd.n14386 vdd.n8309 0.047
R58403 vdd.n14391 vdd.n14390 0.047
R58404 vdd.n14448 vdd.n14444 0.047
R58405 vdd.n14446 vdd.n8229 0.047
R58406 vdd.n14475 vdd.n14474 0.047
R58407 vdd.n14477 vdd.n8195 0.047
R58408 vdd.n14555 vdd.n14536 0.047
R58409 vdd.n14553 vdd.n14537 0.047
R58410 vdd.n14606 vdd.n8178 0.047
R58411 vdd.n13157 vdd.n13156 0.047
R58412 vdd.n13166 vdd.n13165 0.047
R58413 vdd.n13173 vdd.n13171 0.047
R58414 vdd.n13224 vdd.n9196 0.047
R58415 vdd.n13222 vdd.n9198 0.047
R58416 vdd.n13282 vdd.n9138 0.047
R58417 vdd.n13312 vdd.n13309 0.047
R58418 vdd.n13310 vdd.n9110 0.047
R58419 vdd.n9118 vdd.n9115 0.047
R58420 vdd.n9116 vdd.n9076 0.047
R58421 vdd.n9084 vdd.n9082 0.047
R58422 vdd.n13383 vdd.n9059 0.047
R58423 vdd.n13433 vdd.n9026 0.047
R58424 vdd.n13431 vdd.n9027 0.047
R58425 vdd.n13451 vdd.n13449 0.047
R58426 vdd.n13461 vdd.n9008 0.047
R58427 vdd.n13469 vdd.n13468 0.047
R58428 vdd.n13516 vdd.n8974 0.047
R58429 vdd.n13514 vdd.n8976 0.047
R58430 vdd.n13574 vdd.n8916 0.047
R58431 vdd.n13604 vdd.n13601 0.047
R58432 vdd.n13602 vdd.n8889 0.047
R58433 vdd.n8897 vdd.n8894 0.047
R58434 vdd.n8895 vdd.n8856 0.047
R58435 vdd.n8864 vdd.n8862 0.047
R58436 vdd.n13675 vdd.n8839 0.047
R58437 vdd.n13725 vdd.n8806 0.047
R58438 vdd.n13723 vdd.n8807 0.047
R58439 vdd.n10216 vdd.n10215 0.047
R58440 vdd.n10461 vdd.n10286 0.047
R58441 vdd.n10459 vdd.n10287 0.047
R58442 vdd.n10436 vdd.n10303 0.047
R58443 vdd.n10434 vdd.n10304 0.047
R58444 vdd.n10423 vdd.n10422 0.047
R58445 vdd.n10411 vdd.n10313 0.047
R58446 vdd.n10409 vdd.n10323 0.047
R58447 vdd.n10400 vdd.n10399 0.047
R58448 vdd.n10348 vdd.n10335 0.047
R58449 vdd.n10374 vdd.n10373 0.047
R58450 vdd.n10364 vdd.n10361 0.047
R58451 vdd.n10362 vdd.n9295 0.047
R58452 vdd.n13067 vdd.n9304 0.047
R58453 vdd.n13065 vdd.n9305 0.047
R58454 vdd.n13054 vdd.n13053 0.047
R58455 vdd.n9339 vdd.n9338 0.047
R58456 vdd.n13036 vdd.n9351 0.047
R58457 vdd.n9379 vdd.n9377 0.047
R58458 vdd.n9391 vdd.n9365 0.047
R58459 vdd.n13020 vdd.n13019 0.047
R58460 vdd.n13008 vdd.n9396 0.047
R58461 vdd.n13006 vdd.n9404 0.047
R58462 vdd.n9446 vdd.n9426 0.047
R58463 vdd.n12980 vdd.n9450 0.047
R58464 vdd.n12978 vdd.n9451 0.047
R58465 vdd.n12967 vdd.n12966 0.047
R58466 vdd.n9493 vdd.n9489 0.047
R58467 vdd.n9491 vdd.n9480 0.047
R58468 vdd.n9506 vdd.n9505 0.047
R58469 vdd.n12942 vdd.n9514 0.047
R58470 vdd.n9546 vdd.n9530 0.047
R58471 vdd.n12925 vdd.n12924 0.047
R58472 vdd.n12913 vdd.n9551 0.047
R58473 vdd.n12911 vdd.n9559 0.047
R58474 vdd.n9589 vdd.n9587 0.047
R58475 vdd.n9601 vdd.n9576 0.047
R58476 vdd.n12895 vdd.n12894 0.047
R58477 vdd.n9643 vdd.n9639 0.047
R58478 vdd.n9641 vdd.n9627 0.047
R58479 vdd.n9656 vdd.n9655 0.047
R58480 vdd.n12859 vdd.n9664 0.047
R58481 vdd.n12857 vdd.n9665 0.047
R58482 vdd.n12846 vdd.n12845 0.047
R58483 vdd.n9699 vdd.n9698 0.047
R58484 vdd.n12828 vdd.n9711 0.047
R58485 vdd.n9739 vdd.n9737 0.047
R58486 vdd.n9751 vdd.n9725 0.047
R58487 vdd.n12812 vdd.n12811 0.047
R58488 vdd.n12800 vdd.n9756 0.047
R58489 vdd.n12798 vdd.n9764 0.047
R58490 vdd.n9805 vdd.n9786 0.047
R58491 vdd.n12772 vdd.n9809 0.047
R58492 vdd.n12770 vdd.n9810 0.047
R58493 vdd.n12759 vdd.n12758 0.047
R58494 vdd.n9853 vdd.n9849 0.047
R58495 vdd.n9851 vdd.n9840 0.047
R58496 vdd.n9866 vdd.n9865 0.047
R58497 vdd.n12734 vdd.n9874 0.047
R58498 vdd.n9906 vdd.n9891 0.047
R58499 vdd.n12717 vdd.n12716 0.047
R58500 vdd.n12705 vdd.n9911 0.047
R58501 vdd.n12703 vdd.n9918 0.047
R58502 vdd.n9949 vdd.n9947 0.047
R58503 vdd.n9961 vdd.n9935 0.047
R58504 vdd.n12687 vdd.n12686 0.047
R58505 vdd.n10003 vdd.n9999 0.047
R58506 vdd.n10001 vdd.n9987 0.047
R58507 vdd.n10016 vdd.n10015 0.047
R58508 vdd.n12651 vdd.n10024 0.047
R58509 vdd.n12649 vdd.n10025 0.047
R58510 vdd.n12638 vdd.n12637 0.047
R58511 vdd.n10160 vdd.n10149 0.047
R58512 vdd.n24204 vdd.n24203 0.047
R58513 vdd.n16589 vdd.n16588 0.047
R58514 vdd.n16672 vdd.n16671 0.047
R58515 vdd.n19132 vdd.n19130 0.047
R58516 vdd.n19117 vdd.n19115 0.047
R58517 vdd.n19101 vdd.n19099 0.047
R58518 vdd.n19085 vdd.n19083 0.047
R58519 vdd.n19069 vdd.n19067 0.047
R58520 vdd.n19053 vdd.n19051 0.047
R58521 vdd.n19037 vdd.n19035 0.047
R58522 vdd.n19018 vdd.n19006 0.047
R58523 vdd.n19002 vdd.n18990 0.047
R58524 vdd.n18986 vdd.n18974 0.047
R58525 vdd.n18970 vdd.n18958 0.047
R58526 vdd.n18954 vdd.n18942 0.047
R58527 vdd.n18938 vdd.n18926 0.047
R58528 vdd.n18922 vdd.n18910 0.047
R58529 vdd.n18874 vdd.n18872 0.047
R58530 vdd.n18858 vdd.n18856 0.047
R58531 vdd.n18842 vdd.n18840 0.047
R58532 vdd.n18826 vdd.n18824 0.047
R58533 vdd.n18810 vdd.n18808 0.047
R58534 vdd.n18794 vdd.n18792 0.047
R58535 vdd.n18778 vdd.n18776 0.047
R58536 vdd.n18759 vdd.n18747 0.047
R58537 vdd.n18743 vdd.n18731 0.047
R58538 vdd.n18727 vdd.n18715 0.047
R58539 vdd.n18711 vdd.n18699 0.047
R58540 vdd.n18695 vdd.n18683 0.047
R58541 vdd.n18679 vdd.n18667 0.047
R58542 vdd.n18663 vdd.n18651 0.047
R58543 vdd.n18615 vdd.n18613 0.047
R58544 vdd.n18599 vdd.n18597 0.047
R58545 vdd.n18583 vdd.n18581 0.047
R58546 vdd.n18567 vdd.n18565 0.047
R58547 vdd.n18551 vdd.n18549 0.047
R58548 vdd.n18535 vdd.n18533 0.047
R58549 vdd.n18519 vdd.n18517 0.047
R58550 vdd.n21619 vdd.n21599 0.047
R58551 vdd.n21595 vdd.n21583 0.047
R58552 vdd.n21579 vdd.n21567 0.047
R58553 vdd.n21563 vdd.n21551 0.047
R58554 vdd.n21547 vdd.n21535 0.047
R58555 vdd.n21499 vdd.n21497 0.047
R58556 vdd.n21483 vdd.n21481 0.047
R58557 vdd.n21467 vdd.n21465 0.047
R58558 vdd.n21451 vdd.n21449 0.047
R58559 vdd.n21435 vdd.n21433 0.047
R58560 vdd.n21419 vdd.n21417 0.047
R58561 vdd.n21403 vdd.n21401 0.047
R58562 vdd.n21384 vdd.n21372 0.047
R58563 vdd.n21368 vdd.n21356 0.047
R58564 vdd.n21352 vdd.n21340 0.047
R58565 vdd.n21336 vdd.n21324 0.047
R58566 vdd.n21320 vdd.n21308 0.047
R58567 vdd.n21304 vdd.n21292 0.047
R58568 vdd.n21288 vdd.n21276 0.047
R58569 vdd.n21240 vdd.n21238 0.047
R58570 vdd.n21224 vdd.n21222 0.047
R58571 vdd.n21208 vdd.n21206 0.047
R58572 vdd.n21192 vdd.n21190 0.047
R58573 vdd.n21176 vdd.n21174 0.047
R58574 vdd.n21160 vdd.n21158 0.047
R58575 vdd.n21144 vdd.n21142 0.047
R58576 vdd.n21125 vdd.n21113 0.047
R58577 vdd.n21109 vdd.n21097 0.047
R58578 vdd.n16786 vdd.n16785 0.047
R58579 vdd.n15280 vdd.n15279 0.047
R58580 vdd.n15294 vdd.n15293 0.047
R58581 vdd.n15330 vdd.n15329 0.047
R58582 vdd.n15344 vdd.n15343 0.047
R58583 vdd.n15359 vdd.n15358 0.047
R58584 vdd.n15373 vdd.n15372 0.047
R58585 vdd.n15387 vdd.n15386 0.047
R58586 vdd.n15401 vdd.n15400 0.047
R58587 vdd.n15416 vdd.n15415 0.047
R58588 vdd.n15420 vdd.n15419 0.047
R58589 vdd.n15434 vdd.n15433 0.047
R58590 vdd.n15448 vdd.n15447 0.047
R58591 vdd.n15468 vdd.n15467 0.047
R58592 vdd.n15485 vdd.n15484 0.047
R58593 vdd.n15502 vdd.n15501 0.047
R58594 vdd.n15519 vdd.n15518 0.047
R58595 vdd.n15564 vdd.n15563 0.047
R58596 vdd.n15581 vdd.n15580 0.047
R58597 vdd.n15598 vdd.n15597 0.047
R58598 vdd.n15615 vdd.n15614 0.047
R58599 vdd.n15632 vdd.n15631 0.047
R58600 vdd.n15649 vdd.n15648 0.047
R58601 vdd.n15666 vdd.n15665 0.047
R58602 vdd.n15670 vdd.n15669 0.047
R58603 vdd.n15687 vdd.n15686 0.047
R58604 vdd.n15704 vdd.n15703 0.047
R58605 vdd.n15724 vdd.n15723 0.047
R58606 vdd.n15741 vdd.n15740 0.047
R58607 vdd.n15758 vdd.n15757 0.047
R58608 vdd.n15775 vdd.n15774 0.047
R58609 vdd.n15820 vdd.n15819 0.047
R58610 vdd.n15837 vdd.n15836 0.047
R58611 vdd.n15854 vdd.n15853 0.047
R58612 vdd.n15871 vdd.n15870 0.047
R58613 vdd.n15888 vdd.n15887 0.047
R58614 vdd.n15905 vdd.n15904 0.047
R58615 vdd.n15922 vdd.n15921 0.047
R58616 vdd.n15926 vdd.n15925 0.047
R58617 vdd.n15943 vdd.n15942 0.047
R58618 vdd.n15960 vdd.n15959 0.047
R58619 vdd.n15980 vdd.n15979 0.047
R58620 vdd.n15997 vdd.n15996 0.047
R58621 vdd.n16014 vdd.n16013 0.047
R58622 vdd.n16031 vdd.n16030 0.047
R58623 vdd.n16076 vdd.n16075 0.047
R58624 vdd.n16093 vdd.n16092 0.047
R58625 vdd.n16110 vdd.n16109 0.047
R58626 vdd.n16127 vdd.n16126 0.047
R58627 vdd.n16144 vdd.n16143 0.047
R58628 vdd.n16161 vdd.n16160 0.047
R58629 vdd.n16178 vdd.n16177 0.047
R58630 vdd.n16182 vdd.n16181 0.047
R58631 vdd.n16199 vdd.n16198 0.047
R58632 vdd.n16216 vdd.n16215 0.047
R58633 vdd.n16236 vdd.n16235 0.047
R58634 vdd.n16253 vdd.n16252 0.047
R58635 vdd.n16270 vdd.n16269 0.047
R58636 vdd.n16287 vdd.n16286 0.047
R58637 vdd.n16332 vdd.n16331 0.047
R58638 vdd.n16349 vdd.n16348 0.047
R58639 vdd.n16366 vdd.n16365 0.047
R58640 vdd.n16383 vdd.n16382 0.047
R58641 vdd.n16400 vdd.n16399 0.047
R58642 vdd.n16417 vdd.n16416 0.047
R58643 vdd.n16434 vdd.n16433 0.047
R58644 vdd.n16438 vdd.n16437 0.047
R58645 vdd.n16455 vdd.n16454 0.047
R58646 vdd.n16472 vdd.n16471 0.047
R58647 vdd.n16492 vdd.n16491 0.047
R58648 vdd.n16509 vdd.n16508 0.047
R58649 vdd.n16526 vdd.n16525 0.047
R58650 vdd.n16574 vdd.n16542 0.047
R58651 vdd.n34196 vdd.n34160 0.047
R58652 vdd.n35328 vdd.n35292 0.047
R58653 vdd.n34744 vdd.n34708 0.047
R58654 vdd.n5897 vdd.n5861 0.047
R58655 vdd.n5491 vdd.n5455 0.047
R58656 vdd.n4318 vdd.n4282 0.047
R58657 vdd.n25054 vdd.n25052 0.046
R58658 vdd.n27385 vdd.n27384 0.046
R58659 vdd.n4542 vdd.n4541 0.046
R58660 vdd.n802 vdd.n801 0.046
R58661 vdd.n24930 vdd.n24927 0.046
R58662 vdd.n25514 vdd.n25507 0.046
R58663 vdd.n33304 vdd.n33303 0.046
R58664 vdd.n33626 vdd.n33625 0.046
R58665 vdd.n33805 vdd.n33800 0.046
R58666 vdd.n34278 vdd.n34277 0.046
R58667 vdd.n33972 vdd.n33971 0.046
R58668 vdd.n35128 vdd.n35127 0.046
R58669 vdd.n34993 vdd.n34992 0.046
R58670 vdd.n34544 vdd.n34543 0.046
R58671 vdd.n747 vdd.n746 0.046
R58672 vdd.n657 vdd.n656 0.046
R58673 vdd.n833 vdd.n832 0.046
R58674 vdd.n6257 vdd.n6256 0.046
R58675 vdd.n5740 vdd.n5739 0.046
R58676 vdd.n5290 vdd.n5289 0.046
R58677 vdd.n4615 vdd.n4614 0.046
R58678 vdd.n4569 vdd.n4568 0.046
R58679 vdd.n4121 vdd.n4120 0.046
R58680 vdd.n4185 vdd.n4174 0.046
R58681 vdd.n27471 vdd.n27470 0.046
R58682 vdd.n27366 vdd.n27365 0.046
R58683 vdd.n25995 vdd.n25994 0.046
R58684 vdd.n13751 vdd.n13749 0.046
R58685 vdd.n13798 vdd.n8759 0.046
R58686 vdd.n13796 vdd.n8760 0.046
R58687 vdd.n13814 vdd.n13813 0.046
R58688 vdd.n12579 vdd.n10252 0.046
R58689 vdd.n11728 vdd.n11727 0.046
R58690 vdd.n21077 vdd.n21065 0.046
R58691 vdd.n21061 vdd.n21049 0.046
R58692 vdd.n21045 vdd.n21033 0.046
R58693 vdd.n21029 vdd.n21019 0.046
R58694 vdd.n16791 vdd.n16790 0.046
R58695 vdd.n21802 vdd.n21800 0.046
R58696 vdd.n946 vdd.n945 0.046
R58697 vdd.n27242 vdd.n27208 0.046
R58698 vdd.n25650 vdd.n25646 0.046
R58699 vdd.n24540 vdd.n24539 0.046
R58700 vdd.n24962 vdd.n24961 0.046
R58701 vdd.n34133 vdd.n34132 0.046
R58702 vdd.n34964 vdd.n34963 0.046
R58703 vdd.n5711 vdd.n5710 0.046
R58704 vdd.n24889 vdd.n24888 0.046
R58705 vdd.n24924 vdd.n24923 0.046
R58706 vdd.n298 vdd.n297 0.046
R58707 vdd.n25828 vdd.n25827 0.046
R58708 vdd.n27519 vdd.n27518 0.045
R58709 vdd.n27413 vdd.n27412 0.045
R58710 vdd.n35478 vdd.n35477 0.045
R58711 vdd.n5828 vdd.n5827 0.045
R58712 vdd.n25956 vdd.n25955 0.045
R58713 vdd.n25859 vdd.n25858 0.045
R58714 vdd.n33606 vdd.n33603 0.045
R58715 vdd.n650 vdd.n649 0.045
R58716 vdd.n1122 vdd.n1114 0.045
R58717 vdd.n33380 vdd.n33379 0.045
R58718 vdd.n33390 vdd.n33389 0.045
R58719 vdd.n35543 vdd.n35534 0.045
R58720 vdd.n694 vdd.n693 0.045
R58721 vdd.n703 vdd.n702 0.045
R58722 vdd.n492 vdd.n491 0.045
R58723 vdd.n502 vdd.n501 0.045
R58724 vdd.n408 vdd.n407 0.045
R58725 vdd.n125 vdd.n116 0.045
R58726 vdd.n6015 vdd.n6014 0.045
R58727 vdd.n5105 vdd.n5104 0.045
R58728 vdd.n4671 vdd.n4670 0.045
R58729 vdd.n12580 vdd.n10127 0.045
R58730 vdd.n11478 vdd.n11470 0.045
R58731 vdd.n15056 vdd.n15055 0.045
R58732 vdd.n18308 vdd.n18307 0.045
R58733 vdd.n280 vdd.n279 0.045
R58734 vdd.n4850 vdd.n4849 0.045
R58735 vdd.n25585 vdd.n25581 0.044
R58736 vdd.n4541 vdd.n4540 0.044
R58737 vdd.n38217 vdd.n32814 0.044
R58738 vdd.n33420 vdd.n33419 0.044
R58739 vdd.n33503 vdd.n33502 0.044
R58740 vdd.n33303 vdd.n33301 0.044
R58741 vdd.n33303 vdd.n33300 0.044
R58742 vdd.n33637 vdd.n33634 0.044
R58743 vdd.n33674 vdd.n33671 0.044
R58744 vdd.n33817 vdd.n33814 0.044
R58745 vdd.n33835 vdd.n33832 0.044
R58746 vdd.n33806 vdd.n33805 0.044
R58747 vdd.n34116 vdd.n34113 0.044
R58748 vdd.n34277 vdd.n34274 0.044
R58749 vdd.n34292 vdd.n34291 0.044
R58750 vdd.n34312 vdd.n34309 0.044
R58751 vdd.n34173 vdd.n34172 0.044
R58752 vdd.n34169 vdd.n34167 0.044
R58753 vdd.n34210 vdd.n34207 0.044
R58754 vdd.n33914 vdd.n33913 0.044
R58755 vdd.n33886 vdd.n33885 0.044
R58756 vdd.n34021 vdd.n34020 0.044
R58757 vdd.n35318 vdd.n35317 0.044
R58758 vdd.n35314 vdd.n35309 0.044
R58759 vdd.n35578 vdd.n35575 0.044
R58760 vdd.n35558 vdd.n35557 0.044
R58761 vdd.n35543 vdd.n35540 0.044
R58762 vdd.n35532 vdd.n35531 0.044
R58763 vdd.n35111 vdd.n35110 0.044
R58764 vdd.n35060 vdd.n35059 0.044
R58765 vdd.n35331 vdd.n35291 0.044
R58766 vdd.n34992 vdd.n34929 0.044
R58767 vdd.n34908 vdd.n34907 0.044
R58768 vdd.n35001 vdd.n34904 0.044
R58769 vdd.n34723 vdd.n34722 0.044
R58770 vdd.n34738 vdd.n34733 0.044
R58771 vdd.n34747 vdd.n34707 0.044
R58772 vdd.n34473 vdd.n34472 0.044
R58773 vdd.n34524 vdd.n34523 0.044
R58774 vdd.n34607 vdd.n34596 0.044
R58775 vdd.n993 vdd.n992 0.044
R58776 vdd.n657 vdd.n641 0.044
R58777 vdd.n1131 vdd.n1091 0.044
R58778 vdd.n1140 vdd.n1064 0.044
R58779 vdd.n1128 vdd.n1093 0.044
R58780 vdd.n835 vdd.n822 0.044
R58781 vdd.n811 vdd.n810 0.044
R58782 vdd.n539 vdd.n538 0.044
R58783 vdd.n33 vdd.n32 0.044
R58784 vdd.n256 vdd.n255 0.044
R58785 vdd.n5876 vdd.n5875 0.044
R58786 vdd.n5870 vdd.n5868 0.044
R58787 vdd.n6024 vdd.n5947 0.044
R58788 vdd.n5951 vdd.n5950 0.044
R58789 vdd.n6015 vdd.n5972 0.044
R58790 vdd.n5824 vdd.n5821 0.044
R58791 vdd.n6012 vdd.n5973 0.044
R58792 vdd.n6160 vdd.n6159 0.044
R58793 vdd.n6188 vdd.n6187 0.044
R58794 vdd.n6212 vdd.n6205 0.044
R58795 vdd.n5911 vdd.n5908 0.044
R58796 vdd.n5739 vdd.n5676 0.044
R58797 vdd.n5655 vdd.n5654 0.044
R58798 vdd.n5748 vdd.n5651 0.044
R58799 vdd.n5470 vdd.n5469 0.044
R58800 vdd.n5485 vdd.n5480 0.044
R58801 vdd.n5494 vdd.n5454 0.044
R58802 vdd.n5220 vdd.n5219 0.044
R58803 vdd.n5271 vdd.n5270 0.044
R58804 vdd.n5354 vdd.n5343 0.044
R58805 vdd.n4670 vdd.n4653 0.044
R58806 vdd.n4637 vdd.n4636 0.044
R58807 vdd.n4686 vdd.n4635 0.044
R58808 vdd.n5096 vdd.n5095 0.044
R58809 vdd.n4991 vdd.n4990 0.044
R58810 vdd.n4969 vdd.n4968 0.044
R58811 vdd.n4569 vdd.n4503 0.044
R58812 vdd.n4482 vdd.n4481 0.044
R58813 vdd.n4578 vdd.n4478 0.044
R58814 vdd.n4570 vdd.n4569 0.044
R58815 vdd.n4297 vdd.n4296 0.044
R58816 vdd.n4312 vdd.n4307 0.044
R58817 vdd.n4321 vdd.n4281 0.044
R58818 vdd.n4050 vdd.n4049 0.044
R58819 vdd.n4101 vdd.n4100 0.044
R58820 vdd.n27582 vdd.n27570 0.044
R58821 vdd.n27445 vdd.n27443 0.044
R58822 vdd.n27345 vdd.n27343 0.044
R58823 vdd.n25834 vdd.n25833 0.044
R58824 vdd.n25891 vdd.n25889 0.044
R58825 vdd.n25797 vdd.n25795 0.044
R58826 vdd.n25597 vdd.n25593 0.044
R58827 vdd.n2132 vdd.n2131 0.044
R58828 vdd.n10211 vdd.n10210 0.044
R58829 vdd.n22363 vdd.n22344 0.044
R58830 vdd.n22343 vdd.n22342 0.044
R58831 vdd.n24308 vdd.n24307 0.044
R58832 vdd.n24306 vdd.n24305 0.044
R58833 vdd.n24408 vdd.n24407 0.044
R58834 vdd.n16784 vdd.n16783 0.044
R58835 vdd.n25625 vdd.n25624 0.044
R58836 vdd.n25547 vdd.n25546 0.044
R58837 vdd.n25461 vdd.n25460 0.044
R58838 vdd.n160 vdd.n90 0.044
R58839 vdd.n34247 vdd.n34246 0.044
R58840 vdd.n34381 vdd.n34380 0.044
R58841 vdd.n33984 vdd.n33983 0.044
R58842 vdd.n35146 vdd.n35145 0.044
R58843 vdd.n35513 vdd.n35512 0.044
R58844 vdd.n34980 vdd.n34979 0.044
R58845 vdd.n34804 vdd.n34803 0.044
R58846 vdd.n34561 vdd.n34560 0.044
R58847 vdd.n6272 vdd.n6271 0.044
R58848 vdd.n5993 vdd.n5992 0.044
R58849 vdd.n5727 vdd.n5726 0.044
R58850 vdd.n5551 vdd.n5550 0.044
R58851 vdd.n5308 vdd.n5307 0.044
R58852 vdd.n5141 vdd.n5140 0.044
R58853 vdd.n4557 vdd.n4556 0.044
R58854 vdd.n4139 vdd.n4138 0.044
R58855 vdd.n5047 vdd.n5046 0.043
R58856 vdd.n35477 vdd.n35476 0.043
R58857 vdd.n5829 vdd.n5828 0.043
R58858 vdd.n2796 vdd.n2794 0.043
R58859 vdd.n2811 vdd.n2804 0.043
R58860 vdd.n2977 vdd.n2975 0.043
R58861 vdd.n2992 vdd.n2985 0.043
R58862 vdd.n3158 vdd.n3156 0.043
R58863 vdd.n3173 vdd.n3166 0.043
R58864 vdd.n3339 vdd.n3337 0.043
R58865 vdd.n3354 vdd.n3347 0.043
R58866 vdd.n3520 vdd.n3518 0.043
R58867 vdd.n3535 vdd.n3528 0.043
R58868 vdd.n33773 vdd.n33772 0.043
R58869 vdd.n33933 vdd.n33932 0.043
R58870 vdd.n34021 vdd.n34019 0.043
R58871 vdd.n34027 vdd.n34026 0.043
R58872 vdd.n35544 vdd.n35543 0.043
R58873 vdd.n34607 vdd.n34606 0.043
R58874 vdd.n34611 vdd.n34610 0.043
R58875 vdd.n1132 vdd.n1131 0.043
R58876 vdd.n1128 vdd.n1127 0.043
R58877 vdd.n6016 vdd.n6015 0.043
R58878 vdd.n5354 vdd.n5353 0.043
R58879 vdd.n5358 vdd.n5357 0.043
R58880 vdd.n4566 vdd.n4504 0.043
R58881 vdd.n35916 vdd.n35914 0.043
R58882 vdd.n35935 vdd.n35924 0.043
R58883 vdd.n36147 vdd.n36145 0.043
R58884 vdd.n36166 vdd.n36155 0.043
R58885 vdd.n36378 vdd.n36376 0.043
R58886 vdd.n36397 vdd.n36386 0.043
R58887 vdd.n36609 vdd.n36607 0.043
R58888 vdd.n36628 vdd.n36617 0.043
R58889 vdd.n36840 vdd.n36838 0.043
R58890 vdd.n36859 vdd.n36848 0.043
R58891 vdd.n37914 vdd.n37903 0.043
R58892 vdd.n37895 vdd.n37893 0.043
R58893 vdd.n37683 vdd.n37672 0.043
R58894 vdd.n37664 vdd.n37662 0.043
R58895 vdd.n28337 vdd.n28335 0.043
R58896 vdd.n28356 vdd.n28345 0.043
R58897 vdd.n28568 vdd.n28566 0.043
R58898 vdd.n28587 vdd.n28576 0.043
R58899 vdd.n28799 vdd.n28797 0.043
R58900 vdd.n1573 vdd.n1566 0.043
R58901 vdd.n1558 vdd.n1556 0.043
R58902 vdd.n1392 vdd.n1385 0.043
R58903 vdd.n1377 vdd.n1375 0.043
R58904 vdd.n26843 vdd.n26841 0.043
R58905 vdd.n26858 vdd.n26851 0.043
R58906 vdd.n27024 vdd.n27022 0.043
R58907 vdd.n27039 vdd.n27032 0.043
R58908 vdd.n27205 vdd.n27203 0.043
R58909 vdd.n25661 vdd.n25660 0.043
R58910 vdd.n31299 vdd.n31297 0.043
R58911 vdd.n10267 vdd.n10266 0.043
R58912 vdd.n10212 vdd.n10067 0.043
R58913 vdd.n12578 vdd.n12577 0.043
R58914 vdd.n10258 vdd.n10254 0.043
R58915 vdd.n11676 vdd.n11671 0.043
R58916 vdd.n11890 vdd.n11799 0.043
R58917 vdd.n22346 vdd.n22345 0.043
R58918 vdd.n15041 vdd.n15040 0.043
R58919 vdd.n16683 vdd.n16682 0.043
R58920 vdd.n15063 vdd.n15062 0.043
R58921 vdd.n16793 vdd.n16792 0.043
R58922 vdd.n21855 vdd.n21854 0.043
R58923 vdd.n21981 vdd.n21890 0.043
R58924 vdd.n5088 vdd.n5085 0.043
R58925 vdd.n4922 vdd.n4889 0.043
R58926 vdd.n27622 vdd.n27621 0.042
R58927 vdd.n25454 vdd.n25452 0.042
R58928 vdd.n34111 vdd.n34110 0.042
R58929 vdd.n35496 vdd.n35495 0.042
R58930 vdd.n34944 vdd.n34943 0.042
R58931 vdd.n5997 vdd.n5996 0.042
R58932 vdd.n5691 vdd.n5690 0.042
R58933 vdd.n4518 vdd.n4517 0.042
R58934 vdd.n27651 vdd.n27650 0.042
R58935 vdd.n26073 vdd.n26072 0.042
R58936 vdd.n331 vdd.n330 0.042
R58937 vdd.n5117 vdd.n5116 0.042
R58938 vdd.n5105 vdd.n5102 0.042
R58939 vdd.n5013 vdd.n5012 0.042
R58940 vdd.n5007 vdd.n5006 0.042
R58941 vdd.n4665 vdd.n4664 0.042
R58942 vdd.n25604 vdd.n25603 0.042
R58943 vdd.n25559 vdd.n25558 0.042
R58944 vdd.n11762 vdd.n11761 0.042
R58945 vdd.n35212 vdd.n35136 0.042
R58946 vdd.n6336 vdd.n6335 0.042
R58947 vdd.n22364 vdd.n22363 0.042
R58948 vdd.n24309 vdd.n24308 0.042
R58949 vdd.n35597 vdd.n35593 0.042
R58950 vdd.n35333 vdd.n35280 0.042
R58951 vdd.n6032 vdd.n5927 0.042
R58952 vdd.n5914 vdd.n5913 0.042
R58953 vdd.n25538 vdd.n25536 0.042
R58954 vdd.n26043 vdd.n26042 0.042
R58955 vdd.n33337 vdd.n33293 0.042
R58956 vdd.n666 vdd.n614 0.042
R58957 vdd.n555 vdd.n552 0.042
R58958 vdd.n277 vdd.n276 0.041
R58959 vdd.n25913 vdd.n25912 0.041
R58960 vdd.n34250 vdd.n34247 0.041
R58961 vdd.n35516 vdd.n35513 0.041
R58962 vdd.n35436 vdd.n35433 0.041
R58963 vdd.n34983 vdd.n34980 0.041
R58964 vdd.n6006 vdd.n5993 0.041
R58965 vdd.n6116 vdd.n6112 0.041
R58966 vdd.n5730 vdd.n5727 0.041
R58967 vdd.n4742 vdd.n4726 0.041
R58968 vdd.n4560 vdd.n4557 0.041
R58969 vdd.n4413 vdd.n4410 0.041
R58970 vdd.n33638 vdd.n33637 0.041
R58971 vdd.n33626 vdd.n33617 0.041
R58972 vdd.n34266 vdd.n34265 0.041
R58973 vdd.n35113 vdd.n35112 0.041
R58974 vdd.n35391 vdd.n35390 0.041
R58975 vdd.n34989 vdd.n34930 0.041
R58976 vdd.n879 vdd.n876 0.041
R58977 vdd.n6149 vdd.n6148 0.041
R58978 vdd.n6126 vdd.n6125 0.041
R58979 vdd.n5736 vdd.n5677 0.041
R58980 vdd.n4185 vdd.n4184 0.041
R58981 vdd.n4189 vdd.n4188 0.041
R58982 vdd.n27358 vdd.n27357 0.041
R58983 vdd.n25810 vdd.n25809 0.041
R58984 vdd.n31685 vdd.n31684 0.041
R58985 vdd.n10250 vdd.n10249 0.041
R58986 vdd.n12600 vdd.n10095 0.041
R58987 vdd.n10142 vdd.n10136 0.041
R58988 vdd.n22344 vdd.n22343 0.041
R58989 vdd.n22342 vdd.n22341 0.041
R58990 vdd.n22133 vdd.n22132 0.041
R58991 vdd.n24307 vdd.n24306 0.041
R58992 vdd.n24305 vdd.n24304 0.041
R58993 vdd.n16604 vdd.n16603 0.041
R58994 vdd.n16743 vdd.n16741 0.041
R58995 vdd.n4202 vdd.n4126 0.041
R58996 vdd.n4586 vdd.n4458 0.041
R58997 vdd.n4323 vdd.n4270 0.041
R58998 vdd.n29953 vdd.n29952 0.041
R58999 vdd.n33353 vdd.n33352 0.041
R59000 vdd.n33677 vdd.n33676 0.041
R59001 vdd.n34432 vdd.n34431 0.041
R59002 vdd.n34862 vdd.n34861 0.041
R59003 vdd.n5609 vdd.n5608 0.041
R59004 vdd.n4436 vdd.n4435 0.041
R59005 vdd.n27503 vdd.n27502 0.041
R59006 vdd.n27402 vdd.n27401 0.041
R59007 vdd.n27467 vdd.n27466 0.041
R59008 vdd.n25940 vdd.n25939 0.04
R59009 vdd.n25848 vdd.n25847 0.04
R59010 vdd.n2881 vdd.n2879 0.04
R59011 vdd.n2902 vdd.n2900 0.04
R59012 vdd.n3062 vdd.n3060 0.04
R59013 vdd.n3083 vdd.n3081 0.04
R59014 vdd.n3243 vdd.n3241 0.04
R59015 vdd.n3264 vdd.n3262 0.04
R59016 vdd.n3424 vdd.n3422 0.04
R59017 vdd.n3445 vdd.n3443 0.04
R59018 vdd.n3605 vdd.n3603 0.04
R59019 vdd.n3626 vdd.n3624 0.04
R59020 vdd.n33407 vdd.n33406 0.04
R59021 vdd.n33473 vdd.n33471 0.04
R59022 vdd.n33481 vdd.n33477 0.04
R59023 vdd.n33612 vdd.n33611 0.04
R59024 vdd.n34144 vdd.n34099 0.04
R59025 vdd.n34266 vdd.n34263 0.04
R59026 vdd.n34170 vdd.n34169 0.04
R59027 vdd.n33884 vdd.n33881 0.04
R59028 vdd.n33870 vdd.n33866 0.04
R59029 vdd.n34350 vdd.n34346 0.04
R59030 vdd.n34407 vdd.n34406 0.04
R59031 vdd.n34021 vdd.n34009 0.04
R59032 vdd.n35183 vdd.n35171 0.04
R59033 vdd.n35266 vdd.n35260 0.04
R59034 vdd.n35121 vdd.n35117 0.04
R59035 vdd.n35109 vdd.n35106 0.04
R59036 vdd.n35420 vdd.n35419 0.04
R59037 vdd.n35368 vdd.n35364 0.04
R59038 vdd.n35183 vdd.n35181 0.04
R59039 vdd.n35189 vdd.n35188 0.04
R59040 vdd.n34685 vdd.n34676 0.04
R59041 vdd.n34989 vdd.n34988 0.04
R59042 vdd.n34739 vdd.n34738 0.04
R59043 vdd.n34824 vdd.n34823 0.04
R59044 vdd.n34522 vdd.n34519 0.04
R59045 vdd.n34534 vdd.n34530 0.04
R59046 vdd.n34778 vdd.n34774 0.04
R59047 vdd.n34830 vdd.n34829 0.04
R59048 vdd.n34607 vdd.n34595 0.04
R59049 vdd.n731 vdd.n730 0.04
R59050 vdd.n786 vdd.n711 0.04
R59051 vdd.n966 vdd.n962 0.04
R59052 vdd.n648 vdd.n647 0.04
R59053 vdd.n661 vdd.n660 0.04
R59054 vdd.n1105 vdd.n1104 0.04
R59055 vdd.n879 vdd.n878 0.04
R59056 vdd.n487 vdd.n485 0.04
R59057 vdd.n4 vdd.n0 0.04
R59058 vdd.n81 vdd.n15 0.04
R59059 vdd.n422 vdd.n421 0.04
R59060 vdd.n125 vdd.n122 0.04
R59061 vdd.n140 vdd.n139 0.04
R59062 vdd.n334 vdd.n333 0.04
R59063 vdd.n330 vdd.n328 0.04
R59064 vdd.n368 vdd.n365 0.04
R59065 vdd.n6318 vdd.n6306 0.04
R59066 vdd.n5833 vdd.n5804 0.04
R59067 vdd.n6144 vdd.n6140 0.04
R59068 vdd.n6158 vdd.n6155 0.04
R59069 vdd.n6056 vdd.n6052 0.04
R59070 vdd.n6217 vdd.n6216 0.04
R59071 vdd.n6318 vdd.n6317 0.04
R59072 vdd.n6322 vdd.n6321 0.04
R59073 vdd.n5432 vdd.n5423 0.04
R59074 vdd.n5736 vdd.n5735 0.04
R59075 vdd.n5486 vdd.n5485 0.04
R59076 vdd.n5571 vdd.n5570 0.04
R59077 vdd.n5269 vdd.n5266 0.04
R59078 vdd.n5281 vdd.n5277 0.04
R59079 vdd.n5525 vdd.n5521 0.04
R59080 vdd.n5577 vdd.n5576 0.04
R59081 vdd.n5354 vdd.n5342 0.04
R59082 vdd.n5105 vdd.n5103 0.04
R59083 vdd.n4805 vdd.n4801 0.04
R59084 vdd.n4794 vdd.n4790 0.04
R59085 vdd.n4967 vdd.n4964 0.04
R59086 vdd.n4956 vdd.n4952 0.04
R59087 vdd.n4922 vdd.n4898 0.04
R59088 vdd.n4259 vdd.n4253 0.04
R59089 vdd.n4397 vdd.n4396 0.04
R59090 vdd.n4099 vdd.n4096 0.04
R59091 vdd.n4111 vdd.n4107 0.04
R59092 vdd.n4352 vdd.n4348 0.04
R59093 vdd.n4103 vdd.n4102 0.04
R59094 vdd.n4367 vdd.n4366 0.04
R59095 vdd.n4185 vdd.n4173 0.04
R59096 vdd.n36023 vdd.n36021 0.04
R59097 vdd.n36051 vdd.n36049 0.04
R59098 vdd.n36254 vdd.n36252 0.04
R59099 vdd.n36282 vdd.n36280 0.04
R59100 vdd.n36485 vdd.n36483 0.04
R59101 vdd.n36513 vdd.n36511 0.04
R59102 vdd.n36716 vdd.n36714 0.04
R59103 vdd.n36744 vdd.n36742 0.04
R59104 vdd.n36947 vdd.n36945 0.04
R59105 vdd.n38030 vdd.n38028 0.04
R59106 vdd.n38002 vdd.n38000 0.04
R59107 vdd.n37799 vdd.n37797 0.04
R59108 vdd.n37771 vdd.n37769 0.04
R59109 vdd.n28213 vdd.n28211 0.04
R59110 vdd.n28241 vdd.n28239 0.04
R59111 vdd.n28444 vdd.n28442 0.04
R59112 vdd.n28472 vdd.n28470 0.04
R59113 vdd.n28675 vdd.n28673 0.04
R59114 vdd.n28703 vdd.n28701 0.04
R59115 vdd.n1664 vdd.n1662 0.04
R59116 vdd.n1643 vdd.n1641 0.04
R59117 vdd.n1483 vdd.n1481 0.04
R59118 vdd.n1462 vdd.n1460 0.04
R59119 vdd.n1302 vdd.n1300 0.04
R59120 vdd.n26768 vdd.n26766 0.04
R59121 vdd.n26928 vdd.n26926 0.04
R59122 vdd.n26949 vdd.n26947 0.04
R59123 vdd.n27109 vdd.n27107 0.04
R59124 vdd.n27130 vdd.n27128 0.04
R59125 vdd.n27279 vdd.n27278 0.04
R59126 vdd.n27579 vdd.n27576 0.04
R59127 vdd.n27588 vdd.n27584 0.04
R59128 vdd.n25725 vdd.n25724 0.04
R59129 vdd.n25692 vdd.n25689 0.04
R59130 vdd.n26004 vdd.n26000 0.04
R59131 vdd.n25409 vdd.n25408 0.04
R59132 vdd.n25459 vdd.n25458 0.04
R59133 vdd.n25447 vdd.n25446 0.04
R59134 vdd.n12600 vdd.n10077 0.04
R59135 vdd.n11675 vdd.n11672 0.04
R59136 vdd.n11743 vdd.n11725 0.04
R59137 vdd.n11735 vdd.n11725 0.04
R59138 vdd.n11828 vdd.n11827 0.04
R59139 vdd.n11829 vdd.n11828 0.04
R59140 vdd.n22079 vdd.n22078 0.04
R59141 vdd.n16743 vdd.n16691 0.04
R59142 vdd.n21825 vdd.n21820 0.04
R59143 vdd.n21820 vdd.n21812 0.04
R59144 vdd.n21919 vdd.n21918 0.04
R59145 vdd.n21920 vdd.n21919 0.04
R59146 vdd.n25032 vdd.n25030 0.04
R59147 vdd.n25019 vdd.n25017 0.04
R59148 vdd.n24607 vdd.n24605 0.04
R59149 vdd.n24595 vdd.n24593 0.04
R59150 vdd.n5166 vdd.n5069 0.04
R59151 vdd.n4927 vdd.n4878 0.04
R59152 vdd.n4696 vdd.n4693 0.04
R59153 vdd.n33445 vdd.n33392 0.04
R59154 vdd.n563 vdd.n562 0.04
R59155 vdd.n34312 vdd.n34242 0.04
R59156 vdd.n35578 vdd.n35469 0.04
R59157 vdd.n35001 vdd.n34895 0.04
R59158 vdd.n6024 vdd.n5938 0.04
R59159 vdd.n5748 vdd.n5642 0.04
R59160 vdd.n4686 vdd.n4683 0.04
R59161 vdd.n4578 vdd.n4469 0.04
R59162 vdd.n4895 vdd.n4894 0.04
R59163 vdd.n35045 vdd.n35044 0.039
R59164 vdd.n35457 vdd.n35456 0.039
R59165 vdd.n545 vdd.n544 0.039
R59166 vdd.n401 vdd.n400 0.039
R59167 vdd.n74 vdd.n73 0.039
R59168 vdd.n137 vdd.n136 0.039
R59169 vdd.n114 vdd.n113 0.039
R59170 vdd.n303 vdd.n302 0.039
R59171 vdd.n6243 vdd.n6242 0.039
R59172 vdd.n6073 vdd.n6072 0.039
R59173 vdd.n5007 vdd.n5005 0.039
R59174 vdd.n4715 vdd.n4714 0.039
R59175 vdd.n5053 vdd.n5052 0.039
R59176 vdd.n4665 vdd.n4663 0.039
R59177 vdd.n27302 vdd.n27301 0.039
R59178 vdd.n25754 vdd.n25753 0.039
R59179 vdd.n25262 vdd.n25260 0.039
R59180 vdd.n25262 vdd.n25261 0.039
R59181 vdd.n25262 vdd.n7981 0.039
R59182 vdd.n38217 ldomc_0.pmosm_0.vdd 0.039
R59183 vdd.n10143 vdd.n10142 0.039
R59184 vdd.n16706 vdd.n16705 0.039
R59185 vdd.n34051 vdd.n34049 0.039
R59186 vdd.n34625 vdd.n34549 0.039
R59187 vdd.n5372 vdd.n5296 0.039
R59188 vdd.n34331 vdd.n34327 0.039
R59189 vdd.n34213 vdd.n34212 0.039
R59190 vdd.n35009 vdd.n34884 0.039
R59191 vdd.n34749 vdd.n34696 0.039
R59192 vdd.n5756 vdd.n5631 0.039
R59193 vdd.n5496 vdd.n5443 0.039
R59194 vdd.n764 vdd.n760 0.039
R59195 vdd.n459 vdd.n455 0.039
R59196 vdd.n176 vdd.n175 0.039
R59197 vdd.n371 vdd.n370 0.039
R59198 vdd.n60 vdd.n57 0.039
R59199 vdd.n671 vdd.n603 0.039
R59200 vdd.n1142 vdd.n1054 0.039
R59201 vdd.n25516 vdd.n25515 0.038
R59202 vdd.n2785 vdd.n2783 0.038
R59203 vdd.n2822 vdd.n2815 0.038
R59204 vdd.n2966 vdd.n2964 0.038
R59205 vdd.n3003 vdd.n2996 0.038
R59206 vdd.n3147 vdd.n3145 0.038
R59207 vdd.n3184 vdd.n3177 0.038
R59208 vdd.n3328 vdd.n3326 0.038
R59209 vdd.n3365 vdd.n3358 0.038
R59210 vdd.n3509 vdd.n3507 0.038
R59211 vdd.n3546 vdd.n3539 0.038
R59212 vdd.n3657 vdd.n3626 0.038
R59213 vdd.n1759 vdd.n1752 0.038
R59214 vdd.n33314 vdd.n33313 0.038
R59215 vdd.n33557 vdd.n33556 0.038
R59216 vdd.n33773 vdd.n33770 0.038
R59217 vdd.n33875 vdd.n33874 0.038
R59218 vdd.n34423 vdd.n34422 0.038
R59219 vdd.n34526 vdd.n34525 0.038
R59220 vdd.n34793 vdd.n34792 0.038
R59221 vdd.n835 vdd.n815 0.038
R59222 vdd.n5273 vdd.n5272 0.038
R59223 vdd.n5540 vdd.n5539 0.038
R59224 vdd.n4566 vdd.n4565 0.038
R59225 vdd.n4313 vdd.n4312 0.038
R59226 vdd.n4403 vdd.n4402 0.038
R59227 vdd.n4025 vdd.n4024 0.038
R59228 vdd.n4442 vdd.n4441 0.038
R59229 vdd.n38153 vdd.n38143 0.038
R59230 vdd.n35902 vdd.n35900 0.038
R59231 vdd.n35949 vdd.n35939 0.038
R59232 vdd.n36133 vdd.n36131 0.038
R59233 vdd.n36180 vdd.n36170 0.038
R59234 vdd.n36364 vdd.n36362 0.038
R59235 vdd.n36411 vdd.n36401 0.038
R59236 vdd.n36595 vdd.n36593 0.038
R59237 vdd.n36642 vdd.n36632 0.038
R59238 vdd.n36826 vdd.n36824 0.038
R59239 vdd.n36873 vdd.n36863 0.038
R59240 vdd.n38112 vdd.n38110 0.038
R59241 vdd.n37928 vdd.n37918 0.038
R59242 vdd.n37881 vdd.n37879 0.038
R59243 vdd.n37697 vdd.n37687 0.038
R59244 vdd.n37650 vdd.n37648 0.038
R59245 vdd.n28323 vdd.n28321 0.038
R59246 vdd.n28370 vdd.n28360 0.038
R59247 vdd.n28554 vdd.n28552 0.038
R59248 vdd.n28601 vdd.n28591 0.038
R59249 vdd.n28785 vdd.n28783 0.038
R59250 vdd.n1728 vdd.n1726 0.038
R59251 vdd.n1584 vdd.n1577 0.038
R59252 vdd.n1547 vdd.n1545 0.038
R59253 vdd.n1403 vdd.n1396 0.038
R59254 vdd.n1366 vdd.n1364 0.038
R59255 vdd.n26832 vdd.n26830 0.038
R59256 vdd.n26869 vdd.n26862 0.038
R59257 vdd.n27013 vdd.n27011 0.038
R59258 vdd.n27050 vdd.n27043 0.038
R59259 vdd.n27194 vdd.n27192 0.038
R59260 vdd.n25627 vdd.n25626 0.038
R59261 vdd.n25549 vdd.n25548 0.038
R59262 vdd.n25463 vdd.n25462 0.038
R59263 vdd.n31304 vdd.n31014 0.038
R59264 vdd.n31104 vdd.n31102 0.038
R59265 vdd.n12600 vdd.n10071 0.038
R59266 vdd.n10130 vdd.n10129 0.038
R59267 vdd.n12578 vdd.n10126 0.038
R59268 vdd.n11799 vdd.n11798 0.038
R59269 vdd.n11916 vdd.n11662 0.038
R59270 vdd.n16743 vdd.n16596 0.038
R59271 vdd.n16674 vdd.n16673 0.038
R59272 vdd.n15062 vdd.n15061 0.038
R59273 vdd.n21890 vdd.n21889 0.038
R59274 vdd.n22002 vdd.n21878 0.038
R59275 vdd.n24861 bandgapmd_0.bg_stupm_0.vdd 0.038
R59276 vdd.n24876 vdd.n24875 0.038
R59277 vdd.n34051 vdd.n34048 0.038
R59278 vdd.n34625 vdd.n34623 0.038
R59279 vdd.n688 vdd.n687 0.038
R59280 vdd.n5372 vdd.n5370 0.038
R59281 vdd.n764 vdd.n759 0.038
R59282 vdd.n34304 vdd.n34303 0.038
R59283 vdd.n33903 vdd.n33902 0.038
R59284 vdd.n35570 vdd.n35569 0.038
R59285 vdd.n35072 vdd.n35071 0.038
R59286 vdd.n34899 vdd.n34898 0.038
R59287 vdd.n34485 vdd.n34484 0.038
R59288 vdd.n5942 vdd.n5941 0.038
R59289 vdd.n6177 vdd.n6176 0.038
R59290 vdd.n5646 vdd.n5645 0.038
R59291 vdd.n5232 vdd.n5231 0.038
R59292 vdd.n4630 vdd.n4629 0.038
R59293 vdd.n5085 vdd.n5084 0.038
R59294 vdd.n4982 vdd.n4981 0.038
R59295 vdd.n4473 vdd.n4472 0.038
R59296 vdd.n4062 vdd.n4061 0.038
R59297 vdd.n25652 vdd.n25650 0.038
R59298 vdd.n34077 vdd.n34076 0.038
R59299 vdd.n35236 vdd.n35235 0.038
R59300 vdd.n34649 vdd.n34648 0.038
R59301 vdd.n5779 vdd.n5778 0.038
R59302 vdd.n5396 vdd.n5395 0.038
R59303 vdd.n4226 vdd.n4225 0.038
R59304 vdd.n25644 vdd.n25643 0.037
R59305 vdd.n34289 vdd.n34288 0.037
R59306 vdd.n33961 vdd.n33960 0.037
R59307 vdd.n34420 vdd.n34419 0.037
R59308 vdd.n35532 vdd.n35529 0.037
R59309 vdd.n35275 vdd.n35244 0.037
R59310 vdd.n35426 vdd.n35425 0.037
R59311 vdd.n35125 vdd.n35124 0.037
R59312 vdd.n35315 vdd.n35314 0.037
R59313 vdd.n34996 vdd.n34995 0.037
R59314 vdd.n34513 vdd.n34512 0.037
R59315 vdd.n34853 vdd.n34852 0.037
R59316 vdd.n750 vdd.n749 0.037
R59317 vdd.n835 vdd.n823 0.037
R59318 vdd.n5841 vdd.n5840 0.037
R59319 vdd.n6012 vdd.n6011 0.037
R59320 vdd.n6139 vdd.n6138 0.037
R59321 vdd.n6212 vdd.n6211 0.037
R59322 vdd.n5871 vdd.n5870 0.037
R59323 vdd.n5743 vdd.n5742 0.037
R59324 vdd.n5260 vdd.n5259 0.037
R59325 vdd.n5600 vdd.n5599 0.037
R59326 vdd.n4786 vdd.n4785 0.037
R59327 vdd.n4971 vdd.n4970 0.037
R59328 vdd.n32463 vdd.n32433 0.037
R59329 vdd.n32188 vdd.n31563 0.037
R59330 vdd.n31304 vdd.n30998 0.037
R59331 vdd.n31808 vdd.n31719 0.037
R59332 vdd.n31729 vdd.n31728 0.037
R59333 vdd.n12600 vdd.n10089 0.037
R59334 vdd.n11696 vdd.n11695 0.037
R59335 vdd.n11868 vdd.n11810 0.037
R59336 vdd.n11888 vdd.n11887 0.037
R59337 ldomc_0.otaldom_0.vdd vdd.n8151 0.037
R59338 vdd.n22216 vdd.n22215 0.037
R59339 vdd.n16743 vdd.n16731 0.037
R59340 vdd.n19987 bandgapmd_0.otam_1.vdd 0.037
R59341 vdd.n21797 vdd.n21796 0.037
R59342 vdd.n21959 vdd.n21901 0.037
R59343 vdd.n21979 vdd.n21978 0.037
R59344 vdd.n578 vdd.n577 0.037
R59345 vdd.n5166 vdd.n5165 0.037
R59346 vdd.n4927 vdd.n4926 0.037
R59347 vdd.n34331 vdd.n34326 0.037
R59348 vdd.n34213 vdd.n34211 0.037
R59349 vdd.n35009 vdd.n35005 0.037
R59350 vdd.n34749 vdd.n34748 0.037
R59351 vdd.n785 vdd.n784 0.037
R59352 vdd.n5756 vdd.n5752 0.037
R59353 vdd.n5496 vdd.n5495 0.037
R59354 vdd.n33844 vdd.n33843 0.037
R59355 vdd.n459 vdd.n454 0.037
R59356 vdd.n176 vdd.n174 0.037
R59357 vdd.n371 vdd.n369 0.037
R59358 vdd.n671 vdd.n670 0.037
R59359 vdd.n1142 vdd.n1141 0.037
R59360 vdd.n33435 vdd.n33432 0.037
R59361 vdd.n33543 vdd.n33540 0.037
R59362 vdd.n33594 vdd.n33591 0.037
R59363 vdd.n755 vdd.n729 0.037
R59364 vdd.n1019 vdd.n1016 0.037
R59365 vdd.n440 vdd.n389 0.037
R59366 vdd.n32105 vdd.n32104 0.036
R59367 vdd.n32527 vdd.n32526 0.036
R59368 vdd.n27850 vdd.n27849 0.036
R59369 vdd.n25633 vdd.n25631 0.036
R59370 vdd.n33373 vdd.n33372 0.036
R59371 vdd.n33317 vdd.n33316 0.036
R59372 vdd.n33297 vdd.n33296 0.036
R59373 vdd.n33514 vdd.n33513 0.036
R59374 vdd.n33738 vdd.n33737 0.036
R59375 vdd.n33757 vdd.n33738 0.036
R59376 vdd.n33626 vdd.n33623 0.036
R59377 vdd.n33641 vdd.n33640 0.036
R59378 vdd.n33615 vdd.n33614 0.036
R59379 vdd.n33809 vdd.n33808 0.036
R59380 vdd.n33805 vdd.n33803 0.036
R59381 vdd.n33824 vdd.n33821 0.036
R59382 vdd.n33841 vdd.n33838 0.036
R59383 vdd.n34266 vdd.n34264 0.036
R59384 vdd.n34179 vdd.n34178 0.036
R59385 vdd.n34196 vdd.n34193 0.036
R59386 vdd.n34187 vdd.n34186 0.036
R59387 vdd.n34363 vdd.n34359 0.036
R59388 vdd.n34365 vdd.n34364 0.036
R59389 vdd.n34433 vdd.n34421 0.036
R59390 vdd.n34371 vdd.n34370 0.036
R59391 vdd.n33958 vdd.n33957 0.036
R59392 vdd.n34367 vdd.n34366 0.036
R59393 vdd.n35532 vdd.n35530 0.036
R59394 vdd.n35265 vdd.n35264 0.036
R59395 vdd.n35394 vdd.n35393 0.036
R59396 vdd.n35379 vdd.n35375 0.036
R59397 vdd.n35381 vdd.n35380 0.036
R59398 vdd.n35328 vdd.n35303 0.036
R59399 vdd.n35297 vdd.n35296 0.036
R59400 vdd.n35324 vdd.n35323 0.036
R59401 vdd.n34989 vdd.n34931 0.036
R59402 vdd.n34729 vdd.n34728 0.036
R59403 vdd.n34744 vdd.n34719 0.036
R59404 vdd.n34713 vdd.n34712 0.036
R59405 vdd.n34789 vdd.n34785 0.036
R59406 vdd.n34791 vdd.n34790 0.036
R59407 vdd.n34863 vdd.n34794 0.036
R59408 vdd.n34797 vdd.n34796 0.036
R59409 vdd.n34448 vdd.n34447 0.036
R59410 vdd.n34868 vdd.n34867 0.036
R59411 vdd.n595 vdd.n594 0.036
R59412 vdd.n627 vdd.n626 0.036
R59413 vdd.n995 vdd.n994 0.036
R59414 vdd.n896 vdd.n894 0.036
R59415 vdd.n1128 vdd.n1099 0.036
R59416 vdd.n1078 vdd.n1077 0.036
R59417 vdd.n817 vdd.n816 0.036
R59418 vdd.n832 vdd.n827 0.036
R59419 vdd.n841 vdd.n840 0.036
R59420 vdd.n801 vdd.n799 0.036
R59421 vdd.n527 vdd.n526 0.036
R59422 vdd.n583 vdd.n582 0.036
R59423 vdd.n398 vdd.n397 0.036
R59424 vdd.n419 vdd.n418 0.036
R59425 vdd.n401 vdd.n392 0.036
R59426 vdd.n71 vdd.n70 0.036
R59427 vdd.n111 vdd.n110 0.036
R59428 vdd.n114 vdd.n107 0.036
R59429 vdd.n303 vdd.n300 0.036
R59430 vdd.n349 vdd.n346 0.036
R59431 vdd.n358 vdd.n357 0.036
R59432 vdd.n6012 vdd.n5974 0.036
R59433 vdd.n5806 vdd.n5805 0.036
R59434 vdd.n6212 vdd.n6209 0.036
R59435 vdd.n6085 vdd.n6084 0.036
R59436 vdd.n6069 vdd.n6065 0.036
R59437 vdd.n6071 vdd.n6070 0.036
R59438 vdd.n5897 vdd.n5894 0.036
R59439 vdd.n5888 vdd.n5887 0.036
R59440 vdd.n5882 vdd.n5881 0.036
R59441 vdd.n5736 vdd.n5678 0.036
R59442 vdd.n5476 vdd.n5475 0.036
R59443 vdd.n5491 vdd.n5466 0.036
R59444 vdd.n5460 vdd.n5459 0.036
R59445 vdd.n5536 vdd.n5532 0.036
R59446 vdd.n5538 vdd.n5537 0.036
R59447 vdd.n5610 vdd.n5541 0.036
R59448 vdd.n5544 vdd.n5543 0.036
R59449 vdd.n5195 vdd.n5194 0.036
R59450 vdd.n5615 vdd.n5614 0.036
R59451 vdd.n4665 vdd.n4654 0.036
R59452 vdd.n5126 vdd.n5071 0.036
R59453 vdd.n4838 vdd.n4837 0.036
R59454 vdd.n4827 vdd.n4826 0.036
R59455 vdd.n4784 vdd.n4783 0.036
R59456 vdd.n4782 vdd.n4778 0.036
R59457 vdd.n4760 vdd.n4759 0.036
R59458 vdd.n5007 vdd.n5004 0.036
R59459 vdd.n4770 vdd.n4769 0.036
R59460 vdd.n5050 vdd.n5049 0.036
R59461 vdd.n4676 vdd.n4675 0.036
R59462 vdd.n4896 vdd.n4895 0.036
R59463 vdd.n4909 vdd.n4908 0.036
R59464 vdd.n4918 vdd.n4917 0.036
R59465 vdd.n4566 vdd.n4505 0.036
R59466 vdd.n4265 vdd.n4234 0.036
R59467 vdd.n4303 vdd.n4302 0.036
R59468 vdd.n4318 vdd.n4293 0.036
R59469 vdd.n4287 vdd.n4286 0.036
R59470 vdd.n4363 vdd.n4359 0.036
R59471 vdd.n4365 vdd.n4364 0.036
R59472 vdd.n4437 vdd.n4368 0.036
R59473 vdd.n4371 vdd.n4370 0.036
R59474 vdd.n4115 vdd.n4114 0.036
R59475 vdd.n27476 vdd.n27475 0.036
R59476 vdd.n27490 vdd.n27489 0.036
R59477 vdd.n27333 vdd.n27331 0.036
R59478 vdd.n27325 vdd.n27324 0.036
R59479 vdd.n25714 vdd.n25713 0.036
R59480 vdd.n25927 vdd.n25926 0.036
R59481 vdd.n25785 vdd.n25783 0.036
R59482 vdd.n25777 vdd.n25776 0.036
R59483 vdd.n10208 vdd.n10207 0.036
R59484 vdd.n12577 vdd.n10253 0.036
R59485 vdd.n11621 vdd.n11609 0.036
R59486 vdd.n11619 vdd.n11610 0.036
R59487 vdd.n22117 vdd.n22116 0.036
R59488 vdd.n16736 vdd.n16735 0.036
R59489 vdd.n15063 vdd.n15060 0.036
R59490 vdd.n21695 vdd.n21694 0.036
R59491 vdd.n21692 vdd.n21691 0.036
R59492 vdd.n33368 vdd.n33367 0.036
R59493 vdd.n4202 vdd.n4201 0.036
R59494 vdd.n33466 vdd.n33465 0.036
R59495 vdd.n480 vdd.n479 0.036
R59496 vdd.n4696 vdd.n4692 0.036
R59497 vdd.n4586 vdd.n4582 0.036
R59498 vdd.n4323 vdd.n4322 0.036
R59499 vdd.n33445 vdd.n33441 0.036
R59500 vdd.n845 vdd.n843 0.036
R59501 vdd.n33353 vdd.n33351 0.036
R59502 vdd.n33677 vdd.n33675 0.036
R59503 vdd.n563 vdd.n561 0.036
R59504 vdd.n27631 vdd.n27630 0.036
R59505 vdd.n34124 vdd.n34123 0.036
R59506 vdd.n34415 vdd.n34391 0.036
R59507 vdd.n34042 vdd.n34039 0.036
R59508 vdd.n35204 vdd.n35201 0.036
R59509 vdd.n35502 vdd.n35499 0.036
R59510 vdd.n35442 vdd.n35439 0.036
R59511 vdd.n34969 vdd.n34947 0.036
R59512 vdd.n34845 vdd.n34842 0.036
R59513 vdd.n34619 vdd.n34571 0.036
R59514 vdd.n6330 vdd.n6282 0.036
R59515 vdd.n6003 vdd.n6000 0.036
R59516 vdd.n6119 vdd.n6104 0.036
R59517 vdd.n5716 vdd.n5694 0.036
R59518 vdd.n5592 vdd.n5589 0.036
R59519 vdd.n5366 vdd.n5318 0.036
R59520 vdd.n5151 vdd.n5070 0.036
R59521 vdd.n4755 vdd.n4725 0.036
R59522 vdd.n4546 vdd.n4521 0.036
R59523 vdd.n4419 vdd.n4416 0.036
R59524 vdd.n4197 vdd.n4149 0.036
R59525 vdd.n33941 vdd.n33899 0.036
R59526 vdd.n35082 vdd.n35047 0.036
R59527 vdd.n34495 vdd.n34460 0.036
R59528 vdd.n6225 vdd.n6173 0.036
R59529 vdd.n5242 vdd.n5207 0.036
R59530 vdd.n5074 vdd.n5072 0.036
R59531 vdd.n5028 vdd.n5025 0.036
R59532 vdd.n4072 vdd.n4037 0.036
R59533 vdd.n25603 vdd.n25601 0.036
R59534 vdd.n34186 vdd.n34185 0.036
R59535 vdd.n35296 vdd.n35295 0.036
R59536 vdd.n34712 vdd.n34711 0.036
R59537 vdd.n5887 vdd.n5886 0.036
R59538 vdd.n5459 vdd.n5458 0.036
R59539 vdd.n4286 vdd.n4285 0.036
R59540 vdd.n66 vdd.n63 0.035
R59541 vdd.n275 vdd.n273 0.035
R59542 vdd.n26052 vdd.n26051 0.035
R59543 vdd.n29848 vdd.n29847 0.035
R59544 vdd.n29039 vdd.n29038 0.035
R59545 vdd.n2870 vdd.n2868 0.035
R59546 vdd.n2913 vdd.n2911 0.035
R59547 vdd.n3051 vdd.n3049 0.035
R59548 vdd.n3094 vdd.n3092 0.035
R59549 vdd.n3232 vdd.n3230 0.035
R59550 vdd.n3275 vdd.n3273 0.035
R59551 vdd.n3413 vdd.n3411 0.035
R59552 vdd.n3456 vdd.n3454 0.035
R59553 vdd.n3594 vdd.n3592 0.035
R59554 vdd.n33425 vdd.n33424 0.035
R59555 vdd.n33563 vdd.n33562 0.035
R59556 vdd.n33756 vdd.n33755 0.035
R59557 vdd.n33818 vdd.n33817 0.035
R59558 vdd.n34155 vdd.n34154 0.035
R59559 vdd.n33865 vdd.n33864 0.035
R59560 vdd.n33946 vdd.n33945 0.035
R59561 vdd.n34435 vdd.n34434 0.035
R59562 vdd.n34691 vdd.n34657 0.035
R59563 vdd.n34510 vdd.n34509 0.035
R59564 vdd.n34865 vdd.n34864 0.035
R59565 vdd.n34538 vdd.n34537 0.035
R59566 vdd.n653 vdd.n643 0.035
R59567 vdd.n1027 vdd.n1026 0.035
R59568 vdd.n1039 vdd.n1038 0.035
R59569 vdd.n1125 vdd.n1101 0.035
R59570 vdd.n80 vdd.n79 0.035
R59571 vdd.n287 vdd.n286 0.035
R59572 vdd.n5438 vdd.n5404 0.035
R59573 vdd.n5257 vdd.n5256 0.035
R59574 vdd.n5612 vdd.n5611 0.035
R59575 vdd.n5285 vdd.n5284 0.035
R59576 vdd.n4861 vdd.n4860 0.035
R59577 vdd.n5058 vdd.n5057 0.035
R59578 vdd.n4255 vdd.n4254 0.035
R59579 vdd.n4573 vdd.n4572 0.035
R59580 vdd.n4090 vdd.n4089 0.035
R59581 vdd.n4427 vdd.n4426 0.035
R59582 vdd.n36009 vdd.n36007 0.035
R59583 vdd.n36065 vdd.n36063 0.035
R59584 vdd.n36240 vdd.n36238 0.035
R59585 vdd.n36296 vdd.n36294 0.035
R59586 vdd.n36471 vdd.n36469 0.035
R59587 vdd.n36527 vdd.n36525 0.035
R59588 vdd.n36702 vdd.n36700 0.035
R59589 vdd.n36758 vdd.n36756 0.035
R59590 vdd.n36933 vdd.n36931 0.035
R59591 vdd.n38044 vdd.n38042 0.035
R59592 vdd.n37988 vdd.n37986 0.035
R59593 vdd.n37813 vdd.n37811 0.035
R59594 vdd.n37757 vdd.n37755 0.035
R59595 vdd.n28199 vdd.n28197 0.035
R59596 vdd.n28255 vdd.n28253 0.035
R59597 vdd.n28430 vdd.n28428 0.035
R59598 vdd.n28486 vdd.n28484 0.035
R59599 vdd.n28661 vdd.n28659 0.035
R59600 vdd.n28717 vdd.n28715 0.035
R59601 vdd.n1675 vdd.n1673 0.035
R59602 vdd.n1632 vdd.n1630 0.035
R59603 vdd.n1494 vdd.n1492 0.035
R59604 vdd.n1451 vdd.n1449 0.035
R59605 vdd.n1313 vdd.n1311 0.035
R59606 vdd.n26779 vdd.n26777 0.035
R59607 vdd.n26917 vdd.n26915 0.035
R59608 vdd.n26960 vdd.n26958 0.035
R59609 vdd.n27098 vdd.n27096 0.035
R59610 vdd.n27141 vdd.n27139 0.035
R59611 vdd.n10131 vdd.n10124 0.035
R59612 vdd.n12600 vdd.n10085 0.035
R59613 vdd.n11502 vdd.n11501 0.035
R59614 vdd.n11557 vdd.n11556 0.035
R59615 vdd.n10177 vdd.n10176 0.035
R59616 vdd.n16743 vdd.n16719 0.035
R59617 vdd.n16801 vdd.n16800 0.035
R59618 vdd.n18427 vdd.n18426 0.035
R59619 vdd.n16773 vdd.n16772 0.035
R59620 vdd.n25039 vdd.n25037 0.035
R59621 vdd.n25012 vdd.n25010 0.035
R59622 vdd.n24614 vdd.n24612 0.035
R59623 vdd.n24588 vdd.n24586 0.035
R59624 vdd.n24872 vdd.n24865 0.035
R59625 vdd.n35212 vdd.n35211 0.035
R59626 vdd.n6336 vdd.n6334 0.035
R59627 vdd.n35597 vdd.n35592 0.035
R59628 vdd.n35333 vdd.n35332 0.035
R59629 vdd.n6032 vdd.n6028 0.035
R59630 vdd.n5914 vdd.n5912 0.035
R59631 vdd.n845 vdd.n844 0.035
R59632 vdd.n28055 vdd.n28054 0.035
R59633 vdd.n28805 vdd.n28804 0.035
R59634 vdd.n33549 vdd.n33546 0.035
R59635 vdd.n33586 vdd.n33584 0.035
R59636 vdd.n1022 vdd.n1007 0.035
R59637 vdd.n948 vdd.n947 0.035
R59638 vdd.n25643 vdd.n25642 0.035
R59639 vdd.n25668 vdd.n25666 0.035
R59640 vdd.n27975 vdd.n27974 0.035
R59641 vdd.n25452 vdd.n25449 0.034
R59642 vdd.n25536 vdd.n25532 0.034
R59643 vdd.n33944 vdd.n33888 0.034
R59644 vdd.n35095 vdd.n35046 0.034
R59645 vdd.n34508 vdd.n34459 0.034
R59646 vdd.n221 vdd.n220 0.034
R59647 vdd.n6228 vdd.n6162 0.034
R59648 vdd.n5255 vdd.n5206 0.034
R59649 vdd.n4848 vdd.n4846 0.034
R59650 vdd.n5034 vdd.n5031 0.034
R59651 vdd.n4085 vdd.n4036 0.034
R59652 vdd.n33554 vdd.n33553 0.034
R59653 vdd.n34155 vdd.n34152 0.034
R59654 vdd.n33964 vdd.n33963 0.034
R59655 vdd.n33936 vdd.n33935 0.034
R59656 vdd.n34032 vdd.n34031 0.034
R59657 vdd.n35555 vdd.n35554 0.034
R59658 vdd.n35501 vdd.n35500 0.034
R59659 vdd.n35100 vdd.n35099 0.034
R59660 vdd.n35450 vdd.n35449 0.034
R59661 vdd.n35447 vdd.n35446 0.034
R59662 vdd.n35462 vdd.n35461 0.034
R59663 vdd.n35178 vdd.n35177 0.034
R59664 vdd.n35209 vdd.n35208 0.034
R59665 vdd.n34691 vdd.n34690 0.034
R59666 vdd.n34529 vdd.n34528 0.034
R59667 vdd.n34470 vdd.n34469 0.034
R59668 vdd.n34614 vdd.n34613 0.034
R59669 vdd.n653 vdd.n652 0.034
R59670 vdd.n1024 vdd.n1023 0.034
R59671 vdd.n1135 vdd.n1134 0.034
R59672 vdd.n1125 vdd.n1124 0.034
R59673 vdd.n38 vdd.n37 0.034
R59674 vdd.n5995 vdd.n5994 0.034
R59675 vdd.n6019 vdd.n6018 0.034
R59676 vdd.n6092 vdd.n6091 0.034
R59677 vdd.n6060 vdd.n6059 0.034
R59678 vdd.n6246 vdd.n6245 0.034
R59679 vdd.n6124 vdd.n6123 0.034
R59680 vdd.n6314 vdd.n6309 0.034
R59681 vdd.n6269 vdd.n6268 0.034
R59682 vdd.n5438 vdd.n5437 0.034
R59683 vdd.n5276 vdd.n5275 0.034
R59684 vdd.n5217 vdd.n5216 0.034
R59685 vdd.n5361 vdd.n5360 0.034
R59686 vdd.n4773 vdd.n4772 0.034
R59687 vdd.n5036 vdd.n5035 0.034
R59688 vdd.n4087 vdd.n4086 0.034
R59689 vdd.n4439 vdd.n4438 0.034
R59690 vdd.n25645 vdd.n25644 0.034
R59691 vdd.n25483 vdd.n25482 0.034
R59692 vdd.n11756 vdd.n11683 0.034
R59693 vdd.n11888 vdd.n11796 0.034
R59694 vdd.n22239 vdd.n22231 0.034
R59695 vdd.n22116 vdd.n22115 0.034
R59696 vdd.n21836 vdd.n21835 0.034
R59697 vdd.n21979 vdd.n21887 0.034
R59698 vdd.n27657 vdd.n27643 0.034
R59699 vdd.n26079 vdd.n26064 0.034
R59700 vdd.n27824 vdd.n27823 0.034
R59701 vdd.n10094 vdd.n10068 0.034
R59702 vdd.n25555 vdd.n25553 0.034
R59703 vdd.n25469 vdd.n25467 0.034
R59704 vdd.n28991 vdd.n28977 0.034
R59705 vdd.n10178 vdd.n10135 0.033
R59706 vdd.n10259 vdd.n10258 0.033
R59707 vdd.n16777 vdd.n16776 0.033
R59708 vdd.n16794 vdd.n16793 0.033
R59709 vdd.n29904 vdd.n29892 0.033
R59710 vdd.n33552 vdd.n33512 0.033
R59711 vdd.n1036 vdd.n1035 0.033
R59712 vdd.n33512 vdd.n33511 0.033
R59713 vdd.n1037 vdd.n1036 0.033
R59714 vdd.n1783 vdd.n1771 0.033
R59715 vdd.n34130 vdd.n34127 0.033
R59716 vdd.n34418 vdd.n34379 0.033
R59717 vdd.n35491 vdd.n35487 0.033
R59718 vdd.n35448 vdd.n35445 0.033
R59719 vdd.n35210 vdd.n35207 0.033
R59720 vdd.n34966 vdd.n34962 0.033
R59721 vdd.n34851 vdd.n34848 0.033
R59722 vdd.n5826 vdd.n5825 0.033
R59723 vdd.n6122 vdd.n6093 0.033
R59724 vdd.n6333 vdd.n6270 0.033
R59725 vdd.n5713 vdd.n5709 0.033
R59726 vdd.n5598 vdd.n5595 0.033
R59727 vdd.n4768 vdd.n4724 0.033
R59728 vdd.n4543 vdd.n4536 0.033
R59729 vdd.n4425 vdd.n4422 0.033
R59730 vdd.n4200 vdd.n4137 0.033
R59731 vdd.n3673 vdd.n3658 0.033
R59732 vdd.n33375 vdd.n33373 0.033
R59733 vdd.n33623 vdd.n33622 0.033
R59734 vdd.n33768 vdd.n33767 0.033
R59735 vdd.n33803 vdd.n33802 0.033
R59736 vdd.n33838 vdd.n33835 0.033
R59737 vdd.n34143 vdd.n34142 0.033
R59738 vdd.n34436 vdd.n34365 0.033
R59739 vdd.n34400 vdd.n34399 0.033
R59740 vdd.n34000 vdd.n33999 0.033
R59741 vdd.n35162 vdd.n35161 0.033
R59742 vdd.n35098 vdd.n35032 0.033
R59743 vdd.n35414 vdd.n35413 0.033
R59744 vdd.n35458 vdd.n35381 0.033
R59745 vdd.n35097 vdd.n35096 0.033
R59746 vdd.n35454 vdd.n35453 0.033
R59747 vdd.n34678 vdd.n34677 0.033
R59748 vdd.n34869 vdd.n34791 0.033
R59749 vdd.n34818 vdd.n34817 0.033
R59750 vdd.n34582 vdd.n34581 0.033
R59751 vdd.n689 vdd.n595 0.033
R59752 vdd.n981 vdd.n980 0.033
R59753 vdd.n1099 vdd.n1098 0.033
R59754 vdd.n942 vdd.n941 0.033
R59755 vdd.n827 vdd.n826 0.033
R59756 vdd.n585 vdd.n583 0.033
R59757 vdd.n13 vdd.n8 0.033
R59758 vdd.n24 vdd.n21 0.033
R59759 vdd.n401 vdd.n398 0.033
R59760 vdd.n77 vdd.n76 0.033
R59761 vdd.n288 vdd.n256 0.033
R59762 vdd.n114 vdd.n111 0.033
R59763 vdd.n284 vdd.n283 0.033
R59764 vdd.n343 vdd.n342 0.033
R59765 vdd.n6293 vdd.n6292 0.033
R59766 vdd.n6244 vdd.n6161 0.033
R59767 vdd.n6209 vdd.n6208 0.033
R59768 vdd.n6131 vdd.n6071 0.033
R59769 vdd.n6230 vdd.n6229 0.033
R59770 vdd.n6130 vdd.n6129 0.033
R59771 vdd.n5425 vdd.n5424 0.033
R59772 vdd.n5616 vdd.n5538 0.033
R59773 vdd.n5565 vdd.n5564 0.033
R59774 vdd.n5329 vdd.n5328 0.033
R59775 vdd.n5120 vdd.n5119 0.033
R59776 vdd.n4862 vdd.n4827 0.033
R59777 vdd.n5127 vdd.n5126 0.033
R59778 vdd.n4858 vdd.n4857 0.033
R59779 vdd.n4787 vdd.n4784 0.033
R59780 vdd.n5048 vdd.n4972 0.033
R59781 vdd.n5018 vdd.n5017 0.033
R59782 vdd.n5056 vdd.n5055 0.033
R59783 vdd.n4515 vdd.n4514 0.033
R59784 vdd.n4443 vdd.n4365 0.033
R59785 vdd.n4391 vdd.n4390 0.033
R59786 vdd.n4424 vdd.n4423 0.033
R59787 vdd.n4447 vdd.n4446 0.033
R59788 vdd.n4160 vdd.n4159 0.033
R59789 vdd.n4181 vdd.n4175 0.033
R59790 vdd.n4136 vdd.n4135 0.033
R59791 vdd.n25403 vdd.n25399 0.033
R59792 vdd.n25574 vdd.n25573 0.033
R59793 vdd.n25588 vdd.n25587 0.033
R59794 vdd.n25545 vdd.n25544 0.033
R59795 vdd.n32210 vdd.n32209 0.033
R59796 vdd.n24555 vdd.n24554 0.033
R59797 vdd.n33844 vdd.n33842 0.033
R59798 vdd.n25570 vdd.n25569 0.033
R59799 vdd.n25587 vdd.n25585 0.033
R59800 vdd.n34013 vdd.n34012 0.033
R59801 vdd.n34601 vdd.n34600 0.033
R59802 vdd.n5348 vdd.n5347 0.033
R59803 vdd.n4659 vdd.n4658 0.033
R59804 vdd.n25517 vdd.n25516 0.033
R59805 vdd.n30249 vdd.n30248 0.032
R59806 vdd.n29750 vdd.n29749 0.032
R59807 vdd.n30699 vdd.n30698 0.032
R59808 vdd.n25616 vdd.n25615 0.032
R59809 vdd.n4179 vdd.n4178 0.032
R59810 vdd.n29037 vdd.n29036 0.032
R59811 vdd.n2774 vdd.n2772 0.032
R59812 vdd.n2833 vdd.n2826 0.032
R59813 vdd.n2955 vdd.n2953 0.032
R59814 vdd.n3014 vdd.n3007 0.032
R59815 vdd.n3136 vdd.n3134 0.032
R59816 vdd.n3195 vdd.n3188 0.032
R59817 vdd.n3317 vdd.n3315 0.032
R59818 vdd.n3376 vdd.n3369 0.032
R59819 vdd.n3498 vdd.n3496 0.032
R59820 vdd.n3557 vdd.n3550 0.032
R59821 vdd.n33297 vdd.n33294 0.032
R59822 vdd.n33551 vdd.n33550 0.032
R59823 vdd.n33650 vdd.n33649 0.032
R59824 vdd.n33615 vdd.n33608 0.032
R59825 vdd.n33762 vdd.n33761 0.032
R59826 vdd.n34140 vdd.n34139 0.032
R59827 vdd.n34129 vdd.n34128 0.032
R59828 vdd.n34378 vdd.n34377 0.032
R59829 vdd.n34354 vdd.n34353 0.032
R59830 vdd.n34016 vdd.n34014 0.032
R59831 vdd.n34046 vdd.n34045 0.032
R59832 vdd.n35590 vdd.n35589 0.032
R59833 vdd.n35094 vdd.n35093 0.032
R59834 vdd.n34941 vdd.n34940 0.032
R59835 vdd.n34684 vdd.n34683 0.032
R59836 vdd.n34850 vdd.n34849 0.032
R59837 vdd.n34873 vdd.n34872 0.032
R59838 vdd.n34603 vdd.n34597 0.032
R59839 vdd.n34559 vdd.n34558 0.032
R59840 vdd.n1042 vdd.n1041 0.032
R59841 vdd.n910 vdd.n907 0.032
R59842 vdd.n930 vdd.n929 0.032
R59843 vdd.n293 vdd.n292 0.032
R59844 vdd.n5929 vdd.n5928 0.032
R59845 vdd.n6164 vdd.n6163 0.032
R59846 vdd.n5688 vdd.n5687 0.032
R59847 vdd.n5431 vdd.n5430 0.032
R59848 vdd.n5597 vdd.n5596 0.032
R59849 vdd.n5620 vdd.n5619 0.032
R59850 vdd.n5350 vdd.n5344 0.032
R59851 vdd.n5306 vdd.n5305 0.032
R59852 vdd.n5163 vdd.n5162 0.032
R59853 vdd.n5099 vdd.n5098 0.032
R59854 vdd.n4867 vdd.n4866 0.032
R59855 vdd.n4871 vdd.n4809 0.032
R59856 vdd.n4798 vdd.n4797 0.032
R59857 vdd.n4767 vdd.n4766 0.032
R59858 vdd.n4880 vdd.n4879 0.032
R59859 vdd.n4460 vdd.n4459 0.032
R59860 vdd.n4265 vdd.n4264 0.032
R59861 vdd.n4106 vdd.n4105 0.032
R59862 vdd.n4047 vdd.n4046 0.032
R59863 vdd.n4084 vdd.n4083 0.032
R59864 vdd.n4192 vdd.n4191 0.032
R59865 vdd.n35888 vdd.n35886 0.032
R59866 vdd.n35963 vdd.n35953 0.032
R59867 vdd.n36119 vdd.n36117 0.032
R59868 vdd.n36194 vdd.n36184 0.032
R59869 vdd.n36350 vdd.n36348 0.032
R59870 vdd.n36425 vdd.n36415 0.032
R59871 vdd.n36581 vdd.n36579 0.032
R59872 vdd.n36656 vdd.n36646 0.032
R59873 vdd.n36812 vdd.n36810 0.032
R59874 vdd.n36887 vdd.n36877 0.032
R59875 vdd.n38098 vdd.n38096 0.032
R59876 vdd.n37942 vdd.n37932 0.032
R59877 vdd.n37867 vdd.n37865 0.032
R59878 vdd.n37711 vdd.n37701 0.032
R59879 vdd.n37636 vdd.n37634 0.032
R59880 vdd.n28309 vdd.n28307 0.032
R59881 vdd.n28384 vdd.n28374 0.032
R59882 vdd.n28540 vdd.n28538 0.032
R59883 vdd.n28615 vdd.n28605 0.032
R59884 vdd.n28771 vdd.n28769 0.032
R59885 vdd.n1717 vdd.n1715 0.032
R59886 vdd.n1595 vdd.n1588 0.032
R59887 vdd.n1536 vdd.n1534 0.032
R59888 vdd.n1414 vdd.n1407 0.032
R59889 vdd.n1355 vdd.n1353 0.032
R59890 vdd.n26821 vdd.n26819 0.032
R59891 vdd.n26880 vdd.n26873 0.032
R59892 vdd.n27002 vdd.n27000 0.032
R59893 vdd.n27061 vdd.n27054 0.032
R59894 vdd.n27183 vdd.n27181 0.032
R59895 vdd.n25612 vdd.n25609 0.032
R59896 vdd.n25526 vdd.n25525 0.032
R59897 vdd.n25485 vdd.n25484 0.032
R59898 vdd.n10253 vdd.n10125 0.032
R59899 vdd.n11775 vdd.n11665 0.032
R59900 vdd.n11748 vdd.n11747 0.032
R59901 vdd.n11875 vdd.n11805 0.032
R59902 vdd.n11887 vdd.n11801 0.032
R59903 vdd.n11907 vdd.n11787 0.032
R59904 vdd.n22242 vdd.n22241 0.032
R59905 vdd.n15060 vdd.n15059 0.032
R59906 vdd.n21867 vdd.n21866 0.032
R59907 vdd.n21830 vdd.n21829 0.032
R59908 vdd.n21966 vdd.n21896 0.032
R59909 vdd.n21978 vdd.n21892 0.032
R59910 vdd.n21751 vdd.n21750 0.032
R59911 vdd.n25601 vdd.n25600 0.032
R59912 vdd.n25659 vdd.n25658 0.032
R59913 vdd.n29839 vdd.n29829 0.032
R59914 vdd.n33402 vdd.n33401 0.032
R59915 vdd.n33525 vdd.n33524 0.032
R59916 vdd.n33603 vdd.n33602 0.032
R59917 vdd.n723 vdd.n722 0.032
R59918 vdd.n1114 vdd.n1113 0.032
R59919 vdd.n434 vdd.n433 0.032
R59920 vdd.n152 vdd.n151 0.032
R59921 vdd.n346 vdd.n345 0.032
R59922 vdd.n29873 vdd.n29863 0.032
R59923 vdd.n29039 vdd.n29017 0.032
R59924 vdd.n29949 vdd.n29948 0.031
R59925 vdd.n28892 vdd.n28105 0.031
R59926 vdd.n25666 vdd.n25663 0.031
R59927 vdd.n25642 vdd.n25641 0.031
R59928 vdd.n35043 vdd.n35042 0.031
R59929 vdd.n6244 vdd.n6241 0.031
R59930 vdd.n35098 vdd.n35043 0.031
R59931 vdd.n6241 vdd.n6240 0.031
R59932 vdd.n35176 vdd.n35175 0.031
R59933 vdd.n6313 vdd.n6312 0.031
R59934 vdd.n30686 vdd.n30684 0.031
R59935 vdd.n27894 vdd.n27892 0.031
R59936 vdd.n11917 vdd.n11916 0.031
R59937 vdd.n22003 vdd.n22002 0.031
R59938 vdd.n25553 vdd.n25549 0.031
R59939 vdd.n25467 vdd.n25463 0.031
R59940 vdd.n33560 vdd.n33559 0.031
R59941 vdd.n33753 vdd.n33752 0.031
R59942 vdd.n34126 vdd.n34125 0.031
R59943 vdd.n34183 vdd.n34182 0.031
R59944 vdd.n34410 vdd.n34409 0.031
R59945 vdd.n34417 vdd.n34416 0.031
R59946 vdd.n34438 vdd.n34437 0.031
R59947 vdd.n34016 vdd.n34013 0.031
R59948 vdd.n34044 vdd.n34043 0.031
R59949 vdd.n35275 vdd.n35274 0.031
R59950 vdd.n35527 vdd.n35526 0.031
R59951 vdd.n35271 vdd.n35270 0.031
R59952 vdd.n35116 vdd.n35115 0.031
R59953 vdd.n35057 vdd.n35056 0.031
R59954 vdd.n35194 vdd.n35193 0.031
R59955 vdd.n35282 vdd.n35281 0.031
R59956 vdd.n34968 vdd.n34967 0.031
R59957 vdd.n34742 vdd.n34741 0.031
R59958 vdd.n34835 vdd.n34834 0.031
R59959 vdd.n34847 vdd.n34846 0.031
R59960 vdd.n34871 vdd.n34870 0.031
R59961 vdd.n34603 vdd.n34601 0.031
R59962 vdd.n34621 vdd.n34620 0.031
R59963 vdd.n664 vdd.n663 0.031
R59964 vdd.n910 vdd.n909 0.031
R59965 vdd.n68 vdd.n67 0.031
R59966 vdd.n6009 vdd.n5976 0.031
R59967 vdd.n5794 vdd.n5793 0.031
R59968 vdd.n5841 vdd.n5838 0.031
R59969 vdd.n6249 vdd.n6248 0.031
R59970 vdd.n6220 vdd.n6219 0.031
R59971 vdd.n6325 vdd.n6324 0.031
R59972 vdd.n5910 vdd.n5909 0.031
R59973 vdd.n5715 vdd.n5714 0.031
R59974 vdd.n5489 vdd.n5488 0.031
R59975 vdd.n5582 vdd.n5581 0.031
R59976 vdd.n5594 vdd.n5593 0.031
R59977 vdd.n5618 vdd.n5617 0.031
R59978 vdd.n5350 vdd.n5348 0.031
R59979 vdd.n5368 vdd.n5367 0.031
R59980 vdd.n5033 vdd.n5032 0.031
R59981 vdd.n4690 vdd.n4689 0.031
R59982 vdd.n4258 vdd.n4257 0.031
R59983 vdd.n27600 vdd.n27597 0.031
R59984 vdd.n27466 vdd.n27465 0.031
R59985 vdd.n26016 vdd.n26013 0.031
R59986 vdd.n25912 vdd.n25911 0.031
R59987 vdd.n30748 vdd.n30747 0.031
R59988 vdd.n32582 vdd.n32579 0.031
R59989 vdd.n31197 vdd.n31194 0.031
R59990 vdd.n2142 vdd.n2141 0.031
R59991 vdd.n2534 vdd.n2533 0.031
R59992 vdd.n2315 vdd.n2119 0.031
R59993 vdd.n11902 vdd.n11788 0.031
R59994 vdd.n21993 vdd.n21879 0.031
R59995 vdd.n25631 vdd.n25627 0.031
R59996 vdd.n25561 vdd.n25560 0.031
R59997 vdd.n27638 vdd.n27637 0.031
R59998 vdd.n27359 vdd.n27358 0.031
R59999 vdd.n27510 vdd.n27509 0.031
R60000 vdd.n25811 vdd.n25810 0.031
R60001 vdd.n26059 vdd.n26058 0.03
R60002 vdd.n33704 vdd.n33703 0.03
R60003 vdd.n795 vdd.n794 0.03
R60004 vdd.n25947 vdd.n25946 0.03
R60005 vdd.n33439 vdd.n33438 0.03
R60006 vdd.n33548 vdd.n33547 0.03
R60007 vdd.n33569 vdd.n33568 0.03
R60008 vdd.n33593 vdd.n33592 0.03
R60009 vdd.n34324 vdd.n34323 0.03
R60010 vdd.n33890 vdd.n33889 0.03
R60011 vdd.n35262 vdd.n35261 0.03
R60012 vdd.n34886 vdd.n34885 0.03
R60013 vdd.n34507 vdd.n34506 0.03
R60014 vdd.n893 vdd.n892 0.03
R60015 vdd.n550 vdd.n549 0.03
R60016 vdd.n149 vdd.n148 0.03
R60017 vdd.n290 vdd.n289 0.03
R60018 vdd.n5832 vdd.n5831 0.03
R60019 vdd.n5633 vdd.n5632 0.03
R60020 vdd.n5254 vdd.n5253 0.03
R60021 vdd.n5153 vdd.n5152 0.03
R60022 vdd.n5099 vdd.n5090 0.03
R60023 vdd.n4864 vdd.n4863 0.03
R60024 vdd.n4871 vdd.n4870 0.03
R60025 vdd.n4789 vdd.n4788 0.03
R60026 vdd.n4757 vdd.n4756 0.03
R60027 vdd.n4734 vdd.n4733 0.03
R60028 vdd.n4924 vdd.n4923 0.03
R60029 vdd.n4563 vdd.n4507 0.03
R60030 vdd.n4243 vdd.n4242 0.03
R60031 vdd.n4272 vdd.n4271 0.03
R60032 vdd.n27594 vdd.n27592 0.03
R60033 vdd.n27464 vdd.n27463 0.03
R60034 vdd.n26010 vdd.n26008 0.03
R60035 vdd.n25910 vdd.n25909 0.03
R60036 vdd.n25519 vdd.n25518 0.03
R60037 vdd.n10251 vdd.n10250 0.03
R60038 vdd.n10129 vdd.n10124 0.03
R60039 vdd.n11783 vdd.n11779 0.03
R60040 vdd.n22362 vdd.n22350 0.03
R60041 vdd.n22091 vdd.n22079 0.03
R60042 vdd.n16603 vdd.n16602 0.03
R60043 vdd.n21875 vdd.n21872 0.03
R60044 vdd.n30995 vdd.n30991 0.03
R60045 vdd.n27756 vdd.n27755 0.03
R60046 vdd.n2450 vdd.n2449 0.03
R60047 vdd.n27410 vdd.n27409 0.029
R60048 vdd.n25518 vdd.n25517 0.029
R60049 vdd.n27853 vdd.n27852 0.029
R60050 vdd.n28098 vdd.n28097 0.029
R60051 vdd.n2859 vdd.n2857 0.029
R60052 vdd.n2924 vdd.n2922 0.029
R60053 vdd.n3040 vdd.n3038 0.029
R60054 vdd.n3105 vdd.n3103 0.029
R60055 vdd.n3221 vdd.n3219 0.029
R60056 vdd.n3286 vdd.n3284 0.029
R60057 vdd.n3402 vdd.n3400 0.029
R60058 vdd.n3467 vdd.n3465 0.029
R60059 vdd.n3583 vdd.n3581 0.029
R60060 vdd.n33471 vdd.n33470 0.029
R60061 vdd.n33490 vdd.n33485 0.029
R60062 vdd.n33501 vdd.n33497 0.029
R60063 vdd.n33558 vdd.n33503 0.029
R60064 vdd.n33552 vdd.n33515 0.029
R60065 vdd.n33518 vdd.n33517 0.029
R60066 vdd.n33297 vdd.n33295 0.029
R60067 vdd.n33326 vdd.n33325 0.029
R60068 vdd.n33751 vdd.n33746 0.029
R60069 vdd.n33615 vdd.n33612 0.029
R60070 vdd.n33656 vdd.n33653 0.029
R60071 vdd.n33665 vdd.n33664 0.029
R60072 vdd.n33768 vdd.n33765 0.029
R60073 vdd.n33812 vdd.n33809 0.029
R60074 vdd.n34099 vdd.n34098 0.029
R60075 vdd.n34138 vdd.n34108 0.029
R60076 vdd.n34281 vdd.n34280 0.029
R60077 vdd.n34307 vdd.n34304 0.029
R60078 vdd.n34314 vdd.n34313 0.029
R60079 vdd.n34176 vdd.n34173 0.029
R60080 vdd.n34200 vdd.n34199 0.029
R60081 vdd.n33923 vdd.n33922 0.029
R60082 vdd.n33893 vdd.n33892 0.029
R60083 vdd.n33943 vdd.n33942 0.029
R60084 vdd.n33977 vdd.n33976 0.029
R60085 vdd.n35573 vdd.n35570 0.029
R60086 vdd.n35547 vdd.n35546 0.029
R60087 vdd.n35475 vdd.n35473 0.029
R60088 vdd.n35260 vdd.n35259 0.029
R60089 vdd.n35493 vdd.n35492 0.029
R60090 vdd.n35087 vdd.n35086 0.029
R60091 vdd.n35431 vdd.n35430 0.029
R60092 vdd.n35444 vdd.n35443 0.029
R60093 vdd.n35460 vdd.n35459 0.029
R60094 vdd.n35139 vdd.n35138 0.029
R60095 vdd.n35178 vdd.n35176 0.029
R60096 vdd.n35206 vdd.n35205 0.029
R60097 vdd.n35284 vdd.n35283 0.029
R60098 vdd.n35326 vdd.n35325 0.029
R60099 vdd.n35321 vdd.n35318 0.029
R60100 vdd.n34676 vdd.n34675 0.029
R60101 vdd.n34682 vdd.n34680 0.029
R60102 vdd.n34917 vdd.n34916 0.029
R60103 vdd.n34902 vdd.n34899 0.029
R60104 vdd.n35003 vdd.n35002 0.029
R60105 vdd.n34726 vdd.n34723 0.029
R60106 vdd.n34700 vdd.n34699 0.029
R60107 vdd.n34500 vdd.n34499 0.029
R60108 vdd.n34497 vdd.n34496 0.029
R60109 vdd.n34552 vdd.n34551 0.029
R60110 vdd.n711 vdd.n710 0.029
R60111 vdd.n977 vdd.n972 0.029
R60112 vdd.n991 vdd.n987 0.029
R60113 vdd.n1040 vdd.n993 0.029
R60114 vdd.n1037 vdd.n1025 0.029
R60115 vdd.n999 vdd.n998 0.029
R60116 vdd.n653 vdd.n648 0.029
R60117 vdd.n1125 vdd.n1105 0.029
R60118 vdd.n1072 vdd.n1069 0.029
R60119 vdd.n1058 vdd.n1057 0.029
R60120 vdd.n898 vdd.n897 0.029
R60121 vdd.n820 vdd.n817 0.029
R60122 vdd.n485 vdd.n484 0.029
R60123 vdd.n15 vdd.n14 0.029
R60124 vdd.n452 vdd.n451 0.029
R60125 vdd.n85 vdd.n84 0.029
R60126 vdd.n266 vdd.n265 0.029
R60127 vdd.n122 vdd.n121 0.029
R60128 vdd.n155 vdd.n152 0.029
R60129 vdd.n172 vdd.n171 0.029
R60130 vdd.n298 vdd.n236 0.029
R60131 vdd.n328 vdd.n327 0.029
R60132 vdd.n337 vdd.n334 0.029
R60133 vdd.n365 vdd.n359 0.029
R60134 vdd.n5945 vdd.n5942 0.029
R60135 vdd.n5960 vdd.n5959 0.029
R60136 vdd.n5830 vdd.n5816 0.029
R60137 vdd.n5804 vdd.n5803 0.029
R60138 vdd.n6002 vdd.n6001 0.029
R60139 vdd.n6167 vdd.n6166 0.029
R60140 vdd.n6197 vdd.n6196 0.029
R60141 vdd.n6114 vdd.n6113 0.029
R60142 vdd.n6121 vdd.n6120 0.029
R60143 vdd.n6133 vdd.n6132 0.029
R60144 vdd.n6262 vdd.n6261 0.029
R60145 vdd.n6314 vdd.n6313 0.029
R60146 vdd.n6332 vdd.n6331 0.029
R60147 vdd.n5901 vdd.n5900 0.029
R60148 vdd.n5884 vdd.n5883 0.029
R60149 vdd.n5879 vdd.n5876 0.029
R60150 vdd.n5423 vdd.n5422 0.029
R60151 vdd.n5429 vdd.n5427 0.029
R60152 vdd.n5664 vdd.n5663 0.029
R60153 vdd.n5649 vdd.n5646 0.029
R60154 vdd.n5750 vdd.n5749 0.029
R60155 vdd.n5473 vdd.n5470 0.029
R60156 vdd.n5447 vdd.n5446 0.029
R60157 vdd.n5247 vdd.n5246 0.029
R60158 vdd.n5244 vdd.n5243 0.029
R60159 vdd.n5299 vdd.n5298 0.029
R60160 vdd.n4644 vdd.n4643 0.029
R60161 vdd.n4633 vdd.n4630 0.029
R60162 vdd.n5156 vdd.n5155 0.029
R60163 vdd.n4845 vdd.n4844 0.029
R60164 vdd.n4733 vdd.n4727 0.029
R60165 vdd.n4998 vdd.n4997 0.029
R60166 vdd.n4975 vdd.n4974 0.029
R60167 vdd.n5030 vdd.n5029 0.029
R60168 vdd.n4688 vdd.n4687 0.029
R60169 vdd.n4661 vdd.n4660 0.029
R60170 vdd.n4898 vdd.n4896 0.029
R60171 vdd.n4915 vdd.n4912 0.029
R60172 vdd.n4253 vdd.n4252 0.029
R60173 vdd.n4539 vdd.n4537 0.029
R60174 vdd.n4491 vdd.n4490 0.029
R60175 vdd.n4476 vdd.n4473 0.029
R60176 vdd.n4545 vdd.n4544 0.029
R60177 vdd.n4300 vdd.n4297 0.029
R60178 vdd.n4274 vdd.n4273 0.029
R60179 vdd.n4316 vdd.n4315 0.029
R60180 vdd.n4077 vdd.n4076 0.029
R60181 vdd.n4408 vdd.n4407 0.029
R60182 vdd.n4421 vdd.n4420 0.029
R60183 vdd.n4445 vdd.n4444 0.029
R60184 vdd.n4129 vdd.n4128 0.029
R60185 vdd.n4181 vdd.n4179 0.029
R60186 vdd.n4199 vdd.n4198 0.029
R60187 vdd.n35995 vdd.n35993 0.029
R60188 vdd.n36079 vdd.n36077 0.029
R60189 vdd.n36226 vdd.n36224 0.029
R60190 vdd.n36310 vdd.n36308 0.029
R60191 vdd.n36457 vdd.n36455 0.029
R60192 vdd.n36541 vdd.n36539 0.029
R60193 vdd.n36688 vdd.n36686 0.029
R60194 vdd.n36772 vdd.n36770 0.029
R60195 vdd.n36919 vdd.n36917 0.029
R60196 vdd.n38058 vdd.n38056 0.029
R60197 vdd.n37974 vdd.n37972 0.029
R60198 vdd.n37827 vdd.n37825 0.029
R60199 vdd.n37743 vdd.n37741 0.029
R60200 vdd.n28185 vdd.n28183 0.029
R60201 vdd.n28269 vdd.n28267 0.029
R60202 vdd.n28416 vdd.n28414 0.029
R60203 vdd.n28500 vdd.n28498 0.029
R60204 vdd.n28647 vdd.n28645 0.029
R60205 vdd.n28731 vdd.n28729 0.029
R60206 vdd.n1686 vdd.n1684 0.029
R60207 vdd.n1621 vdd.n1619 0.029
R60208 vdd.n1505 vdd.n1503 0.029
R60209 vdd.n1440 vdd.n1438 0.029
R60210 vdd.n1324 vdd.n1322 0.029
R60211 vdd.n26790 vdd.n26788 0.029
R60212 vdd.n26906 vdd.n26904 0.029
R60213 vdd.n26971 vdd.n26969 0.029
R60214 vdd.n27087 vdd.n27085 0.029
R60215 vdd.n27152 vdd.n27150 0.029
R60216 vdd.n27609 vdd.n27608 0.029
R60217 vdd.n27550 vdd.n27549 0.029
R60218 vdd.n27441 vdd.n27438 0.029
R60219 vdd.n27318 vdd.n27315 0.029
R60220 vdd.n27336 vdd.n27335 0.029
R60221 vdd.n26030 vdd.n26029 0.029
R60222 vdd.n25987 vdd.n25986 0.029
R60223 vdd.n25887 vdd.n25884 0.029
R60224 vdd.n25770 vdd.n25767 0.029
R60225 vdd.n25788 vdd.n25787 0.029
R60226 vdd.n30902 vdd.n30901 0.029
R60227 vdd.n29598 vdd.n29597 0.029
R60228 vdd.n27691 vdd.n27690 0.029
R60229 vdd.n22339 vdd.n22331 0.029
R60230 vdd.n25047 vdd.n25046 0.029
R60231 vdd.n25046 vdd.n25044 0.029
R60232 vdd.n25005 vdd.n25003 0.029
R60233 vdd.n24581 vdd.n24579 0.029
R60234 vdd.n25856 vdd.n25855 0.029
R60235 vdd.n1819 vdd.n1817 0.029
R60236 vdd.n28130 vdd.n28129 0.028
R60237 vdd.n33349 vdd.n33348 0.028
R60238 vdd.n33759 vdd.n33758 0.028
R60239 vdd.n34301 vdd.n34300 0.028
R60240 vdd.n34261 vdd.n34252 0.028
R60241 vdd.n34146 vdd.n34145 0.028
R60242 vdd.n34261 vdd.n34260 0.028
R60243 vdd.n34149 vdd.n34148 0.028
R60244 vdd.n34198 vdd.n34197 0.028
R60245 vdd.n34209 vdd.n34208 0.028
R60246 vdd.n34986 vdd.n34933 0.028
R60247 vdd.n34666 vdd.n34665 0.028
R60248 vdd.n34999 vdd.n34998 0.028
R60249 vdd.n34986 vdd.n34985 0.028
R60250 vdd.n34687 vdd.n34686 0.028
R60251 vdd.n34698 vdd.n34697 0.028
R60252 vdd.n34746 vdd.n34745 0.028
R60253 vdd.n721 vdd.n720 0.028
R60254 vdd.n753 vdd.n752 0.028
R60255 vdd.n757 vdd.n756 0.028
R60256 vdd.n1006 vdd.n1005 0.028
R60257 vdd.n1046 vdd.n970 0.028
R60258 vdd.n1021 vdd.n1020 0.028
R60259 vdd.n1046 vdd.n1045 0.028
R60260 vdd.n1116 vdd.n1115 0.028
R60261 vdd.n1118 vdd.n1117 0.028
R60262 vdd.n807 vdd.n804 0.028
R60263 vdd.n807 vdd.n805 0.028
R60264 vdd.n559 vdd.n558 0.028
R60265 vdd.n65 vdd.n64 0.028
R60266 vdd.n105 vdd.n104 0.028
R60267 vdd.n5733 vdd.n5680 0.028
R60268 vdd.n5413 vdd.n5412 0.028
R60269 vdd.n5746 vdd.n5745 0.028
R60270 vdd.n5733 vdd.n5732 0.028
R60271 vdd.n5434 vdd.n5433 0.028
R60272 vdd.n5445 vdd.n5444 0.028
R60273 vdd.n5493 vdd.n5492 0.028
R60274 vdd.n4580 vdd.n4579 0.028
R60275 vdd.n4074 vdd.n4073 0.028
R60276 vdd.n27352 vdd.n27351 0.028
R60277 vdd.n25804 vdd.n25803 0.028
R60278 vdd.n30878 vdd.n30875 0.028
R60279 vdd.n13741 ldomc_0.otaldom_0.pdiffm_0.vdd 0.028
R60280 ldomc_0.otaldom_0.pmosbm_0.vdd vdd.n14974 0.028
R60281 vdd.n22030 vdd.n22029 0.028
R60282 vdd.n22033 vdd.n22032 0.028
R60283 vdd.n24387 vdd.n24386 0.028
R60284 vdd.n24390 vdd.n24389 0.028
R60285 bandgapmd_0.otam_1.pdiffm_0.vdd vdd.n21092 0.028
R60286 vdd.n20026 bandgapmd_0.otam_1.pmosbm_0.vdd 0.028
R60287 vdd.n24892 vdd.n24891 0.028
R60288 vdd.n24749 vdd.n24745 0.028
R60289 vdd.n24750 vdd.n24749 0.028
R60290 vdd.n25166 vdd.n25165 0.028
R60291 vdd.n25165 vdd.n25161 0.028
R60292 vdd.n10180 vdd.n10179 0.028
R60293 vdd.n16775 vdd.n16774 0.028
R60294 vdd.n13138 vdd.n13137 0.028
R60295 vdd.n21688 vdd.n21687 0.028
R60296 vdd.n25473 vdd.n25472 0.028
R60297 vdd.n29953 vdd.n29849 0.027
R60298 vdd.n25557 vdd.n25556 0.027
R60299 vdd.n11680 vdd.n11679 0.027
R60300 vdd.n21762 vdd.n21758 0.027
R60301 vdd.n2763 vdd.n2761 0.027
R60302 vdd.n2844 vdd.n2837 0.027
R60303 vdd.n2944 vdd.n2942 0.027
R60304 vdd.n3025 vdd.n3018 0.027
R60305 vdd.n3125 vdd.n3123 0.027
R60306 vdd.n3206 vdd.n3199 0.027
R60307 vdd.n3306 vdd.n3304 0.027
R60308 vdd.n3387 vdd.n3380 0.027
R60309 vdd.n3487 vdd.n3485 0.027
R60310 vdd.n3568 vdd.n3561 0.027
R60311 vdd.n33568 vdd.n33567 0.027
R60312 vdd.n33673 vdd.n33672 0.027
R60313 vdd.n33606 vdd.n33605 0.027
R60314 vdd.n35580 vdd.n35579 0.027
R60315 vdd.n35515 vdd.n35514 0.027
R60316 vdd.n35272 vdd.n35271 0.027
R60317 vdd.n35084 vdd.n35083 0.027
R60318 vdd.n35441 vdd.n35440 0.027
R60319 vdd.n35203 vdd.n35202 0.027
R60320 vdd.n605 vdd.n604 0.027
R60321 vdd.n442 vdd.n441 0.027
R60322 vdd.n431 vdd.n430 0.027
R60323 vdd.n83 vdd.n82 0.027
R60324 vdd.n162 vdd.n161 0.027
R60325 vdd.n298 vdd.n296 0.027
R60326 vdd.n5984 vdd.n5983 0.027
R60327 vdd.n5836 vdd.n5794 0.027
R60328 vdd.n6026 vdd.n6025 0.027
R60329 vdd.n6103 vdd.n6102 0.027
R60330 vdd.n6227 vdd.n6226 0.027
R60331 vdd.n6281 vdd.n6280 0.027
R60332 vdd.n4661 vdd.n4659 0.027
R60333 vdd.n4681 vdd.n4680 0.027
R60334 vdd.n4920 vdd.n4919 0.027
R60335 vdd.n4559 vdd.n4558 0.027
R60336 vdd.n4262 vdd.n4243 0.027
R60337 vdd.n4418 vdd.n4417 0.027
R60338 vdd.n4148 vdd.n4147 0.027
R60339 vdd.n35874 vdd.n35872 0.027
R60340 vdd.n35977 vdd.n35967 0.027
R60341 vdd.n36105 vdd.n36103 0.027
R60342 vdd.n36208 vdd.n36198 0.027
R60343 vdd.n36336 vdd.n36334 0.027
R60344 vdd.n36439 vdd.n36429 0.027
R60345 vdd.n36567 vdd.n36565 0.027
R60346 vdd.n36670 vdd.n36660 0.027
R60347 vdd.n36798 vdd.n36796 0.027
R60348 vdd.n36901 vdd.n36891 0.027
R60349 vdd.n38084 vdd.n38082 0.027
R60350 vdd.n37956 vdd.n37946 0.027
R60351 vdd.n37853 vdd.n37851 0.027
R60352 vdd.n37725 vdd.n37715 0.027
R60353 vdd.n37622 vdd.n37620 0.027
R60354 vdd.n28295 vdd.n28293 0.027
R60355 vdd.n28398 vdd.n28388 0.027
R60356 vdd.n28526 vdd.n28524 0.027
R60357 vdd.n28629 vdd.n28619 0.027
R60358 vdd.n28757 vdd.n28755 0.027
R60359 vdd.n1706 vdd.n1704 0.027
R60360 vdd.n1606 vdd.n1599 0.027
R60361 vdd.n1525 vdd.n1523 0.027
R60362 vdd.n1425 vdd.n1418 0.027
R60363 vdd.n1344 vdd.n1342 0.027
R60364 vdd.n26810 vdd.n26808 0.027
R60365 vdd.n26891 vdd.n26884 0.027
R60366 vdd.n26991 vdd.n26989 0.027
R60367 vdd.n27072 vdd.n27065 0.027
R60368 vdd.n27172 vdd.n27170 0.027
R60369 vdd.n11677 vdd.n11669 0.027
R60370 vdd.n21856 vdd.n21847 0.027
R60371 vdd.n24970 vdd.n24956 0.027
R60372 vdd.n24901 vdd.n24900 0.027
R60373 vdd.n24920 vdd.n24919 0.027
R60374 vdd.n24681 vdd.n24673 0.027
R60375 vdd.n25099 vdd.n25091 0.027
R60376 vdd.n10198 vdd.n10197 0.027
R60377 vdd.n10203 vdd.n10198 0.027
R60378 vdd.n10205 vdd.n10204 0.027
R60379 vdd.n16779 vdd.n16778 0.027
R60380 vdd.n16780 vdd.n16779 0.027
R60381 vdd.n16782 vdd.n16781 0.027
R60382 vdd.n31935 vdd.n31934 0.027
R60383 vdd.n27516 vdd.n27515 0.026
R60384 vdd.n33329 vdd.n33328 0.026
R60385 vdd.n33653 vdd.n33652 0.026
R60386 vdd.n33821 vdd.n33820 0.026
R60387 vdd.n618 vdd.n617 0.026
R60388 vdd.n1069 vdd.n1068 0.026
R60389 vdd.n842 vdd.n841 0.026
R60390 vdd.n520 vdd.n519 0.026
R60391 vdd.n49 vdd.n48 0.026
R60392 vdd.n102 vdd.n101 0.026
R60393 vdd.n27641 vdd.n27255 0.026
R60394 vdd.n24903 vdd.n24894 0.026
R60395 vdd.n33430 vdd.n33429 0.026
R60396 vdd.n33437 vdd.n33436 0.026
R60397 vdd.n33545 vdd.n33544 0.026
R60398 vdd.n33569 vdd.n33566 0.026
R60399 vdd.n33588 vdd.n33587 0.026
R60400 vdd.n33830 vdd.n33829 0.026
R60401 vdd.n35567 vdd.n35566 0.026
R60402 vdd.n35527 vdd.n35518 0.026
R60403 vdd.n35268 vdd.n35267 0.026
R60404 vdd.n35081 vdd.n35080 0.026
R60405 vdd.n35330 vdd.n35329 0.026
R60406 vdd.n668 vdd.n667 0.026
R60407 vdd.n557 vdd.n556 0.026
R60408 vdd.n62 vdd.n61 0.026
R60409 vdd.n86 vdd.n85 0.026
R60410 vdd.n105 vdd.n95 0.026
R60411 vdd.n236 vdd.n235 0.026
R60412 vdd.n367 vdd.n366 0.026
R60413 vdd.n6022 vdd.n6021 0.026
R60414 vdd.n6009 vdd.n6008 0.026
R60415 vdd.n5835 vdd.n5834 0.026
R60416 vdd.n6175 vdd.n6174 0.026
R60417 vdd.n5899 vdd.n5898 0.026
R60418 vdd.n5150 vdd.n5149 0.026
R60419 vdd.n4754 vdd.n4753 0.026
R60420 vdd.n4576 vdd.n4575 0.026
R60421 vdd.n4563 vdd.n4562 0.026
R60422 vdd.n4261 vdd.n4260 0.026
R60423 vdd.n4320 vdd.n4319 0.026
R60424 vdd.n31104 vdd.n31103 0.026
R60425 vdd.n11761 vdd.n11680 0.026
R60426 vdd.n11760 vdd.n11678 0.026
R60427 vdd.n11886 vdd.n11881 0.026
R60428 vdd.n11899 vdd.n11794 0.026
R60429 vdd.n21763 vdd.n21762 0.026
R60430 vdd.n21841 vdd.n21840 0.026
R60431 vdd.n21977 vdd.n21972 0.026
R60432 vdd.n21990 vdd.n21885 0.026
R60433 vdd.n24886 vdd.n24885 0.026
R60434 vdd.n10179 vdd.n10178 0.026
R60435 vdd.n16776 vdd.n16775 0.026
R60436 vdd.n26062 vdd.n25677 0.026
R60437 vdd.n25953 vdd.n25952 0.026
R60438 vdd.n11890 vdd.n11889 0.025
R60439 vdd.n21981 vdd.n21980 0.025
R60440 vdd.n25484 vdd.n25483 0.025
R60441 vdd.n27347 vdd.n27345 0.025
R60442 vdd.n31852 vdd.n31697 0.025
R60443 vdd.n25799 vdd.n25797 0.025
R60444 vdd.n25478 vdd.n25477 0.025
R60445 vdd.n30508 vdd.n30323 0.025
R60446 vdd.n24965 vdd.n24964 0.025
R60447 vdd.n11881 vdd.n11800 0.025
R60448 vdd.n21972 vdd.n21891 0.025
R60449 vdd.n33414 vdd.n33413 0.025
R60450 vdd.n33339 vdd.n33338 0.025
R60451 vdd.n33715 vdd.n33711 0.025
R60452 vdd.n33703 vdd.n33702 0.025
R60453 vdd.n33634 vdd.n33633 0.025
R60454 vdd.n33671 vdd.n33666 0.025
R60455 vdd.n33814 vdd.n33812 0.025
R60456 vdd.n34088 vdd.n34084 0.025
R60457 vdd.n34274 vdd.n34273 0.025
R60458 vdd.n34309 vdd.n34307 0.025
R60459 vdd.n34249 vdd.n34248 0.025
R60460 vdd.n34150 vdd.n34146 0.025
R60461 vdd.n34244 vdd.n34243 0.025
R60462 vdd.n34150 vdd.n34149 0.025
R60463 vdd.n34167 vdd.n34166 0.025
R60464 vdd.n34193 vdd.n34188 0.025
R60465 vdd.n34207 vdd.n34201 0.025
R60466 vdd.n33962 vdd.n33886 0.025
R60467 vdd.n34390 vdd.n34389 0.025
R60468 vdd.n33939 vdd.n33938 0.025
R60469 vdd.n34414 vdd.n34413 0.025
R60470 vdd.n33973 vdd.n33972 0.025
R60471 vdd.n34037 vdd.n34036 0.025
R60472 vdd.n34038 vdd.n34037 0.025
R60473 vdd.n34041 vdd.n34040 0.025
R60474 vdd.n35309 vdd.n35308 0.025
R60475 vdd.n35575 vdd.n35573 0.025
R60476 vdd.n35540 vdd.n35539 0.025
R60477 vdd.n35249 vdd.n35245 0.025
R60478 vdd.n35114 vdd.n35111 0.025
R60479 vdd.n35303 vdd.n35298 0.025
R60480 vdd.n35291 vdd.n35285 0.025
R60481 vdd.n34662 vdd.n34658 0.025
R60482 vdd.n34929 vdd.n34928 0.025
R60483 vdd.n34904 vdd.n34902 0.025
R60484 vdd.n34982 vdd.n34981 0.025
R60485 vdd.n34688 vdd.n34666 0.025
R60486 vdd.n34971 vdd.n34970 0.025
R60487 vdd.n34688 vdd.n34687 0.025
R60488 vdd.n34733 vdd.n34732 0.025
R60489 vdd.n34719 vdd.n34714 0.025
R60490 vdd.n34707 vdd.n34701 0.025
R60491 vdd.n34527 vdd.n34524 0.025
R60492 vdd.n34482 vdd.n34481 0.025
R60493 vdd.n34841 vdd.n34840 0.025
R60494 vdd.n34844 vdd.n34843 0.025
R60495 vdd.n34545 vdd.n34544 0.025
R60496 vdd.n34570 vdd.n34569 0.025
R60497 vdd.n34617 vdd.n34616 0.025
R60498 vdd.n34618 vdd.n34617 0.025
R60499 vdd.n740 vdd.n739 0.025
R60500 vdd.n705 vdd.n694 0.025
R60501 vdd.n704 vdd.n703 0.025
R60502 vdd.n970 vdd.n969 0.025
R60503 vdd.n1045 vdd.n1044 0.025
R60504 vdd.n905 vdd.n901 0.025
R60505 vdd.n794 vdd.n793 0.025
R60506 vdd.n1091 vdd.n1090 0.025
R60507 vdd.n1064 vdd.n1059 0.025
R60508 vdd.n1056 vdd.n1055 0.025
R60509 vdd.n1122 vdd.n1107 0.025
R60510 vdd.n1139 vdd.n1138 0.025
R60511 vdd.n1138 vdd.n1137 0.025
R60512 vdd.n1122 vdd.n1121 0.025
R60513 vdd.n822 vdd.n820 0.025
R60514 vdd.n75 vdd.n26 0.025
R60515 vdd.n411 vdd.n410 0.025
R60516 vdd.n232 vdd.n228 0.025
R60517 vdd.n282 vdd.n264 0.025
R60518 vdd.n129 vdd.n128 0.025
R60519 vdd.n5868 vdd.n5867 0.025
R60520 vdd.n5947 vdd.n5945 0.025
R60521 vdd.n5972 vdd.n5971 0.025
R60522 vdd.n5790 vdd.n5786 0.025
R60523 vdd.n6247 vdd.n6160 0.025
R60524 vdd.n5894 vdd.n5889 0.025
R60525 vdd.n5908 vdd.n5902 0.025
R60526 vdd.n5409 vdd.n5405 0.025
R60527 vdd.n5676 vdd.n5675 0.025
R60528 vdd.n5651 vdd.n5649 0.025
R60529 vdd.n5729 vdd.n5728 0.025
R60530 vdd.n5435 vdd.n5413 0.025
R60531 vdd.n5718 vdd.n5717 0.025
R60532 vdd.n5435 vdd.n5434 0.025
R60533 vdd.n5480 vdd.n5479 0.025
R60534 vdd.n5466 vdd.n5461 0.025
R60535 vdd.n5454 vdd.n5448 0.025
R60536 vdd.n5274 vdd.n5271 0.025
R60537 vdd.n5229 vdd.n5228 0.025
R60538 vdd.n5588 vdd.n5587 0.025
R60539 vdd.n5591 vdd.n5590 0.025
R60540 vdd.n5291 vdd.n5290 0.025
R60541 vdd.n5317 vdd.n5316 0.025
R60542 vdd.n5364 vdd.n5363 0.025
R60543 vdd.n5365 vdd.n5364 0.025
R60544 vdd.n4653 vdd.n4652 0.025
R60545 vdd.n4635 vdd.n4633 0.025
R60546 vdd.n5099 vdd.n5096 0.025
R60547 vdd.n4833 vdd.n4830 0.025
R60548 vdd.n4856 vdd.n4835 0.025
R60549 vdd.n4825 vdd.n4819 0.025
R60550 vdd.n4814 vdd.n4810 0.025
R60551 vdd.n5088 vdd.n5087 0.025
R60552 vdd.n5087 vdd.n5086 0.025
R60553 vdd.n5054 vdd.n4969 0.025
R60554 vdd.n5027 vdd.n5026 0.025
R60555 vdd.n4239 vdd.n4235 0.025
R60556 vdd.n4503 vdd.n4502 0.025
R60557 vdd.n4478 vdd.n4476 0.025
R60558 vdd.n4307 vdd.n4306 0.025
R60559 vdd.n4293 vdd.n4288 0.025
R60560 vdd.n4281 vdd.n4275 0.025
R60561 vdd.n4104 vdd.n4101 0.025
R60562 vdd.n4071 vdd.n4070 0.025
R60563 vdd.n32492 vdd.n32416 0.025
R60564 vdd.n32075 vdd.n32074 0.025
R60565 vdd.n32104 vdd.n32103 0.025
R60566 vdd.n32245 vdd.n32241 0.025
R60567 vdd.n32520 vdd.n32518 0.025
R60568 vdd.n27296 vdd.n27295 0.025
R60569 vdd.n27443 vdd.n27441 0.025
R60570 vdd.n27331 vdd.n27326 0.025
R60571 vdd.n27343 vdd.n27337 0.025
R60572 vdd.n25748 vdd.n25747 0.025
R60573 vdd.n25889 vdd.n25887 0.025
R60574 vdd.n25783 vdd.n25778 0.025
R60575 vdd.n25795 vdd.n25789 0.025
R60576 vdd.n25500 vdd.n25499 0.025
R60577 vdd.n25623 vdd.n25622 0.025
R60578 vdd.n25615 vdd.n25614 0.025
R60579 vdd.n25495 vdd.n25492 0.025
R60580 vdd.n31788 vdd.n31731 0.025
R60581 vdd.n10207 vdd.n10206 0.025
R60582 vdd.n10213 vdd.n10212 0.025
R60583 vdd.n22241 vdd.n22240 0.025
R60584 vdd.n22215 vdd.n22214 0.025
R60585 vdd.n22107 vdd.n22106 0.025
R60586 vdd.n22067 vdd.n22066 0.025
R60587 vdd.n24309 vdd.n22061 0.025
R60588 vdd.n16735 vdd.n16734 0.025
R60589 vdd.n16684 vdd.n16683 0.025
R60590 vdd.n25496 vdd.n25495 0.025
R60591 vdd.n31615 vdd.n31611 0.025
R60592 vdd.n26703 vdd.n26693 0.025
R60593 vdd.n25516 vdd.n25514 0.025
R60594 vdd.n207 vdd.n206 0.025
R60595 vdd.n10094 vdd.n10092 0.025
R60596 vdd.n16740 vdd.n16739 0.025
R60597 vdd.n25674 vdd.n25673 0.025
R60598 vdd.n34232 vdd.n34158 0.025
R60599 bandgapmd_0.pnp_groupm_0.vdd vdd.n22471 0.024
R60600 vdd.n4347 vdd.n4265 0.024
R60601 vdd.n34773 vdd.n34691 0.024
R60602 vdd.n5520 vdd.n5438 0.024
R60603 vdd.n35357 vdd.n35275 0.024
R60604 vdd.n2097 vdd.n2096 0.024
R60605 vdd.n2754 vdd.n2752 0.024
R60606 vdd.n2848 vdd.n2846 0.024
R60607 vdd.n2935 vdd.n2933 0.024
R60608 vdd.n3029 vdd.n3027 0.024
R60609 vdd.n3116 vdd.n3114 0.024
R60610 vdd.n3210 vdd.n3208 0.024
R60611 vdd.n3297 vdd.n3295 0.024
R60612 vdd.n3391 vdd.n3389 0.024
R60613 vdd.n3478 vdd.n3476 0.024
R60614 vdd.n3572 vdd.n3570 0.024
R60615 vdd.n33434 vdd.n33433 0.024
R60616 vdd.n33538 vdd.n33537 0.024
R60617 vdd.n33566 vdd.n33565 0.024
R60618 vdd.n33542 vdd.n33541 0.024
R60619 vdd.n33663 vdd.n33662 0.024
R60620 vdd.n33662 vdd.n33661 0.024
R60621 vdd.n33606 vdd.n33596 0.024
R60622 vdd.n33605 vdd.n33604 0.024
R60623 vdd.n33763 vdd.n33762 0.024
R60624 vdd.n33767 vdd.n33766 0.024
R60625 vdd.n33840 vdd.n33839 0.024
R60626 vdd.n33901 vdd.n33900 0.024
R60627 vdd.n35577 vdd.n35576 0.024
R60628 vdd.n35516 vdd.n35515 0.024
R60629 vdd.n35463 vdd.n35462 0.024
R60630 vdd.n34494 vdd.n34493 0.024
R60631 vdd.n493 vdd.n492 0.024
R60632 vdd.n503 vdd.n502 0.024
R60633 vdd.n86 vdd.n83 0.024
R60634 vdd.n296 vdd.n295 0.024
R60635 vdd.n356 vdd.n355 0.024
R60636 vdd.n355 vdd.n354 0.024
R60637 vdd.n5940 vdd.n5939 0.024
R60638 vdd.n6006 vdd.n5984 0.024
R60639 vdd.n6134 vdd.n6060 0.024
R60640 vdd.n5241 vdd.n5240 0.024
R60641 vdd.n5139 vdd.n5138 0.024
R60642 vdd.n5138 vdd.n5137 0.024
R60643 vdd.n4744 vdd.n4743 0.024
R60644 vdd.n5023 vdd.n5022 0.024
R60645 vdd.n4616 vdd.n4615 0.024
R60646 vdd.n4471 vdd.n4470 0.024
R60647 vdd.n4560 vdd.n4559 0.024
R60648 vdd.n4548 vdd.n4547 0.024
R60649 vdd.n4262 vdd.n4261 0.024
R60650 vdd.n4059 vdd.n4058 0.024
R60651 vdd.n4415 vdd.n4414 0.024
R60652 vdd.n4448 vdd.n4447 0.024
R60653 vdd.n4195 vdd.n4194 0.024
R60654 vdd.n4196 vdd.n4195 0.024
R60655 vdd.n35862 vdd.n35860 0.024
R60656 vdd.n35981 vdd.n35979 0.024
R60657 vdd.n36093 vdd.n36091 0.024
R60658 vdd.n36212 vdd.n36210 0.024
R60659 vdd.n36324 vdd.n36322 0.024
R60660 vdd.n36443 vdd.n36441 0.024
R60661 vdd.n36555 vdd.n36553 0.024
R60662 vdd.n36674 vdd.n36672 0.024
R60663 vdd.n36786 vdd.n36784 0.024
R60664 vdd.n36905 vdd.n36903 0.024
R60665 vdd.n38072 vdd.n38070 0.024
R60666 vdd.n37960 vdd.n37958 0.024
R60667 vdd.n37841 vdd.n37839 0.024
R60668 vdd.n37729 vdd.n37727 0.024
R60669 vdd.n37610 vdd.n37608 0.024
R60670 vdd.n28283 vdd.n28281 0.024
R60671 vdd.n28402 vdd.n28400 0.024
R60672 vdd.n28514 vdd.n28512 0.024
R60673 vdd.n28633 vdd.n28631 0.024
R60674 vdd.n28745 vdd.n28743 0.024
R60675 vdd.n1697 vdd.n1695 0.024
R60676 vdd.n1610 vdd.n1608 0.024
R60677 vdd.n1516 vdd.n1514 0.024
R60678 vdd.n1429 vdd.n1427 0.024
R60679 vdd.n1335 vdd.n1333 0.024
R60680 vdd.n26801 vdd.n26799 0.024
R60681 vdd.n26895 vdd.n26893 0.024
R60682 vdd.n26982 vdd.n26980 0.024
R60683 vdd.n27076 vdd.n27074 0.024
R60684 vdd.n27163 vdd.n27161 0.024
R60685 vdd.n26547 vdd.n26546 0.024
R60686 vdd.n31693 vdd.n31691 0.024
R60687 vdd.n31852 vdd.n31699 0.024
R60688 vdd.n32276 vdd.n32275 0.024
R60689 vdd.n11743 vdd.n11721 0.024
R60690 vdd.n13211 vdd.n9174 0.024
R60691 vdd.n14402 vdd.n14401 0.024
R60692 vdd.n14707 vdd.n8116 0.024
R60693 vdd.n14708 vdd.n14707 0.024
R60694 vdd.n14795 vdd.n14794 0.024
R60695 vdd.n14880 vdd.n8027 0.024
R60696 vdd.n14881 vdd.n14880 0.024
R60697 vdd.n20629 vdd.n20628 0.024
R60698 vdd.n20392 vdd.n20391 0.024
R60699 vdd.n20391 vdd.n20385 0.024
R60700 vdd.n20271 vdd.n20270 0.024
R60701 vdd.n20156 vdd.n20155 0.024
R60702 vdd.n20155 vdd.n20149 0.024
R60703 vdd.n19423 vdd.n19422 0.024
R60704 vdd.n21825 vdd.n21824 0.024
R60705 vdd.n24909 vdd.n24908 0.024
R60706 vdd.n24946 vdd.n24945 0.024
R60707 vdd.n24562 vdd.n24561 0.024
R60708 vdd.n24574 vdd.n24572 0.024
R60709 vdd.n25830 vdd.n25828 0.024
R60710 vdd.n34071 vdd.n33974 0.024
R60711 vdd.n34646 vdd.n34548 0.024
R60712 vdd.n5393 vdd.n5295 0.024
R60713 vdd.n33701 vdd.n33572 0.024
R60714 vdd.n11768 vdd.n11767 0.024
R60715 vdd.n21853 vdd.n21852 0.024
R60716 vdd.n31981 vdd.n31635 0.024
R60717 vdd.n30203 vdd.n30202 0.024
R60718 vdd.n27936 vdd.n27935 0.024
R60719 vdd.n24969 vdd.n24968 0.024
R60720 vdd.n34156 vdd.n34155 0.024
R60721 vdd.n5848 vdd.n5841 0.023
R60722 vdd.n11745 vdd.n11723 0.023
R60723 vdd.n21827 vdd.n21804 0.023
R60724 vdd.n4711 vdd.n4608 0.023
R60725 vdd.n25560 vdd.n25559 0.023
R60726 vdd.n33381 vdd.n33380 0.023
R60727 vdd.n33391 vdd.n33390 0.023
R60728 vdd.n33940 vdd.n33939 0.023
R60729 vdd.n35504 vdd.n35503 0.023
R60730 vdd.n35272 vdd.n35268 0.023
R60731 vdd.n35069 vdd.n35068 0.023
R60732 vdd.n35438 vdd.n35437 0.023
R60733 vdd.n35199 vdd.n35198 0.023
R60734 vdd.n35200 vdd.n35199 0.023
R60735 vdd.n34483 vdd.n34482 0.023
R60736 vdd.n439 vdd.n438 0.023
R60737 vdd.n6005 vdd.n6004 0.023
R60738 vdd.n5836 vdd.n5835 0.023
R60739 vdd.n6223 vdd.n6222 0.023
R60740 vdd.n6118 vdd.n6117 0.023
R60741 vdd.n6328 vdd.n6327 0.023
R60742 vdd.n6329 vdd.n6328 0.023
R60743 vdd.n5230 vdd.n5229 0.023
R60744 vdd.n5088 vdd.n5076 0.023
R60745 vdd.n5076 vdd.n5075 0.023
R60746 vdd.n4868 vdd.n4867 0.023
R60747 vdd.n4809 vdd.n4808 0.023
R60748 vdd.n5024 vdd.n5023 0.023
R60749 vdd.n4799 vdd.n4798 0.023
R60750 vdd.n4685 vdd.n4684 0.023
R60751 vdd.n4891 vdd.n4890 0.023
R60752 vdd.n4122 vdd.n4121 0.023
R60753 vdd.n29491 vdd.n29482 0.023
R60754 vdd.n32812 vdd.n6391 0.023
R60755 vdd.n26092 vdd.n25358 0.023
R60756 vdd.n30975 vdd.n30974 0.023
R60757 vdd.n31356 vdd.n31352 0.023
R60758 vdd.n31337 vdd.n31332 0.023
R60759 vdd.n30883 vdd.n30882 0.023
R60760 vdd.n30905 vdd.n30904 0.023
R60761 vdd.n30711 vdd.n30703 0.023
R60762 vdd.n30711 vdd.n30710 0.023
R60763 vdd.n32605 vdd.n32604 0.023
R60764 vdd.n30145 vdd.n30144 0.023
R60765 vdd.n29578 vdd.n29570 0.023
R60766 vdd.n29578 vdd.n29577 0.023
R60767 vdd.n29601 vdd.n29600 0.023
R60768 vdd.n7173 vdd.n7157 0.023
R60769 vdd.n32739 vdd.n7137 0.023
R60770 vdd.n29380 vdd.n29379 0.023
R60771 vdd.n29359 vdd.n29358 0.023
R60772 vdd.n27673 vdd.n27672 0.023
R60773 vdd.n27695 vdd.n27694 0.023
R60774 vdd.n26524 vdd.n26480 0.023
R60775 vdd.n26241 vdd.n26232 0.023
R60776 vdd.n26241 vdd.n26240 0.023
R60777 vdd.n25344 vdd.n25340 0.023
R60778 vdd.n26083 vdd.n26081 0.023
R60779 vdd.n26711 vdd.n26630 0.023
R60780 vdd.n26407 vdd.n26362 0.023
R60781 vdd.n29464 vdd.n29446 0.023
R60782 vdd.n32703 vdd.n32691 0.023
R60783 vdd.n32703 vdd.n32686 0.023
R60784 vdd.n29671 vdd.n29652 0.023
R60785 vdd.n30125 vdd.n30113 0.023
R60786 vdd.n32563 vdd.n32545 0.023
R60787 vdd.n30924 vdd.n30923 0.023
R60788 vdd.n29619 vdd.n29618 0.023
R60789 vdd.n7173 vdd.n7162 0.023
R60790 vdd.n29336 vdd.n29324 0.023
R60791 vdd.n29336 vdd.n29320 0.023
R60792 vdd.n29101 vdd.n29054 0.023
R60793 vdd.n27713 vdd.n27712 0.023
R60794 vdd.n26524 vdd.n26490 0.023
R60795 vdd.n26217 vdd.n26105 0.023
R60796 vdd.n30767 vdd.n30759 0.023
R60797 vdd.n30767 vdd.n30750 0.023
R60798 vdd.n30813 vdd.n30791 0.023
R60799 vdd.n30860 vdd.n30855 0.023
R60800 vdd.n32563 vdd.n32558 0.023
R60801 vdd.n29995 vdd.n29991 0.023
R60802 vdd.n29671 vdd.n29666 0.023
R60803 vdd.n29530 vdd.n29523 0.023
R60804 vdd.n7173 vdd.n7168 0.023
R60805 vdd.n29464 vdd.n29459 0.023
R60806 vdd.n26472 vdd.n26449 0.023
R60807 vdd.n26407 vdd.n26375 0.023
R60808 vdd.n26181 vdd.n26144 0.023
R60809 vdd.n31002 vdd.n31001 0.023
R60810 vdd.n30831 vdd.n30823 0.023
R60811 vdd.n30104 vdd.n30096 0.023
R60812 vdd.n7173 vdd.n7165 0.023
R60813 vdd.n29552 vdd.n29544 0.023
R60814 vdd.n29311 vdd.n29303 0.023
R60815 vdd.n26524 vdd.n26494 0.023
R60816 vdd.n26673 vdd.n26650 0.023
R60817 vdd.n25370 vdd.n25368 0.023
R60818 vdd.n31300 vdd.n31299 0.023
R60819 vdd.n31225 vdd.n31217 0.023
R60820 vdd.n31225 vdd.n31224 0.023
R60821 vdd.n30767 vdd.n30760 0.023
R60822 vdd.n30860 vdd.n30856 0.023
R60823 vdd.n31428 vdd.n31426 0.023
R60824 vdd.n32563 vdd.n32559 0.023
R60825 vdd.n29995 vdd.n29992 0.023
R60826 vdd.n29671 vdd.n29667 0.023
R60827 vdd.n32678 vdd.n32676 0.023
R60828 vdd.n32703 vdd.n32699 0.023
R60829 vdd.n7173 vdd.n7169 0.023
R60830 vdd.n29432 vdd.n29430 0.023
R60831 vdd.n29464 vdd.n29460 0.023
R60832 vdd.n29336 vdd.n29332 0.023
R60833 vdd.n29097 vdd.n29076 0.023
R60834 vdd.n29101 vdd.n29061 0.023
R60835 vdd.n29093 vdd.n29079 0.023
R60836 vdd.n26524 vdd.n26499 0.023
R60837 vdd.n26320 vdd.n26284 0.023
R60838 vdd.n26407 vdd.n26376 0.023
R60839 vdd.n26217 vdd.n26098 0.023
R60840 vdd.n4000 vdd.n3736 0.023
R60841 vdd.n3959 vdd.n3773 0.023
R60842 vdd.n31718 vdd.n31717 0.023
R60843 vdd.n29311 vdd.n29286 0.023
R60844 vdd.n29464 vdd.n29414 0.023
R60845 vdd.n7173 vdd.n7156 0.023
R60846 vdd.n29530 vdd.n29500 0.023
R60847 vdd.n29671 vdd.n29634 0.023
R60848 vdd.n30104 vdd.n30079 0.023
R60849 vdd.n30767 vdd.n30735 0.023
R60850 vdd.n31236 vdd.n31189 0.023
R60851 vdd.n31247 vdd.n31017 0.023
R60852 vdd.n31302 vdd.n31016 0.023
R60853 vdd.n26472 vdd.n26455 0.023
R60854 vdd.n26407 vdd.n26352 0.023
R60855 vdd.n26673 vdd.n26657 0.023
R60856 vdd.n11867 vdd.n11811 0.023
R60857 vdd.n13086 vdd.n9270 0.023
R60858 vdd.n14495 vdd.n14494 0.023
R60859 vdd.n14652 vdd.n8151 0.023
R60860 vdd.n14974 vdd.n7982 0.023
R60861 vdd.n24192 vdd.n24190 0.023
R60862 vdd.n23984 vdd.n23982 0.023
R60863 vdd.n23960 vdd.n23958 0.023
R60864 vdd.n23752 vdd.n23750 0.023
R60865 vdd.n23728 vdd.n23726 0.023
R60866 vdd.n23064 vdd.n23062 0.023
R60867 vdd.n23272 vdd.n23270 0.023
R60868 vdd.n23296 vdd.n23294 0.023
R60869 vdd.n23504 vdd.n23502 0.023
R60870 vdd.n23528 vdd.n23526 0.023
R60871 vdd.n22485 vdd.n22483 0.023
R60872 vdd.n22693 vdd.n22691 0.023
R60873 vdd.n22717 vdd.n22715 0.023
R60874 vdd.n22925 vdd.n22923 0.023
R60875 vdd.n22949 vdd.n22947 0.023
R60876 vdd.n20547 vdd.n19969 0.023
R60877 vdd.n20467 vdd.n19987 0.023
R60878 vdd.n20065 vdd.n20026 0.023
R60879 vdd.n19338 vdd.n19299 0.023
R60880 vdd.n21958 vdd.n21902 0.023
R60881 vdd.n24935 vdd.n24934 0.023
R60882 vdd.n24947 vdd.n24946 0.023
R60883 vdd.n24561 vdd.n24560 0.023
R60884 vdd.n10210 vdd.n10205 0.023
R60885 vdd.n16783 vdd.n16782 0.023
R60886 vdd.n32492 vdd.n32491 0.023
R60887 vdd.n2353 vdd.n2107 0.023
R60888 vdd.n1799 vdd.n1260 0.023
R60889 vdd.n27592 vdd.n27591 0.023
R60890 vdd.n26008 vdd.n26007 0.023
R60891 vdd.n27803 vdd.n27802 0.022
R60892 vdd.n35528 vdd.n35527 0.022
R60893 vdd.n6010 vdd.n6009 0.022
R60894 vdd.n30820 vdd.n30817 0.022
R60895 vdd.n26387 vdd.n26386 0.022
R60896 vdd.n4662 vdd.n4661 0.022
R60897 vdd.n24543 vdd.n24542 0.022
R60898 vdd.n27387 vdd.n27385 0.022
R60899 vdd.n4564 vdd.n4563 0.022
R60900 vdd.n27815 vdd.n27803 0.022
R60901 vdd.n22471 vdd.n22470 0.022
R60902 vdd.n26023 vdd.n26022 0.022
R60903 vdd.n27607 vdd.n27606 0.022
R60904 vdd.n34262 vdd.n34261 0.022
R60905 vdd.n34987 vdd.n34986 0.022
R60906 vdd.n5734 vdd.n5733 0.022
R60907 vdd.n4223 vdd.n4125 0.022
R60908 vdd.n32463 vdd.n32462 0.022
R60909 vdd.n30013 vdd.n30012 0.022
R60910 vdd.n33394 vdd.n33393 0.022
R60911 vdd.n33395 vdd.n33394 0.022
R60912 vdd.n33405 vdd.n33402 0.022
R60913 vdd.n33492 vdd.n33491 0.022
R60914 vdd.n33517 vdd.n33516 0.022
R60915 vdd.n33528 vdd.n33525 0.022
R60916 vdd.n33307 vdd.n33306 0.022
R60917 vdd.n33332 vdd.n33329 0.022
R60918 vdd.n33341 vdd.n33340 0.022
R60919 vdd.n33726 vdd.n33725 0.022
R60920 vdd.n33590 vdd.n33589 0.022
R60921 vdd.n33602 vdd.n33601 0.022
R60922 vdd.n33630 vdd.n33629 0.022
R60923 vdd.n33644 vdd.n33641 0.022
R60924 vdd.n34097 vdd.n34092 0.022
R60925 vdd.n34106 vdd.n34103 0.022
R60926 vdd.n34246 vdd.n34245 0.022
R60927 vdd.n34295 vdd.n34292 0.022
R60928 vdd.n34317 vdd.n34316 0.022
R60929 vdd.n34316 vdd.n34315 0.022
R60930 vdd.n34302 vdd.n34301 0.022
R60931 vdd.n34250 vdd.n34249 0.022
R60932 vdd.n34311 vdd.n34310 0.022
R60933 vdd.n34250 vdd.n34244 0.022
R60934 vdd.n34197 vdd.n34196 0.022
R60935 vdd.n34370 vdd.n34369 0.022
R60936 vdd.n34382 vdd.n34381 0.022
R60937 vdd.n33904 vdd.n33903 0.022
R60938 vdd.n33892 vdd.n33891 0.022
R60939 vdd.n33962 vdd.n33873 0.022
R60940 vdd.n33872 vdd.n33871 0.022
R60941 vdd.n34439 vdd.n34354 0.022
R60942 vdd.n34413 vdd.n34412 0.022
R60943 vdd.n34439 vdd.n34438 0.022
R60944 vdd.n33976 vdd.n33975 0.022
R60945 vdd.n33985 vdd.n33984 0.022
R60946 vdd.n33991 vdd.n33986 0.022
R60947 vdd.n33996 vdd.n33993 0.022
R60948 vdd.n34008 vdd.n34007 0.022
R60949 vdd.n35170 vdd.n35169 0.022
R60950 vdd.n35158 vdd.n35155 0.022
R60951 vdd.n35147 vdd.n35146 0.022
R60952 vdd.n35153 vdd.n35148 0.022
R60953 vdd.n35583 vdd.n35582 0.022
R60954 vdd.n35582 vdd.n35581 0.022
R60955 vdd.n35561 vdd.n35558 0.022
R60956 vdd.n35512 vdd.n35511 0.022
R60957 vdd.n35511 vdd.n35510 0.022
R60958 vdd.n35486 vdd.n35485 0.022
R60959 vdd.n35258 vdd.n35253 0.022
R60960 vdd.n35123 vdd.n35122 0.022
R60961 vdd.n35114 vdd.n35031 0.022
R60962 vdd.n35086 vdd.n35085 0.022
R60963 vdd.n35073 vdd.n35072 0.022
R60964 vdd.n35401 vdd.n35400 0.022
R60965 vdd.n35393 vdd.n35392 0.022
R60966 vdd.n35070 vdd.n35069 0.022
R60967 vdd.n35129 vdd.n35128 0.022
R60968 vdd.n35138 vdd.n35137 0.022
R60969 vdd.n34674 vdd.n34669 0.022
R60970 vdd.n34961 vdd.n34957 0.022
R60971 vdd.n34979 vdd.n34978 0.022
R60972 vdd.n34978 vdd.n34977 0.022
R60973 vdd.n34911 vdd.n34908 0.022
R60974 vdd.n34889 vdd.n34888 0.022
R60975 vdd.n34888 vdd.n34887 0.022
R60976 vdd.n34897 vdd.n34896 0.022
R60977 vdd.n34983 vdd.n34982 0.022
R60978 vdd.n35000 vdd.n34999 0.022
R60979 vdd.n34983 vdd.n34971 0.022
R60980 vdd.n34745 vdd.n34744 0.022
R60981 vdd.n34796 vdd.n34795 0.022
R60982 vdd.n34805 vdd.n34804 0.022
R60983 vdd.n34486 vdd.n34485 0.022
R60984 vdd.n34499 vdd.n34498 0.022
R60985 vdd.n34527 vdd.n34445 0.022
R60986 vdd.n34536 vdd.n34535 0.022
R60987 vdd.n34840 vdd.n34839 0.022
R60988 vdd.n34874 vdd.n34871 0.022
R60989 vdd.n34874 vdd.n34873 0.022
R60990 vdd.n34551 vdd.n34550 0.022
R60991 vdd.n34562 vdd.n34561 0.022
R60992 vdd.n34568 vdd.n34563 0.022
R60993 vdd.n34576 vdd.n34573 0.022
R60994 vdd.n34592 vdd.n34591 0.022
R60995 vdd.n713 vdd.n712 0.022
R60996 vdd.n714 vdd.n713 0.022
R60997 vdd.n726 vdd.n723 0.022
R60998 vdd.n728 vdd.n727 0.022
R60999 vdd.n754 vdd.n753 0.022
R61000 vdd.n979 vdd.n978 0.022
R61001 vdd.n998 vdd.n997 0.022
R61002 vdd.n1011 vdd.n1008 0.022
R61003 vdd.n636 vdd.n635 0.022
R61004 vdd.n621 vdd.n618 0.022
R61005 vdd.n607 vdd.n606 0.022
R61006 vdd.n1015 vdd.n1014 0.022
R61007 vdd.n667 vdd.n666 0.022
R61008 vdd.n1018 vdd.n1017 0.022
R61009 vdd.n890 vdd.n889 0.022
R61010 vdd.n950 vdd.n949 0.022
R61011 vdd.n1113 vdd.n1112 0.022
R61012 vdd.n1087 vdd.n1086 0.022
R61013 vdd.n1081 vdd.n1078 0.022
R61014 vdd.n1107 vdd.n1106 0.022
R61015 vdd.n899 vdd.n893 0.022
R61016 vdd.n907 vdd.n906 0.022
R61017 vdd.n1121 vdd.n1120 0.022
R61018 vdd.n899 vdd.n898 0.022
R61019 vdd.n909 vdd.n908 0.022
R61020 vdd.n512 vdd.n511 0.022
R61021 vdd.n523 vdd.n520 0.022
R61022 vdd.n534 vdd.n533 0.022
R61023 vdd.n41 vdd.n40 0.022
R61024 vdd.n42 vdd.n41 0.022
R61025 vdd.n437 vdd.n434 0.022
R61026 vdd.n445 vdd.n444 0.022
R61027 vdd.n444 vdd.n443 0.022
R61028 vdd.n245 vdd.n244 0.022
R61029 vdd.n133 vdd.n132 0.022
R61030 vdd.n143 vdd.n140 0.022
R61031 vdd.n170 vdd.n165 0.022
R61032 vdd.n164 vdd.n163 0.022
R61033 vdd.n339 vdd.n337 0.022
R61034 vdd.n6303 vdd.n6302 0.022
R61035 vdd.n6287 vdd.n6284 0.022
R61036 vdd.n6273 vdd.n6272 0.022
R61037 vdd.n6279 vdd.n6274 0.022
R61038 vdd.n5932 vdd.n5931 0.022
R61039 vdd.n5931 vdd.n5930 0.022
R61040 vdd.n5954 vdd.n5951 0.022
R61041 vdd.n5992 vdd.n5991 0.022
R61042 vdd.n5991 vdd.n5990 0.022
R61043 vdd.n5814 vdd.n5811 0.022
R61044 vdd.n5802 vdd.n5797 0.022
R61045 vdd.n6146 vdd.n6145 0.022
R61046 vdd.n6247 vdd.n6147 0.022
R61047 vdd.n6166 vdd.n6165 0.022
R61048 vdd.n6178 vdd.n6177 0.022
R61049 vdd.n6095 vdd.n6094 0.022
R61050 vdd.n6084 vdd.n6083 0.022
R61051 vdd.n6224 vdd.n6223 0.022
R61052 vdd.n6258 vdd.n6257 0.022
R61053 vdd.n6261 vdd.n6260 0.022
R61054 vdd.n5421 vdd.n5416 0.022
R61055 vdd.n5708 vdd.n5704 0.022
R61056 vdd.n5726 vdd.n5725 0.022
R61057 vdd.n5725 vdd.n5724 0.022
R61058 vdd.n5658 vdd.n5655 0.022
R61059 vdd.n5636 vdd.n5635 0.022
R61060 vdd.n5635 vdd.n5634 0.022
R61061 vdd.n5644 vdd.n5643 0.022
R61062 vdd.n5730 vdd.n5729 0.022
R61063 vdd.n5747 vdd.n5746 0.022
R61064 vdd.n5730 vdd.n5718 0.022
R61065 vdd.n5492 vdd.n5491 0.022
R61066 vdd.n5543 vdd.n5542 0.022
R61067 vdd.n5552 vdd.n5551 0.022
R61068 vdd.n5233 vdd.n5232 0.022
R61069 vdd.n5246 vdd.n5245 0.022
R61070 vdd.n5274 vdd.n5192 0.022
R61071 vdd.n5283 vdd.n5282 0.022
R61072 vdd.n5587 vdd.n5586 0.022
R61073 vdd.n5621 vdd.n5618 0.022
R61074 vdd.n5621 vdd.n5620 0.022
R61075 vdd.n5298 vdd.n5297 0.022
R61076 vdd.n5309 vdd.n5308 0.022
R61077 vdd.n5315 vdd.n5310 0.022
R61078 vdd.n5323 vdd.n5320 0.022
R61079 vdd.n5339 vdd.n5338 0.022
R61080 vdd.n4640 vdd.n4637 0.022
R61081 vdd.n5155 vdd.n5154 0.022
R61082 vdd.n5148 vdd.n5143 0.022
R61083 vdd.n5142 vdd.n5141 0.022
R61084 vdd.n5132 vdd.n5129 0.022
R61085 vdd.n5113 vdd.n5112 0.022
R61086 vdd.n5084 vdd.n5083 0.022
R61087 vdd.n4837 vdd.n4836 0.022
R61088 vdd.n4759 vdd.n4758 0.022
R61089 vdd.n4746 vdd.n4745 0.022
R61090 vdd.n4983 vdd.n4982 0.022
R61091 vdd.n4974 vdd.n4973 0.022
R61092 vdd.n5054 vdd.n5051 0.022
R61093 vdd.n4958 vdd.n4957 0.022
R61094 vdd.n4622 vdd.n4621 0.022
R61095 vdd.n4623 vdd.n4622 0.022
R61096 vdd.n4888 vdd.n4883 0.022
R61097 vdd.n4883 vdd.n4882 0.022
R61098 vdd.n4882 vdd.n4881 0.022
R61099 vdd.n4251 vdd.n4246 0.022
R61100 vdd.n4535 vdd.n4531 0.022
R61101 vdd.n4556 vdd.n4555 0.022
R61102 vdd.n4555 vdd.n4554 0.022
R61103 vdd.n4485 vdd.n4482 0.022
R61104 vdd.n4463 vdd.n4462 0.022
R61105 vdd.n4462 vdd.n4461 0.022
R61106 vdd.n4370 vdd.n4369 0.022
R61107 vdd.n4378 vdd.n4377 0.022
R61108 vdd.n4063 vdd.n4062 0.022
R61109 vdd.n4076 vdd.n4075 0.022
R61110 vdd.n4104 vdd.n4022 0.022
R61111 vdd.n4113 vdd.n4112 0.022
R61112 vdd.n4060 vdd.n4059 0.022
R61113 vdd.n4128 vdd.n4127 0.022
R61114 vdd.n4140 vdd.n4139 0.022
R61115 vdd.n4146 vdd.n4141 0.022
R61116 vdd.n4154 vdd.n4151 0.022
R61117 vdd.n4170 vdd.n4169 0.022
R61118 vdd.n27610 vdd.n27609 0.022
R61119 vdd.n27621 vdd.n27620 0.022
R61120 vdd.n27619 vdd.n27618 0.022
R61121 vdd.n27630 vdd.n27629 0.022
R61122 vdd.n27491 vdd.n27490 0.022
R61123 vdd.n27502 vdd.n27501 0.022
R61124 vdd.n27538 vdd.n27537 0.022
R61125 vdd.n27549 vdd.n27548 0.022
R61126 vdd.n27373 vdd.n27372 0.022
R61127 vdd.n27384 vdd.n27380 0.022
R61128 vdd.n27401 vdd.n27400 0.022
R61129 vdd.n27400 vdd.n27399 0.022
R61130 vdd.n27432 vdd.n27429 0.022
R61131 vdd.n27449 vdd.n27448 0.022
R61132 vdd.n27448 vdd.n27447 0.022
R61133 vdd.n27311 vdd.n27309 0.022
R61134 vdd.n26031 vdd.n26030 0.022
R61135 vdd.n26042 vdd.n26041 0.022
R61136 vdd.n26040 vdd.n26039 0.022
R61137 vdd.n26051 vdd.n26050 0.022
R61138 vdd.n25928 vdd.n25927 0.022
R61139 vdd.n25939 vdd.n25938 0.022
R61140 vdd.n25975 vdd.n25974 0.022
R61141 vdd.n25986 vdd.n25985 0.022
R61142 vdd.n25741 vdd.n25740 0.022
R61143 vdd.n25827 vdd.n25823 0.022
R61144 vdd.n25847 vdd.n25846 0.022
R61145 vdd.n25846 vdd.n25845 0.022
R61146 vdd.n25878 vdd.n25875 0.022
R61147 vdd.n25895 vdd.n25894 0.022
R61148 vdd.n25894 vdd.n25893 0.022
R61149 vdd.n25763 vdd.n25761 0.022
R61150 vdd.n25499 vdd.n25498 0.022
R61151 vdd.n25658 vdd.n25657 0.022
R61152 vdd.n25408 vdd.n25407 0.022
R61153 vdd.n25624 vdd.n25623 0.022
R61154 vdd.n25573 vdd.n25572 0.022
R61155 vdd.n25546 vdd.n25545 0.022
R61156 vdd.n25460 vdd.n25459 0.022
R61157 vdd.n31959 vdd.n31958 0.022
R61158 vdd.n32055 vdd.n32054 0.022
R61159 vdd.n10251 vdd.n10124 0.022
R61160 vdd.n10214 vdd.n10213 0.022
R61161 vdd.n11492 vdd.n11467 0.022
R61162 vdd.n11498 vdd.n11497 0.022
R61163 vdd.n11508 vdd.n11507 0.022
R61164 vdd.n11555 vdd.n11553 0.022
R61165 vdd.n11592 vdd.n11591 0.022
R61166 vdd.n11623 vdd.n11622 0.022
R61167 vdd.n12622 vdd.n10052 0.022
R61168 vdd.n11768 vdd.n11671 0.022
R61169 vdd.n24104 vdd.n24094 0.022
R61170 vdd.n24080 vdd.n24078 0.022
R61171 vdd.n23872 vdd.n23862 0.022
R61172 vdd.n23848 vdd.n23846 0.022
R61173 vdd.n23640 vdd.n23630 0.022
R61174 vdd.n23160 vdd.n23158 0.022
R61175 vdd.n23184 vdd.n23174 0.022
R61176 vdd.n23392 vdd.n23390 0.022
R61177 vdd.n23416 vdd.n23406 0.022
R61178 vdd.n23624 vdd.n23622 0.022
R61179 vdd.n22581 vdd.n22579 0.022
R61180 vdd.n22605 vdd.n22595 0.022
R61181 vdd.n22813 vdd.n22811 0.022
R61182 vdd.n22837 vdd.n22827 0.022
R61183 vdd.n23045 vdd.n23043 0.022
R61184 vdd.n16685 vdd.n16684 0.022
R61185 vdd.n18312 vdd.n18311 0.022
R61186 vdd.n18317 vdd.n18316 0.022
R61187 vdd.n18334 vdd.n18333 0.022
R61188 vdd.n18391 vdd.n18390 0.022
R61189 vdd.n18407 vdd.n18406 0.022
R61190 vdd.n21648 vdd.n21647 0.022
R61191 vdd.n16756 vdd.n16755 0.022
R61192 vdd.n21855 vdd.n21853 0.022
R61193 vdd.n24936 vdd.n24935 0.022
R61194 vdd.n11744 vdd.n11743 0.022
R61195 vdd.n21826 vdd.n21825 0.022
R61196 vdd.n31967 vdd.n31647 0.022
R61197 vdd.n26620 vdd.n26586 0.022
R61198 vdd.n4800 vdd.n4711 0.022
R61199 vdd.n33780 vdd.n33773 0.022
R61200 vdd.n388 vdd.n383 0.022
R61201 vdd.n25556 vdd.n25555 0.022
R61202 vdd.n28099 vdd.n28098 0.022
R61203 vdd.n33860 vdd.n33859 0.022
R61204 vdd.n961 vdd.n960 0.022
R61205 vdd.n27843 vdd.n27842 0.021
R61206 vdd.n28105 vdd.n28104 0.021
R61207 vdd.n10197 vdd.n10135 0.021
R61208 vdd.n12574 vdd.n10259 0.021
R61209 vdd.n16778 vdd.n16777 0.021
R61210 vdd.n16795 vdd.n16794 0.021
R61211 vdd.n29315 vdd.n29314 0.021
R61212 vdd.n7155 vdd.n7153 0.021
R61213 vdd.n30108 vdd.n30107 0.021
R61214 vdd.n30833 vdd.n30728 0.021
R61215 vdd.n30771 vdd.n30770 0.021
R61216 vdd.n26710 vdd.n26642 0.021
R61217 vdd.n29185 vdd.n29184 0.021
R61218 vdd.n29534 vdd.n29533 0.021
R61219 vdd.n32645 vdd.n32644 0.021
R61220 vdd.n29961 vdd.n29960 0.021
R61221 vdd.n32538 vdd.n32537 0.021
R61222 vdd.n30816 vdd.n30815 0.021
R61223 vdd.n29044 vdd.n29043 0.021
R61224 vdd.n26476 vdd.n26475 0.021
R61225 vdd.n210 vdd.n86 0.021
R61226 vdd.n32737 vdd.n27682 0.021
R61227 vdd.n35233 vdd.n35135 0.021
R61228 vdd.n6356 vdd.n6259 0.021
R61229 vdd.n27755 vdd.n27754 0.021
R61230 vdd.n10167 vdd.n10166 0.021
R61231 vdd.n16769 vdd.n16582 0.021
R61232 vdd.n34071 vdd.n34070 0.021
R61233 vdd.n2752 vdd.n2750 0.021
R61234 vdd.n2855 vdd.n2848 0.021
R61235 vdd.n2933 vdd.n2931 0.021
R61236 vdd.n3036 vdd.n3029 0.021
R61237 vdd.n3114 vdd.n3112 0.021
R61238 vdd.n3217 vdd.n3210 0.021
R61239 vdd.n3295 vdd.n3293 0.021
R61240 vdd.n3398 vdd.n3391 0.021
R61241 vdd.n3476 vdd.n3474 0.021
R61242 vdd.n3579 vdd.n3572 0.021
R61243 vdd.n33431 vdd.n33430 0.021
R61244 vdd.n33338 vdd.n33337 0.021
R61245 vdd.n33539 vdd.n33538 0.021
R61246 vdd.n33596 vdd.n33595 0.021
R61247 vdd.n33763 vdd.n33759 0.021
R61248 vdd.n33765 vdd.n33764 0.021
R61249 vdd.n33831 vdd.n33830 0.021
R61250 vdd.n35526 vdd.n35525 0.021
R61251 vdd.n35244 vdd.n35243 0.021
R61252 vdd.n35126 vdd.n35125 0.021
R61253 vdd.n35435 vdd.n35434 0.021
R61254 vdd.n35294 vdd.n35293 0.021
R61255 vdd.n556 vdd.n555 0.021
R61256 vdd.n432 vdd.n431 0.021
R61257 vdd.n59 vdd.n58 0.021
R61258 vdd.n161 vdd.n160 0.021
R61259 vdd.n104 vdd.n103 0.021
R61260 vdd.n93 vdd.n92 0.021
R61261 vdd.n5976 vdd.n5975 0.021
R61262 vdd.n5840 vdd.n5839 0.021
R61263 vdd.n6250 vdd.n6139 0.021
R61264 vdd.n6111 vdd.n6110 0.021
R61265 vdd.n5896 vdd.n5895 0.021
R61266 vdd.n4868 vdd.n4864 0.021
R61267 vdd.n4870 vdd.n4869 0.021
R61268 vdd.n4799 vdd.n4789 0.021
R61269 vdd.n4743 vdd.n4742 0.021
R61270 vdd.n4682 vdd.n4681 0.021
R61271 vdd.n4921 vdd.n4920 0.021
R61272 vdd.n4577 vdd.n4576 0.021
R61273 vdd.n4560 vdd.n4548 0.021
R61274 vdd.n4319 vdd.n4318 0.021
R61275 vdd.n4414 vdd.n4413 0.021
R61276 vdd.n4448 vdd.n4445 0.021
R61277 vdd.n35860 vdd.n35858 0.021
R61278 vdd.n35991 vdd.n35981 0.021
R61279 vdd.n36091 vdd.n36089 0.021
R61280 vdd.n36222 vdd.n36212 0.021
R61281 vdd.n36322 vdd.n36320 0.021
R61282 vdd.n36453 vdd.n36443 0.021
R61283 vdd.n36553 vdd.n36551 0.021
R61284 vdd.n36684 vdd.n36674 0.021
R61285 vdd.n36784 vdd.n36782 0.021
R61286 vdd.n36915 vdd.n36905 0.021
R61287 vdd.n38070 vdd.n38068 0.021
R61288 vdd.n37970 vdd.n37960 0.021
R61289 vdd.n37839 vdd.n37837 0.021
R61290 vdd.n37739 vdd.n37729 0.021
R61291 vdd.n37608 vdd.n37606 0.021
R61292 vdd.n28281 vdd.n28279 0.021
R61293 vdd.n28412 vdd.n28402 0.021
R61294 vdd.n28512 vdd.n28510 0.021
R61295 vdd.n28643 vdd.n28633 0.021
R61296 vdd.n28743 vdd.n28741 0.021
R61297 vdd.n1695 vdd.n1693 0.021
R61298 vdd.n1617 vdd.n1610 0.021
R61299 vdd.n1514 vdd.n1512 0.021
R61300 vdd.n1436 vdd.n1429 0.021
R61301 vdd.n1333 vdd.n1331 0.021
R61302 vdd.n26799 vdd.n26797 0.021
R61303 vdd.n26902 vdd.n26895 0.021
R61304 vdd.n26980 vdd.n26978 0.021
R61305 vdd.n27083 vdd.n27076 0.021
R61306 vdd.n27161 vdd.n27159 0.021
R61307 vdd.n31245 vdd.n31244 0.021
R61308 vdd.n3695 vdd.n2695 0.021
R61309 vdd.n32500 vdd.n32499 0.021
R61310 vdd.n10209 vdd.n10208 0.021
R61311 vdd.n10218 vdd.n10217 0.021
R61312 vdd.n10232 vdd.n10074 0.021
R61313 vdd.n10226 vdd.n10130 0.021
R61314 vdd.n11491 vdd.n11490 0.021
R61315 vdd.n11496 vdd.n11463 0.021
R61316 vdd.n11593 vdd.n11588 0.021
R61317 vdd.n16737 vdd.n16736 0.021
R61318 vdd.n16590 vdd.n16589 0.021
R61319 vdd.n16676 vdd.n16674 0.021
R61320 vdd.n16808 vdd.n16807 0.021
R61321 vdd.n16804 vdd.n16803 0.021
R61322 vdd.n18430 vdd.n18429 0.021
R61323 vdd.n25001 vdd.n24998 0.021
R61324 vdd.n24577 vdd.n24574 0.021
R61325 vdd.n24693 vdd.n24685 0.021
R61326 vdd.n24705 vdd.n24697 0.021
R61327 vdd.n24717 vdd.n24709 0.021
R61328 vdd.n24744 vdd.n24734 0.021
R61329 vdd.n24760 vdd.n24758 0.021
R61330 vdd.n24772 vdd.n24770 0.021
R61331 vdd.n24784 vdd.n24782 0.021
R61332 vdd.n24796 vdd.n24794 0.021
R61333 vdd.n24808 vdd.n24806 0.021
R61334 vdd.n24820 vdd.n24818 0.021
R61335 vdd.n24832 vdd.n24830 0.021
R61336 vdd.n25238 vdd.n25236 0.021
R61337 vdd.n25226 vdd.n25224 0.021
R61338 vdd.n25214 vdd.n25212 0.021
R61339 vdd.n25202 vdd.n25200 0.021
R61340 vdd.n25190 vdd.n25188 0.021
R61341 vdd.n25178 vdd.n25176 0.021
R61342 vdd.n25160 vdd.n25152 0.021
R61343 vdd.n25135 vdd.n25127 0.021
R61344 vdd.n25123 vdd.n25115 0.021
R61345 vdd.n25111 vdd.n25103 0.021
R61346 vdd.n24927 vdd.n24926 0.021
R61347 vdd.n1172 vdd.n1046 0.021
R61348 vdd.n25532 vdd.n25531 0.021
R61349 vdd.n2334 vdd.n2109 0.021
R61350 vdd.n3859 vdd.n3829 0.021
R61351 vdd.n5186 vdd.n5185 0.021
R61352 vdd.n10168 vdd.n10167 0.021
R61353 vdd.n16769 vdd.n16768 0.021
R61354 vdd.n29162 vdd.n29160 0.021
R61355 vdd.n30933 vdd.n30932 0.021
R61356 vdd.n30890 vdd.n30889 0.021
R61357 vdd.n30867 vdd.n30866 0.021
R61358 vdd.n30001 vdd.n30000 0.021
R61359 vdd.n29586 vdd.n29585 0.021
R61360 vdd.n29584 vdd.n29583 0.021
R61361 vdd.n29471 vdd.n29470 0.021
R61362 vdd.n29388 vdd.n29387 0.021
R61363 vdd.n29386 vdd.n29385 0.021
R61364 vdd.n29344 vdd.n29343 0.021
R61365 vdd.n29342 vdd.n29341 0.021
R61366 vdd.n29213 vdd.n29212 0.021
R61367 vdd.n29109 vdd.n29108 0.021
R61368 vdd.n29107 vdd.n29106 0.021
R61369 vdd.n27722 vdd.n27721 0.021
R61370 vdd.n26436 vdd.n26435 0.021
R61371 vdd.n26247 vdd.n26246 0.021
R61372 vdd.n25352 vdd.n25351 0.021
R61373 vdd.n25350 vdd.n25349 0.021
R61374 vdd.n31345 vdd.n31344 0.021
R61375 vdd.n31343 vdd.n31342 0.021
R61376 vdd.n31398 vdd.n31397 0.021
R61377 vdd.n31396 vdd.n31395 0.021
R61378 vdd.n30913 vdd.n30912 0.021
R61379 vdd.n30911 vdd.n30910 0.021
R61380 vdd.n30718 vdd.n30717 0.021
R61381 vdd.n30716 vdd.n30715 0.021
R61382 vdd.n30171 vdd.n30170 0.021
R61383 vdd.n30169 vdd.n30168 0.021
R61384 vdd.n32591 vdd.n32590 0.021
R61385 vdd.n32589 vdd.n32588 0.021
R61386 vdd.n30153 vdd.n30152 0.021
R61387 vdd.n30151 vdd.n30150 0.021
R61388 vdd.n30066 vdd.n30065 0.021
R61389 vdd.n30064 vdd.n30063 0.021
R61390 vdd.n30033 vdd.n30032 0.021
R61391 vdd.n30031 vdd.n30030 0.021
R61392 vdd.n32632 vdd.n32631 0.021
R61393 vdd.n32630 vdd.n32629 0.021
R61394 vdd.n32729 vdd.n32728 0.021
R61395 vdd.n32727 vdd.n32726 0.021
R61396 vdd.n29608 vdd.n29607 0.021
R61397 vdd.n29606 vdd.n29605 0.021
R61398 vdd.n29559 vdd.n29558 0.021
R61399 vdd.n29557 vdd.n29556 0.021
R61400 vdd.n29490 vdd.n29489 0.021
R61401 vdd.n29488 vdd.n29487 0.021
R61402 vdd.n29404 vdd.n29403 0.021
R61403 vdd.n29402 vdd.n29401 0.021
R61404 vdd.n29365 vdd.n29364 0.021
R61405 vdd.n29363 vdd.n29362 0.021
R61406 vdd.n29265 vdd.n29264 0.021
R61407 vdd.n29263 vdd.n29262 0.021
R61408 vdd.n29247 vdd.n29246 0.021
R61409 vdd.n29245 vdd.n29244 0.021
R61410 vdd.n29143 vdd.n29142 0.021
R61411 vdd.n29141 vdd.n29140 0.021
R61412 vdd.n27742 vdd.n27741 0.021
R61413 vdd.n27740 vdd.n27739 0.021
R61414 vdd.n27702 vdd.n27701 0.021
R61415 vdd.n27700 vdd.n27699 0.021
R61416 vdd.n26532 vdd.n26531 0.021
R61417 vdd.n26530 vdd.n26529 0.021
R61418 vdd.n26556 vdd.n26555 0.021
R61419 vdd.n26554 vdd.n26553 0.021
R61420 vdd.n26265 vdd.n26264 0.021
R61421 vdd.n26263 vdd.n26262 0.021
R61422 vdd.n26576 vdd.n26575 0.021
R61423 vdd.n26574 vdd.n26573 0.021
R61424 vdd.n26224 vdd.n26223 0.021
R61425 vdd.n26222 vdd.n26221 0.021
R61426 vdd.n26090 vdd.n26089 0.021
R61427 vdd.n30940 vdd.n30939 0.021
R61428 vdd.n31369 vdd.n31368 0.021
R61429 vdd.n30837 vdd.n30835 0.021
R61430 vdd.n32541 vdd.n32539 0.021
R61431 vdd.n32544 vdd.n32542 0.021
R61432 vdd.n30110 vdd.n30109 0.021
R61433 vdd.n30112 vdd.n30111 0.021
R61434 vdd.n30046 vdd.n30045 0.021
R61435 vdd.n29979 vdd.n29977 0.021
R61436 vdd.n29648 vdd.n29647 0.021
R61437 vdd.n29651 vdd.n29649 0.021
R61438 vdd.n32683 vdd.n32682 0.021
R61439 vdd.n32685 vdd.n32684 0.021
R61440 vdd.n32716 vdd.n32715 0.021
R61441 vdd.n29537 vdd.n29536 0.021
R61442 vdd.n29442 vdd.n29440 0.021
R61443 vdd.n29445 vdd.n29443 0.021
R61444 vdd.n29317 vdd.n29316 0.021
R61445 vdd.n29319 vdd.n29318 0.021
R61446 vdd.n29257 vdd.n29256 0.021
R61447 vdd.n29189 vdd.n29188 0.021
R61448 vdd.n29234 vdd.n29233 0.021
R61449 vdd.n29159 vdd.n29158 0.021
R61450 vdd.n29123 vdd.n29122 0.021
R61451 vdd.n29049 vdd.n29048 0.021
R61452 vdd.n27729 vdd.n27728 0.021
R61453 vdd.n26484 vdd.n26481 0.021
R61454 vdd.n26428 vdd.n26426 0.021
R61455 vdd.n26358 vdd.n26356 0.021
R61456 vdd.n26361 vdd.n26359 0.021
R61457 vdd.n26627 vdd.n26626 0.021
R61458 vdd.n26629 vdd.n26628 0.021
R61459 vdd.n26112 vdd.n26111 0.021
R61460 vdd.n31318 vdd.n31317 0.021
R61461 vdd.n30973 vdd.n30971 0.021
R61462 vdd.n30841 vdd.n30839 0.021
R61463 vdd.n30846 vdd.n30844 0.021
R61464 vdd.n32549 vdd.n32547 0.021
R61465 vdd.n30048 vdd.n30047 0.021
R61466 vdd.n30050 vdd.n30049 0.021
R61467 vdd.n29984 vdd.n29982 0.021
R61468 vdd.n29657 vdd.n29655 0.021
R61469 vdd.n7159 vdd.n7158 0.021
R61470 vdd.n29540 vdd.n29539 0.021
R61471 vdd.n29450 vdd.n29448 0.021
R61472 vdd.n29232 vdd.n29231 0.021
R61473 vdd.n29193 vdd.n29192 0.021
R61474 vdd.n29230 vdd.n29229 0.021
R61475 vdd.n29125 vdd.n29124 0.021
R61476 vdd.n29127 vdd.n29126 0.021
R61477 vdd.n26488 vdd.n26487 0.021
R61478 vdd.n26366 vdd.n26364 0.021
R61479 vdd.n26110 vdd.n26109 0.021
R61480 vdd.n25365 vdd.n25363 0.021
R61481 vdd.n25674 vdd.n25671 0.021
R61482 vdd.n30826 vdd.n30825 0.021
R61483 vdd.n30849 vdd.n30847 0.021
R61484 vdd.n31424 vdd.n31423 0.021
R61485 vdd.n32552 vdd.n32550 0.021
R61486 vdd.n30099 vdd.n30098 0.021
R61487 vdd.n30053 vdd.n30052 0.021
R61488 vdd.n30055 vdd.n30054 0.021
R61489 vdd.n30117 vdd.n30116 0.021
R61490 vdd.n29660 vdd.n29658 0.021
R61491 vdd.n32674 vdd.n32673 0.021
R61492 vdd.n32689 vdd.n32688 0.021
R61493 vdd.n32693 vdd.n32692 0.021
R61494 vdd.n29510 vdd.n29509 0.021
R61495 vdd.n29547 vdd.n29546 0.021
R61496 vdd.n7164 vdd.n7163 0.021
R61497 vdd.n29428 vdd.n29427 0.021
R61498 vdd.n29453 vdd.n29451 0.021
R61499 vdd.n29306 vdd.n29305 0.021
R61500 vdd.n29323 vdd.n29322 0.021
R61501 vdd.n29326 vdd.n29325 0.021
R61502 vdd.n29226 vdd.n29225 0.021
R61503 vdd.n29224 vdd.n29223 0.021
R61504 vdd.n29198 vdd.n29196 0.021
R61505 vdd.n29130 vdd.n29129 0.021
R61506 vdd.n29132 vdd.n29131 0.021
R61507 vdd.n29074 vdd.n29073 0.021
R61508 vdd.n29053 vdd.n29052 0.021
R61509 vdd.n26464 vdd.n26463 0.021
R61510 vdd.n26496 vdd.n26495 0.021
R61511 vdd.n26498 vdd.n26497 0.021
R61512 vdd.n26383 vdd.n26382 0.021
R61513 vdd.n26282 vdd.n26281 0.021
R61514 vdd.n26369 vdd.n26367 0.021
R61515 vdd.n26648 vdd.n26647 0.021
R61516 vdd.n26102 vdd.n26101 0.021
R61517 vdd.n26100 vdd.n26099 0.021
R61518 vdd.n26634 vdd.n26633 0.021
R61519 vdd.n30802 vdd.n30801 0.021
R61520 vdd.n30852 vdd.n30851 0.021
R61521 vdd.n30854 vdd.n30853 0.021
R61522 vdd.n32555 vdd.n32554 0.021
R61523 vdd.n32557 vdd.n32556 0.021
R61524 vdd.n31422 vdd.n31421 0.021
R61525 vdd.n30119 vdd.n30118 0.021
R61526 vdd.n30121 vdd.n30120 0.021
R61527 vdd.n29988 vdd.n29987 0.021
R61528 vdd.n29990 vdd.n29989 0.021
R61529 vdd.n29663 vdd.n29662 0.021
R61530 vdd.n29665 vdd.n29664 0.021
R61531 vdd.n32696 vdd.n32695 0.021
R61532 vdd.n32698 vdd.n32697 0.021
R61533 vdd.n32661 vdd.n32660 0.021
R61534 vdd.n32672 vdd.n32671 0.021
R61535 vdd.n29526 vdd.n29525 0.021
R61536 vdd.n7167 vdd.n7166 0.021
R61537 vdd.n29456 vdd.n29455 0.021
R61538 vdd.n29458 vdd.n29457 0.021
R61539 vdd.n29426 vdd.n29425 0.021
R61540 vdd.n29329 vdd.n29328 0.021
R61541 vdd.n29331 vdd.n29330 0.021
R61542 vdd.n29200 vdd.n29199 0.021
R61543 vdd.n29202 vdd.n29201 0.021
R61544 vdd.n29153 vdd.n29152 0.021
R61545 vdd.n29151 vdd.n29150 0.021
R61546 vdd.n29058 vdd.n29057 0.021
R61547 vdd.n29060 vdd.n29059 0.021
R61548 vdd.n29082 vdd.n29081 0.021
R61549 vdd.n29072 vdd.n29071 0.021
R61550 vdd.n26447 vdd.n26446 0.021
R61551 vdd.n26507 vdd.n26506 0.021
R61552 vdd.n26493 vdd.n26492 0.021
R61553 vdd.n26372 vdd.n26371 0.021
R61554 vdd.n26374 vdd.n26373 0.021
R61555 vdd.n26280 vdd.n26279 0.021
R61556 vdd.n26636 vdd.n26635 0.021
R61557 vdd.n26638 vdd.n26637 0.021
R61558 vdd.n26142 vdd.n26141 0.021
R61559 vdd.n26104 vdd.n26103 0.021
R61560 vdd.n30765 vdd.n30763 0.021
R61561 vdd.n30829 vdd.n30827 0.021
R61562 vdd.n30812 vdd.n30804 0.021
R61563 vdd.n30858 vdd.n30857 0.021
R61564 vdd.n32561 vdd.n32560 0.021
R61565 vdd.n30102 vdd.n30100 0.021
R61566 vdd.n30058 vdd.n30056 0.021
R61567 vdd.n30123 vdd.n30122 0.021
R61568 vdd.n29994 vdd.n29993 0.021
R61569 vdd.n29669 vdd.n29668 0.021
R61570 vdd.n32701 vdd.n32700 0.021
R61571 vdd.n29512 vdd.n29511 0.021
R61572 vdd.n29550 vdd.n29548 0.021
R61573 vdd.n29528 vdd.n29527 0.021
R61574 vdd.n7171 vdd.n7170 0.021
R61575 vdd.n29462 vdd.n29461 0.021
R61576 vdd.n29309 vdd.n29307 0.021
R61577 vdd.n29334 vdd.n29333 0.021
R61578 vdd.n29222 vdd.n29220 0.021
R61579 vdd.n29204 vdd.n29203 0.021
R61580 vdd.n29149 vdd.n29148 0.021
R61581 vdd.n29135 vdd.n29133 0.021
R61582 vdd.n29063 vdd.n29062 0.021
R61583 vdd.n26502 vdd.n26500 0.021
R61584 vdd.n26445 vdd.n26444 0.021
R61585 vdd.n26381 vdd.n26380 0.021
R61586 vdd.n26378 vdd.n26377 0.021
R61587 vdd.n26646 vdd.n26644 0.021
R61588 vdd.n26097 vdd.n26095 0.021
R61589 vdd.n26640 vdd.n26639 0.021
R61590 vdd.n26130 vdd.n26129 0.021
R61591 vdd.n26726 vdd.n26724 0.021
R61592 vdd.n30977 vdd.n30976 0.021
R61593 vdd.n31324 vdd.n31323 0.021
R61594 vdd.n26088 vdd.n26087 0.021
R61595 vdd.n29182 vdd.n29181 0.021
R61596 vdd.n29273 vdd.n29272 0.021
R61597 vdd.n29417 vdd.n29416 0.021
R61598 vdd.n29413 vdd.n29412 0.021
R61599 vdd.n32651 vdd.n32650 0.021
R61600 vdd.n32648 vdd.n32647 0.021
R61601 vdd.n32641 vdd.n32640 0.021
R61602 vdd.n29633 vdd.n29632 0.021
R61603 vdd.n29959 vdd.n29958 0.021
R61604 vdd.n30075 vdd.n30074 0.021
R61605 vdd.n31413 vdd.n31412 0.021
R61606 vdd.n31410 vdd.n31409 0.021
R61607 vdd.n30727 vdd.n30726 0.021
R61608 vdd.n30733 vdd.n30731 0.021
R61609 vdd.n31191 vdd.n31190 0.021
R61610 vdd.n29047 vdd.n29045 0.021
R61611 vdd.n29090 vdd.n29088 0.021
R61612 vdd.n29066 vdd.n29064 0.021
R61613 vdd.n26516 vdd.n26514 0.021
R61614 vdd.n26479 vdd.n26477 0.021
R61615 vdd.n26355 vdd.n26353 0.021
R61616 vdd.n26273 vdd.n26271 0.021
R61617 vdd.n26625 vdd.n26623 0.021
R61618 vdd.n26118 vdd.n26116 0.021
R61619 vdd.n26115 vdd.n26113 0.021
R61620 vdd.n26722 vdd.n26721 0.021
R61621 vdd.n29236 vdd.n29235 0.021
R61622 vdd.n30980 vdd.n30979 0.021
R61623 vdd.n30982 vdd.n30981 0.021
R61624 vdd.n31360 vdd.n31359 0.021
R61625 vdd.n31358 vdd.n31357 0.021
R61626 vdd.n30931 vdd.n30930 0.021
R61627 vdd.n30929 vdd.n30928 0.021
R61628 vdd.n30887 vdd.n30886 0.021
R61629 vdd.n30885 vdd.n30884 0.021
R61630 vdd.n30864 vdd.n30863 0.021
R61631 vdd.n30862 vdd.n30861 0.021
R61632 vdd.n32567 vdd.n32566 0.021
R61633 vdd.n32565 vdd.n32564 0.021
R61634 vdd.n32609 vdd.n32608 0.021
R61635 vdd.n32607 vdd.n32606 0.021
R61636 vdd.n30129 vdd.n30128 0.021
R61637 vdd.n30127 vdd.n30126 0.021
R61638 vdd.n29999 vdd.n29998 0.021
R61639 vdd.n29997 vdd.n29996 0.021
R61640 vdd.n29675 vdd.n29674 0.021
R61641 vdd.n29673 vdd.n29672 0.021
R61642 vdd.n32707 vdd.n32706 0.021
R61643 vdd.n32705 vdd.n32704 0.021
R61644 vdd.n29625 vdd.n29624 0.021
R61645 vdd.n29623 vdd.n29622 0.021
R61646 vdd.n29582 vdd.n29581 0.021
R61647 vdd.n29580 vdd.n29579 0.021
R61648 vdd.n7215 vdd.n7214 0.021
R61649 vdd.n29468 vdd.n29467 0.021
R61650 vdd.n29466 vdd.n29465 0.021
R61651 vdd.n29384 vdd.n29383 0.021
R61652 vdd.n29382 vdd.n29381 0.021
R61653 vdd.n29340 vdd.n29339 0.021
R61654 vdd.n29338 vdd.n29337 0.021
R61655 vdd.n29210 vdd.n29209 0.021
R61656 vdd.n29208 vdd.n29207 0.021
R61657 vdd.n29169 vdd.n29168 0.021
R61658 vdd.n29167 vdd.n29166 0.021
R61659 vdd.n29105 vdd.n29104 0.021
R61660 vdd.n29103 vdd.n29102 0.021
R61661 vdd.n27719 vdd.n27718 0.021
R61662 vdd.n27717 vdd.n27716 0.021
R61663 vdd.n27677 vdd.n27676 0.021
R61664 vdd.n27675 vdd.n27674 0.021
R61665 vdd.n26433 vdd.n26432 0.021
R61666 vdd.n26431 vdd.n26430 0.021
R61667 vdd.n26411 vdd.n26410 0.021
R61668 vdd.n26409 vdd.n26408 0.021
R61669 vdd.n26245 vdd.n26244 0.021
R61670 vdd.n26243 vdd.n26242 0.021
R61671 vdd.n26715 vdd.n26714 0.021
R61672 vdd.n26713 vdd.n26712 0.021
R61673 vdd.n25348 vdd.n25347 0.021
R61674 vdd.n25346 vdd.n25345 0.021
R61675 vdd.n31339 vdd.n31338 0.021
R61676 vdd.n31394 vdd.n31393 0.021
R61677 vdd.n30909 vdd.n30908 0.021
R61678 vdd.n30907 vdd.n30906 0.021
R61679 vdd.n30713 vdd.n30712 0.021
R61680 vdd.n30166 vdd.n30165 0.021
R61681 vdd.n32587 vdd.n32586 0.021
R61682 vdd.n32585 vdd.n32584 0.021
R61683 vdd.n30149 vdd.n30148 0.021
R61684 vdd.n30147 vdd.n30146 0.021
R61685 vdd.n30062 vdd.n30061 0.021
R61686 vdd.n30029 vdd.n30028 0.021
R61687 vdd.n30027 vdd.n30026 0.021
R61688 vdd.n32628 vdd.n32627 0.021
R61689 vdd.n32626 vdd.n32625 0.021
R61690 vdd.n32725 vdd.n32724 0.021
R61691 vdd.n32723 vdd.n32722 0.021
R61692 vdd.n29604 vdd.n29603 0.021
R61693 vdd.n29554 vdd.n29553 0.021
R61694 vdd.n29486 vdd.n29485 0.021
R61695 vdd.n29484 vdd.n29483 0.021
R61696 vdd.n29260 vdd.n29259 0.021
R61697 vdd.n29242 vdd.n29241 0.021
R61698 vdd.n29139 vdd.n29138 0.021
R61699 vdd.n27737 vdd.n27736 0.021
R61700 vdd.n27697 vdd.n27696 0.021
R61701 vdd.n26528 vdd.n26527 0.021
R61702 vdd.n26526 vdd.n26525 0.021
R61703 vdd.n26551 vdd.n26550 0.021
R61704 vdd.n26261 vdd.n26260 0.021
R61705 vdd.n26572 vdd.n26571 0.021
R61706 vdd.n26570 vdd.n26569 0.021
R61707 vdd.n26220 vdd.n26219 0.021
R61708 vdd.n26085 vdd.n26084 0.021
R61709 vdd.n31341 vdd.n31340 0.021
R61710 vdd.n4151 vdd.n4150 0.021
R61711 vdd.n4386 vdd.n4385 0.021
R61712 vdd.n4513 vdd.n4512 0.021
R61713 vdd.n5320 vdd.n5319 0.021
R61714 vdd.n5560 vdd.n5559 0.021
R61715 vdd.n5686 vdd.n5685 0.021
R61716 vdd.n6284 vdd.n6283 0.021
R61717 vdd.n6106 vdd.n6105 0.021
R61718 vdd.n5982 vdd.n5981 0.021
R61719 vdd.n34573 vdd.n34572 0.021
R61720 vdd.n34813 vdd.n34812 0.021
R61721 vdd.n34939 vdd.n34938 0.021
R61722 vdd.n35155 vdd.n35154 0.021
R61723 vdd.n35409 vdd.n35408 0.021
R61724 vdd.n35524 vdd.n35523 0.021
R61725 vdd.n33993 vdd.n33992 0.021
R61726 vdd.n34393 vdd.n34392 0.021
R61727 vdd.n34258 vdd.n34257 0.021
R61728 vdd.n6137 vdd.n6045 0.02
R61729 vdd.n30697 vdd.n30693 0.02
R61730 vdd.n11787 vdd.n11786 0.02
R61731 vdd.n21752 vdd.n21751 0.02
R61732 vdd.n35355 vdd.n35354 0.02
R61733 vdd.n34771 vdd.n34770 0.02
R61734 vdd.n5518 vdd.n5517 0.02
R61735 vdd.n4345 vdd.n4344 0.02
R61736 vdd.n33570 vdd.n33569 0.02
R61737 vdd.n27457 vdd.n27456 0.02
R61738 vdd.n25903 vdd.n25902 0.02
R61739 vdd.n4951 vdd.n4871 0.02
R61740 vdd.n4602 vdd.n4448 0.02
R61741 vdd.n35233 vdd.n35232 0.02
R61742 vdd.n34646 vdd.n34645 0.02
R61743 vdd.n5393 vdd.n5392 0.02
R61744 vdd.n4711 vdd.n4710 0.02
R61745 vdd.n4223 vdd.n4222 0.02
R61746 vdd.n33336 vdd.n33335 0.02
R61747 vdd.n33564 vdd.n33563 0.02
R61748 vdd.n33594 vdd.n33593 0.02
R61749 vdd.n35568 vdd.n35567 0.02
R61750 vdd.n35516 vdd.n35504 0.02
R61751 vdd.n35437 vdd.n35436 0.02
R61752 vdd.n35463 vdd.n35460 0.02
R61753 vdd.n35329 vdd.n35328 0.02
R61754 vdd.n554 vdd.n553 0.02
R61755 vdd.n56 vdd.n55 0.02
R61756 vdd.n61 vdd.n60 0.02
R61757 vdd.n95 vdd.n94 0.02
R61758 vdd.n93 vdd.n91 0.02
R61759 vdd.n159 vdd.n158 0.02
R61760 vdd.n294 vdd.n293 0.02
R61761 vdd.n6023 vdd.n6022 0.02
R61762 vdd.n6006 vdd.n6005 0.02
R61763 vdd.n6117 vdd.n6116 0.02
R61764 vdd.n6134 vdd.n6133 0.02
R61765 vdd.n5898 vdd.n5897 0.02
R61766 vdd.n4741 vdd.n4740 0.02
R61767 vdd.n5059 vdd.n5058 0.02
R61768 vdd.n4507 vdd.n4506 0.02
R61769 vdd.n4234 vdd.n4233 0.02
R61770 vdd.n4284 vdd.n4283 0.02
R61771 vdd.n4116 vdd.n4115 0.02
R61772 vdd.n4412 vdd.n4411 0.02
R61773 vdd.n26318 vdd.n26297 0.02
R61774 vdd.n32166 vdd.n32165 0.02
R61775 vdd.n10219 vdd.n10218 0.02
R61776 vdd.n10202 vdd.n10201 0.02
R61777 vdd.n11695 vdd.n11682 0.02
R61778 vdd.n11869 vdd.n11868 0.02
R61779 vdd.n24178 vdd.n24176 0.02
R61780 vdd.n23998 vdd.n23996 0.02
R61781 vdd.n23946 vdd.n23944 0.02
R61782 vdd.n23766 vdd.n23764 0.02
R61783 vdd.n23714 vdd.n23712 0.02
R61784 vdd.n23078 vdd.n23076 0.02
R61785 vdd.n23258 vdd.n23256 0.02
R61786 vdd.n23310 vdd.n23308 0.02
R61787 vdd.n23490 vdd.n23488 0.02
R61788 vdd.n23542 vdd.n23540 0.02
R61789 vdd.n22499 vdd.n22497 0.02
R61790 vdd.n22679 vdd.n22677 0.02
R61791 vdd.n22731 vdd.n22729 0.02
R61792 vdd.n22911 vdd.n22909 0.02
R61793 vdd.n22963 vdd.n22961 0.02
R61794 vdd.n16591 vdd.n16590 0.02
R61795 vdd.n16695 vdd.n16694 0.02
R61796 vdd.n21798 vdd.n21797 0.02
R61797 vdd.n21960 vdd.n21959 0.02
R61798 vdd.n24998 vdd.n24996 0.02
R61799 vdd.n24945 vdd.n24944 0.02
R61800 vdd.n24563 vdd.n24562 0.02
R61801 vdd.n35025 vdd.n34874 0.02
R61802 vdd.n5772 vdd.n5621 0.02
R61803 vdd.n29506 vdd.n29505 0.02
R61804 vdd.n880 vdd.n879 0.02
R61805 vdd.n26213 vdd.n26184 0.02
R61806 vdd.n35611 vdd.n35610 0.02
R61807 vdd.n33367 vdd.n33366 0.02
R61808 vdd.n33698 vdd.n33697 0.02
R61809 vdd.n33789 vdd.n33782 0.02
R61810 vdd.n577 vdd.n576 0.02
R61811 vdd.n6350 vdd.n6347 0.02
R61812 vdd.n33474 vdd.n33391 0.02
R61813 vdd.n787 vdd.n705 0.02
R61814 vdd.n1170 vdd.n1169 0.02
R61815 vdd.n35024 vdd.n35023 0.019
R61816 vdd.n5771 vdd.n5770 0.019
R61817 vdd.n4601 vdd.n4600 0.019
R61818 vdd.n784 vdd.n781 0.019
R61819 vdd.n30699 vdd.n30692 0.019
R61820 vdd.n27884 vdd.n27873 0.019
R61821 vdd.n26061 vdd.n26059 0.019
R61822 vdd.n25964 vdd.n25963 0.019
R61823 vdd.n32811 vdd.n32810 0.019
R61824 vdd.n32806 vdd.n32805 0.019
R61825 vdd.n32801 vdd.n32800 0.019
R61826 vdd.n32798 vdd.n32797 0.019
R61827 vdd.n32795 vdd.n32794 0.019
R61828 vdd.n32792 vdd.n32791 0.019
R61829 vdd.n32787 vdd.n32786 0.019
R61830 vdd.n32784 vdd.n32783 0.019
R61831 vdd.n32777 vdd.n32776 0.019
R61832 vdd.n32774 vdd.n32773 0.019
R61833 vdd.n32771 vdd.n32770 0.019
R61834 vdd.n32768 vdd.n32767 0.019
R61835 vdd.n32765 vdd.n32764 0.019
R61836 vdd.n32762 vdd.n32761 0.019
R61837 vdd.n32759 vdd.n32758 0.019
R61838 vdd.n32756 vdd.n32755 0.019
R61839 vdd.n32753 vdd.n32752 0.019
R61840 vdd.n32750 vdd.n32749 0.019
R61841 vdd.n32747 vdd.n32746 0.019
R61842 vdd.n32744 vdd.n32743 0.019
R61843 vdd.n32741 vdd.n32740 0.019
R61844 vdd.n25334 vdd.n25333 0.019
R61845 vdd.n25331 vdd.n25330 0.019
R61846 vdd.n25328 vdd.n25327 0.019
R61847 vdd.n25325 vdd.n25324 0.019
R61848 vdd.n25322 vdd.n25321 0.019
R61849 vdd.n25317 vdd.n25316 0.019
R61850 vdd.n25314 vdd.n25313 0.019
R61851 vdd.n25311 vdd.n25310 0.019
R61852 vdd.n25308 vdd.n25307 0.019
R61853 vdd.n25305 vdd.n25304 0.019
R61854 vdd.n25300 vdd.n25299 0.019
R61855 vdd.n25295 vdd.n25294 0.019
R61856 vdd.n25290 vdd.n25289 0.019
R61857 vdd.n25283 vdd.n25282 0.019
R61858 vdd.n25280 vdd.n25279 0.019
R61859 vdd.n25277 vdd.n25276 0.019
R61860 vdd.n25274 vdd.n25273 0.019
R61861 vdd.n25271 vdd.n25270 0.019
R61862 vdd.n25268 vdd.n25267 0.019
R61863 vdd.n29863 vdd.n29862 0.019
R61864 vdd.n25478 vdd.n25475 0.019
R61865 vdd.n25949 vdd.n25947 0.019
R61866 vdd.n25867 vdd.n25866 0.019
R61867 vdd.n6918 vdd.n6917 0.019
R61868 vdd.n6949 vdd.n6948 0.019
R61869 vdd.n6975 vdd.n6974 0.019
R61870 vdd.n7006 vdd.n7005 0.019
R61871 vdd.n7031 vdd.n7030 0.019
R61872 vdd.n7085 vdd.n7084 0.019
R61873 vdd.n7284 vdd.n7283 0.019
R61874 vdd.n7824 vdd.n7823 0.019
R61875 vdd.n7850 vdd.n7849 0.019
R61876 vdd.n7881 vdd.n7880 0.019
R61877 vdd.n7907 vdd.n7906 0.019
R61878 vdd.n7935 vdd.n7934 0.019
R61879 vdd.n6779 vdd.n6778 0.019
R61880 vdd.n6719 vdd.n6718 0.019
R61881 vdd.n6667 vdd.n6666 0.019
R61882 vdd.n6554 vdd.n6553 0.019
R61883 vdd.n6496 vdd.n6495 0.019
R61884 vdd.n6439 vdd.n6438 0.019
R61885 vdd.n6373 vdd.n6365 0.019
R61886 vdd.n26706 vdd.n26687 0.019
R61887 vdd.n25874 vdd.n25873 0.019
R61888 vdd.n25760 vdd.n25759 0.019
R61889 vdd.n26064 vdd.n26062 0.019
R61890 vdd.n25957 vdd.n25956 0.019
R61891 vdd.n25955 vdd.n25953 0.019
R61892 vdd.n25860 vdd.n25859 0.019
R61893 vdd.n2765 vdd.n2763 0.019
R61894 vdd.n2837 vdd.n2835 0.019
R61895 vdd.n2946 vdd.n2944 0.019
R61896 vdd.n3018 vdd.n3016 0.019
R61897 vdd.n3127 vdd.n3125 0.019
R61898 vdd.n3199 vdd.n3197 0.019
R61899 vdd.n3308 vdd.n3306 0.019
R61900 vdd.n3380 vdd.n3378 0.019
R61901 vdd.n3489 vdd.n3487 0.019
R61902 vdd.n3561 vdd.n3559 0.019
R61903 vdd.n34313 vdd.n34312 0.019
R61904 vdd.n34252 vdd.n34251 0.019
R61905 vdd.n34152 vdd.n34151 0.019
R61906 vdd.n34260 vdd.n34259 0.019
R61907 vdd.n34154 vdd.n34153 0.019
R61908 vdd.n34184 vdd.n34183 0.019
R61909 vdd.n34195 vdd.n34194 0.019
R61910 vdd.n33965 vdd.n33865 0.019
R61911 vdd.n34398 vdd.n34397 0.019
R61912 vdd.n33965 vdd.n33964 0.019
R61913 vdd.n34411 vdd.n34410 0.019
R61914 vdd.n34933 vdd.n34932 0.019
R61915 vdd.n34657 vdd.n34656 0.019
R61916 vdd.n35002 vdd.n35001 0.019
R61917 vdd.n34985 vdd.n34984 0.019
R61918 vdd.n34690 vdd.n34689 0.019
R61919 vdd.n34710 vdd.n34709 0.019
R61920 vdd.n34743 vdd.n34742 0.019
R61921 vdd.n34539 vdd.n34529 0.019
R61922 vdd.n34836 vdd.n34835 0.019
R61923 vdd.n34539 vdd.n34538 0.019
R61924 vdd.n34838 vdd.n34837 0.019
R61925 vdd.n756 vdd.n755 0.019
R61926 vdd.n616 vdd.n615 0.019
R61927 vdd.n1043 vdd.n981 0.019
R61928 vdd.n665 vdd.n664 0.019
R61929 vdd.n1020 vdd.n1019 0.019
R61930 vdd.n1043 vdd.n1042 0.019
R61931 vdd.n1119 vdd.n1116 0.019
R61932 vdd.n1119 vdd.n1118 0.019
R61933 vdd.n5680 vdd.n5679 0.019
R61934 vdd.n5404 vdd.n5403 0.019
R61935 vdd.n5749 vdd.n5748 0.019
R61936 vdd.n5732 vdd.n5731 0.019
R61937 vdd.n5437 vdd.n5436 0.019
R61938 vdd.n5457 vdd.n5456 0.019
R61939 vdd.n5490 vdd.n5489 0.019
R61940 vdd.n5286 vdd.n5276 0.019
R61941 vdd.n5583 vdd.n5582 0.019
R61942 vdd.n5286 vdd.n5285 0.019
R61943 vdd.n5585 vdd.n5584 0.019
R61944 vdd.n35876 vdd.n35874 0.019
R61945 vdd.n35967 vdd.n35965 0.019
R61946 vdd.n36107 vdd.n36105 0.019
R61947 vdd.n36198 vdd.n36196 0.019
R61948 vdd.n36338 vdd.n36336 0.019
R61949 vdd.n36429 vdd.n36427 0.019
R61950 vdd.n36569 vdd.n36567 0.019
R61951 vdd.n36660 vdd.n36658 0.019
R61952 vdd.n36800 vdd.n36798 0.019
R61953 vdd.n36891 vdd.n36889 0.019
R61954 vdd.n38086 vdd.n38084 0.019
R61955 vdd.n37946 vdd.n37944 0.019
R61956 vdd.n37855 vdd.n37853 0.019
R61957 vdd.n37715 vdd.n37713 0.019
R61958 vdd.n37624 vdd.n37622 0.019
R61959 vdd.n28297 vdd.n28295 0.019
R61960 vdd.n28388 vdd.n28386 0.019
R61961 vdd.n28528 vdd.n28526 0.019
R61962 vdd.n28619 vdd.n28617 0.019
R61963 vdd.n28759 vdd.n28757 0.019
R61964 vdd.n1708 vdd.n1706 0.019
R61965 vdd.n1599 vdd.n1597 0.019
R61966 vdd.n1527 vdd.n1525 0.019
R61967 vdd.n1418 vdd.n1416 0.019
R61968 vdd.n1346 vdd.n1344 0.019
R61969 vdd.n26812 vdd.n26810 0.019
R61970 vdd.n26884 vdd.n26882 0.019
R61971 vdd.n26993 vdd.n26991 0.019
R61972 vdd.n27065 vdd.n27063 0.019
R61973 vdd.n27174 vdd.n27172 0.019
R61974 vdd.n31389 vdd.n31387 0.019
R61975 vdd.n31389 vdd.n31388 0.019
R61976 vdd.n30161 vdd.n30160 0.019
R61977 vdd.n30163 vdd.n30162 0.019
R61978 vdd.n32719 vdd.n32718 0.019
R61979 vdd.n2387 vdd.n2371 0.019
R61980 vdd.n1957 vdd.n1956 0.019
R61981 vdd.n32480 vdd.n32479 0.019
R61982 vdd.n10199 vdd.n10078 0.019
R61983 vdd.n11488 vdd.n11467 0.019
R61984 vdd.n11532 vdd.n11455 0.019
R61985 vdd.n11953 vdd.n11450 0.019
R61986 vdd.n11514 vdd.n11511 0.019
R61987 vdd.n11456 vdd.n11452 0.019
R61988 vdd.n11952 vdd.n11951 0.019
R61989 vdd.n11898 vdd.n11793 0.019
R61990 vdd.n11827 vdd.n11816 0.019
R61991 vdd.n11867 vdd.n11807 0.019
R61992 vdd.n24118 vdd.n24108 0.019
R61993 vdd.n24066 vdd.n24064 0.019
R61994 vdd.n23886 vdd.n23876 0.019
R61995 vdd.n23834 vdd.n23832 0.019
R61996 vdd.n23654 vdd.n23644 0.019
R61997 vdd.n23146 vdd.n23144 0.019
R61998 vdd.n23198 vdd.n23188 0.019
R61999 vdd.n23378 vdd.n23376 0.019
R62000 vdd.n23430 vdd.n23420 0.019
R62001 vdd.n23610 vdd.n23608 0.019
R62002 vdd.n22567 vdd.n22565 0.019
R62003 vdd.n22619 vdd.n22609 0.019
R62004 vdd.n22799 vdd.n22797 0.019
R62005 vdd.n22851 vdd.n22841 0.019
R62006 vdd.n23031 vdd.n23029 0.019
R62007 vdd.n18311 vdd.n18310 0.019
R62008 vdd.n18369 vdd.n18358 0.019
R62009 vdd.n18382 vdd.n18378 0.019
R62010 vdd.n18420 vdd.n18419 0.019
R62011 vdd.n18424 vdd.n18423 0.019
R62012 vdd.n21989 vdd.n21884 0.019
R62013 vdd.n21918 vdd.n21907 0.019
R62014 vdd.n21958 vdd.n21898 0.019
R62015 vdd.n24881 vdd.n24880 0.019
R62016 vdd.n5048 vdd.n5047 0.019
R62017 vdd.n32034 vdd.n32032 0.019
R62018 vdd.n26337 vdd.n26323 0.019
R62019 vdd.n34340 vdd.n34339 0.019
R62020 vdd.n3873 vdd.n3867 0.019
R62021 vdd.n2501 vdd.n2446 0.019
R62022 vdd.n35227 vdd.n35224 0.019
R62023 vdd.n34640 vdd.n34637 0.019
R62024 vdd.n5387 vdd.n5384 0.019
R62025 vdd.n4217 vdd.n4214 0.019
R62026 vdd.n26054 vdd.n26052 0.019
R62027 vdd.n2514 vdd.n2435 0.019
R62028 vdd.n1854 vdd.n1853 0.019
R62029 vdd.n6468 vdd.n6467 0.019
R62030 vdd.n6522 vdd.n6521 0.019
R62031 vdd.n6665 vdd.n6664 0.019
R62032 vdd.n6746 vdd.n6745 0.019
R62033 vdd.n6777 vdd.n6776 0.019
R62034 vdd.n7255 vdd.n7254 0.019
R62035 vdd.n7424 vdd.n7423 0.019
R62036 vdd.n7594 vdd.n7593 0.019
R62037 vdd.n7651 vdd.n7650 0.019
R62038 vdd.n7708 vdd.n7707 0.019
R62039 vdd.n7763 vdd.n7762 0.019
R62040 vdd.n7792 vdd.n7791 0.019
R62041 vdd.n7980 vdd.n7979 0.019
R62042 vdd.n7898 vdd.n7897 0.019
R62043 vdd.n7784 vdd.n7783 0.019
R62044 vdd.n7727 vdd.n7726 0.019
R62045 vdd.n7670 vdd.n7669 0.019
R62046 vdd.n7613 vdd.n7612 0.019
R62047 vdd.n7497 vdd.n7496 0.019
R62048 vdd.n7494 vdd.n7493 0.019
R62049 vdd.n7444 vdd.n7443 0.019
R62050 vdd.n7387 vdd.n7386 0.019
R62051 vdd.n7328 vdd.n7327 0.019
R62052 vdd.n7276 vdd.n7275 0.019
R62053 vdd.n7273 vdd.n7272 0.019
R62054 vdd.n7140 vdd.n7139 0.019
R62055 vdd.n7107 vdd.n7106 0.019
R62056 vdd.n7050 vdd.n7049 0.019
R62057 vdd.n6937 vdd.n6936 0.019
R62058 vdd.n6882 vdd.n6881 0.019
R62059 vdd.n6826 vdd.n6825 0.019
R62060 vdd.n6765 vdd.n6764 0.019
R62061 vdd.n6708 vdd.n6707 0.019
R62062 vdd.n6655 vdd.n6654 0.019
R62063 vdd.n6597 vdd.n6596 0.019
R62064 vdd.n6543 vdd.n6542 0.019
R62065 vdd.n6484 vdd.n6483 0.019
R62066 vdd.n7929 vdd.n7928 0.019
R62067 vdd.n7874 vdd.n7873 0.019
R62068 vdd.n7817 vdd.n7816 0.019
R62069 vdd.n7757 vdd.n7756 0.019
R62070 vdd.n7702 vdd.n7701 0.019
R62071 vdd.n7645 vdd.n7644 0.019
R62072 vdd.n7588 vdd.n7587 0.019
R62073 vdd.n7531 vdd.n7530 0.019
R62074 vdd.n7418 vdd.n7417 0.019
R62075 vdd.n7362 vdd.n7361 0.019
R62076 vdd.n7306 vdd.n7305 0.019
R62077 vdd.n7249 vdd.n7248 0.019
R62078 vdd.n6690 vdd.n6689 0.019
R62079 vdd.n6632 vdd.n6631 0.019
R62080 vdd.n6397 vdd.n6396 0.019
R62081 vdd.n7924 vdd.n7923 0.019
R62082 vdd.n7868 vdd.n7867 0.019
R62083 vdd.n7812 vdd.n7811 0.019
R62084 vdd.n7752 vdd.n7751 0.019
R62085 vdd.n7697 vdd.n7696 0.019
R62086 vdd.n7640 vdd.n7639 0.019
R62087 vdd.n7582 vdd.n7581 0.019
R62088 vdd.n7526 vdd.n7525 0.019
R62089 vdd.n7413 vdd.n7412 0.019
R62090 vdd.n7356 vdd.n7355 0.019
R62091 vdd.n7302 vdd.n7301 0.019
R62092 vdd.n7244 vdd.n7243 0.019
R62093 vdd.n6686 vdd.n6685 0.019
R62094 vdd.n6626 vdd.n6625 0.019
R62095 vdd.n6458 vdd.n6457 0.019
R62096 vdd.n6390 vdd.n6388 0.019
R62097 vdd.n7974 vdd.n7972 0.019
R62098 vdd.n7954 vdd.n7953 0.019
R62099 vdd.n24927 vdd.n24921 0.019
R62100 vdd.n24931 vdd.n24918 0.019
R62101 vdd.n29036 vdd.n29035 0.019
R62102 vdd.n4949 vdd.n4948 0.019
R62103 vdd.n7926 vdd.n7925 0.019
R62104 vdd.n7872 vdd.n7871 0.019
R62105 vdd.n7870 vdd.n7869 0.019
R62106 vdd.n7814 vdd.n7813 0.019
R62107 vdd.n7754 vdd.n7753 0.019
R62108 vdd.n7699 vdd.n7698 0.019
R62109 vdd.n7642 vdd.n7641 0.019
R62110 vdd.n7586 vdd.n7585 0.019
R62111 vdd.n7584 vdd.n7583 0.019
R62112 vdd.n7528 vdd.n7527 0.019
R62113 vdd.n7415 vdd.n7414 0.019
R62114 vdd.n7360 vdd.n7359 0.019
R62115 vdd.n7358 vdd.n7357 0.019
R62116 vdd.n7247 vdd.n7246 0.019
R62117 vdd.n7077 vdd.n7076 0.019
R62118 vdd.n7025 vdd.n7024 0.019
R62119 vdd.n7023 vdd.n7022 0.019
R62120 vdd.n6969 vdd.n6968 0.019
R62121 vdd.n6967 vdd.n6966 0.019
R62122 vdd.n6854 vdd.n6853 0.019
R62123 vdd.n6801 vdd.n6800 0.019
R62124 vdd.n6799 vdd.n6798 0.019
R62125 vdd.n6739 vdd.n6738 0.019
R62126 vdd.n6629 vdd.n6628 0.019
R62127 vdd.n6572 vdd.n6571 0.019
R62128 vdd.n6515 vdd.n6514 0.019
R62129 vdd.n6462 vdd.n6461 0.019
R62130 vdd.n6460 vdd.n6459 0.019
R62131 vdd.n6393 vdd.n6392 0.019
R62132 vdd.n7901 vdd.n7900 0.019
R62133 vdd.n7877 vdd.n7876 0.019
R62134 vdd.n7844 vdd.n7843 0.019
R62135 vdd.n7820 vdd.n7819 0.019
R62136 vdd.n7787 vdd.n7786 0.019
R62137 vdd.n7760 vdd.n7759 0.019
R62138 vdd.n7730 vdd.n7729 0.019
R62139 vdd.n7705 vdd.n7704 0.019
R62140 vdd.n7673 vdd.n7672 0.019
R62141 vdd.n7648 vdd.n7647 0.019
R62142 vdd.n7616 vdd.n7615 0.019
R62143 vdd.n7591 vdd.n7590 0.019
R62144 vdd.n7558 vdd.n7557 0.019
R62145 vdd.n7534 vdd.n7533 0.019
R62146 vdd.n7501 vdd.n7500 0.019
R62147 vdd.n7499 vdd.n7498 0.019
R62148 vdd.n7447 vdd.n7446 0.019
R62149 vdd.n7421 vdd.n7420 0.019
R62150 vdd.n7390 vdd.n7389 0.019
R62151 vdd.n7364 vdd.n7363 0.019
R62152 vdd.n7366 vdd.n7365 0.019
R62153 vdd.n7308 vdd.n7307 0.019
R62154 vdd.n7310 vdd.n7309 0.019
R62155 vdd.n7251 vdd.n7250 0.019
R62156 vdd.n7253 vdd.n7252 0.019
R62157 vdd.n7149 vdd.n7148 0.019
R62158 vdd.n7143 vdd.n7142 0.019
R62159 vdd.n7082 vdd.n7081 0.019
R62160 vdd.n7054 vdd.n7053 0.019
R62161 vdd.n7052 vdd.n7051 0.019
R62162 vdd.n6998 vdd.n6997 0.019
R62163 vdd.n6996 vdd.n6995 0.019
R62164 vdd.n6941 vdd.n6940 0.019
R62165 vdd.n6913 vdd.n6912 0.019
R62166 vdd.n6915 vdd.n6914 0.019
R62167 vdd.n6859 vdd.n6858 0.019
R62168 vdd.n6829 vdd.n6828 0.019
R62169 vdd.n6805 vdd.n6804 0.019
R62170 vdd.n6770 vdd.n6769 0.019
R62171 vdd.n6742 vdd.n6741 0.019
R62172 vdd.n6768 vdd.n6767 0.019
R62173 vdd.n6712 vdd.n6711 0.019
R62174 vdd.n6659 vdd.n6658 0.019
R62175 vdd.n6657 vdd.n6656 0.019
R62176 vdd.n6600 vdd.n6599 0.019
R62177 vdd.n6577 vdd.n6576 0.019
R62178 vdd.n6546 vdd.n6545 0.019
R62179 vdd.n6520 vdd.n6519 0.019
R62180 vdd.n6488 vdd.n6487 0.019
R62181 vdd.n6486 vdd.n6485 0.019
R62182 vdd.n6433 vdd.n6432 0.019
R62183 vdd.n6395 vdd.n6394 0.019
R62184 vdd.n6431 vdd.n6430 0.019
R62185 vdd.n7904 vdd.n7903 0.019
R62186 vdd.n7847 vdd.n7846 0.019
R62187 vdd.n7790 vdd.n7789 0.019
R62188 vdd.n7733 vdd.n7732 0.019
R62189 vdd.n7676 vdd.n7675 0.019
R62190 vdd.n7619 vdd.n7618 0.019
R62191 vdd.n7561 vdd.n7560 0.019
R62192 vdd.n7503 vdd.n7502 0.019
R62193 vdd.n7505 vdd.n7504 0.019
R62194 vdd.n7450 vdd.n7449 0.019
R62195 vdd.n7393 vdd.n7392 0.019
R62196 vdd.n7335 vdd.n7334 0.019
R62197 vdd.n7281 vdd.n7280 0.019
R62198 vdd.n7225 vdd.n7224 0.019
R62199 vdd.n7147 vdd.n7146 0.019
R62200 vdd.n7111 vdd.n7110 0.019
R62201 vdd.n7113 vdd.n7112 0.019
R62202 vdd.n7057 vdd.n7056 0.019
R62203 vdd.n7059 vdd.n7058 0.019
R62204 vdd.n7001 vdd.n7000 0.019
R62205 vdd.n7003 vdd.n7002 0.019
R62206 vdd.n6944 vdd.n6943 0.019
R62207 vdd.n6946 vdd.n6945 0.019
R62208 vdd.n6887 vdd.n6886 0.019
R62209 vdd.n6889 vdd.n6888 0.019
R62210 vdd.n6832 vdd.n6831 0.019
R62211 vdd.n6834 vdd.n6833 0.019
R62212 vdd.n6773 vdd.n6772 0.019
R62213 vdd.n6775 vdd.n6774 0.019
R62214 vdd.n6716 vdd.n6715 0.019
R62215 vdd.n6663 vdd.n6662 0.019
R62216 vdd.n6602 vdd.n6601 0.019
R62217 vdd.n6604 vdd.n6603 0.019
R62218 vdd.n6549 vdd.n6548 0.019
R62219 vdd.n6551 vdd.n6550 0.019
R62220 vdd.n6491 vdd.n6490 0.019
R62221 vdd.n6493 vdd.n6492 0.019
R62222 vdd.n6436 vdd.n6435 0.019
R62223 vdd.n6399 vdd.n6398 0.019
R62224 vdd.n7960 vdd.n7959 0.019
R62225 vdd.n7922 vdd.n7921 0.019
R62226 vdd.n7866 vdd.n7865 0.019
R62227 vdd.n7810 vdd.n7809 0.019
R62228 vdd.n7750 vdd.n7749 0.019
R62229 vdd.n7695 vdd.n7694 0.019
R62230 vdd.n7638 vdd.n7637 0.019
R62231 vdd.n7580 vdd.n7579 0.019
R62232 vdd.n7524 vdd.n7523 0.019
R62233 vdd.n7467 vdd.n7466 0.019
R62234 vdd.n7492 vdd.n7491 0.019
R62235 vdd.n7411 vdd.n7410 0.019
R62236 vdd.n7354 vdd.n7353 0.019
R62237 vdd.n7300 vdd.n7299 0.019
R62238 vdd.n7242 vdd.n7241 0.019
R62239 vdd.n7136 vdd.n7135 0.019
R62240 vdd.n7073 vdd.n7072 0.019
R62241 vdd.n7103 vdd.n7102 0.019
R62242 vdd.n7019 vdd.n7018 0.019
R62243 vdd.n7047 vdd.n7046 0.019
R62244 vdd.n6963 vdd.n6962 0.019
R62245 vdd.n6992 vdd.n6991 0.019
R62246 vdd.n6906 vdd.n6905 0.019
R62247 vdd.n6935 vdd.n6934 0.019
R62248 vdd.n6850 vdd.n6849 0.019
R62249 vdd.n6879 vdd.n6878 0.019
R62250 vdd.n6795 vdd.n6794 0.019
R62251 vdd.n6823 vdd.n6822 0.019
R62252 vdd.n6735 vdd.n6734 0.019
R62253 vdd.n6763 vdd.n6762 0.019
R62254 vdd.n6684 vdd.n6683 0.019
R62255 vdd.n6624 vdd.n6623 0.019
R62256 vdd.n6568 vdd.n6567 0.019
R62257 vdd.n6594 vdd.n6593 0.019
R62258 vdd.n6511 vdd.n6510 0.019
R62259 vdd.n6540 vdd.n6539 0.019
R62260 vdd.n6456 vdd.n6455 0.019
R62261 vdd.n6426 vdd.n6425 0.019
R62262 vdd.n7920 vdd.n7919 0.019
R62263 vdd.n7950 vdd.n7948 0.019
R62264 vdd.n7864 vdd.n7863 0.019
R62265 vdd.n7893 vdd.n7892 0.019
R62266 vdd.n7808 vdd.n7807 0.019
R62267 vdd.n7837 vdd.n7836 0.019
R62268 vdd.n7777 vdd.n7776 0.019
R62269 vdd.n7779 vdd.n7778 0.019
R62270 vdd.n7693 vdd.n7692 0.019
R62271 vdd.n7722 vdd.n7721 0.019
R62272 vdd.n7578 vdd.n7577 0.019
R62273 vdd.n7607 vdd.n7606 0.019
R62274 vdd.n7634 vdd.n7633 0.019
R62275 vdd.n7665 vdd.n7664 0.019
R62276 vdd.n7521 vdd.n7520 0.019
R62277 vdd.n7549 vdd.n7548 0.019
R62278 vdd.n7551 vdd.n7550 0.019
R62279 vdd.n7489 vdd.n7488 0.019
R62280 vdd.n7409 vdd.n7408 0.019
R62281 vdd.n7439 vdd.n7438 0.019
R62282 vdd.n7352 vdd.n7351 0.019
R62283 vdd.n7382 vdd.n7381 0.019
R62284 vdd.n7298 vdd.n7297 0.019
R62285 vdd.n7325 vdd.n7324 0.019
R62286 vdd.n7238 vdd.n7237 0.019
R62287 vdd.n7240 vdd.n7239 0.019
R62288 vdd.n7270 vdd.n7269 0.019
R62289 vdd.n7134 vdd.n7132 0.019
R62290 vdd.n6988 vdd.n6987 0.019
R62291 vdd.n6990 vdd.n6989 0.019
R62292 vdd.n7045 vdd.n7044 0.019
R62293 vdd.n7071 vdd.n7070 0.019
R62294 vdd.n7099 vdd.n7098 0.019
R62295 vdd.n7101 vdd.n7100 0.019
R62296 vdd.n6932 vdd.n6931 0.019
R62297 vdd.n6960 vdd.n6959 0.019
R62298 vdd.n6876 vdd.n6875 0.019
R62299 vdd.n6903 vdd.n6902 0.019
R62300 vdd.n6820 vdd.n6819 0.019
R62301 vdd.n6847 vdd.n6846 0.019
R62302 vdd.n6792 vdd.n6791 0.019
R62303 vdd.n6731 vdd.n6730 0.019
R62304 vdd.n6733 vdd.n6732 0.019
R62305 vdd.n6620 vdd.n6619 0.019
R62306 vdd.n6622 vdd.n6621 0.019
R62307 vdd.n6680 vdd.n6679 0.019
R62308 vdd.n6682 vdd.n6681 0.019
R62309 vdd.n6508 vdd.n6507 0.019
R62310 vdd.n6538 vdd.n6537 0.019
R62311 vdd.n6566 vdd.n6565 0.019
R62312 vdd.n6591 vdd.n6590 0.019
R62313 vdd.n6454 vdd.n6453 0.019
R62314 vdd.n6422 vdd.n6421 0.019
R62315 vdd.n6424 vdd.n6423 0.019
R62316 vdd.n7890 vdd.n7889 0.019
R62317 vdd.n7916 vdd.n7915 0.019
R62318 vdd.n7834 vdd.n7833 0.019
R62319 vdd.n7860 vdd.n7859 0.019
R62320 vdd.n7775 vdd.n7774 0.019
R62321 vdd.n7804 vdd.n7803 0.019
R62322 vdd.n7719 vdd.n7718 0.019
R62323 vdd.n7745 vdd.n7744 0.019
R62324 vdd.n7662 vdd.n7661 0.019
R62325 vdd.n7689 vdd.n7688 0.019
R62326 vdd.n7605 vdd.n7604 0.019
R62327 vdd.n7632 vdd.n7631 0.019
R62328 vdd.n7547 vdd.n7546 0.019
R62329 vdd.n7574 vdd.n7573 0.019
R62330 vdd.n7487 vdd.n7486 0.019
R62331 vdd.n7518 vdd.n7517 0.019
R62332 vdd.n7436 vdd.n7435 0.019
R62333 vdd.n7462 vdd.n7461 0.019
R62334 vdd.n7379 vdd.n7378 0.019
R62335 vdd.n7405 vdd.n7404 0.019
R62336 vdd.n7322 vdd.n7321 0.019
R62337 vdd.n7348 vdd.n7347 0.019
R62338 vdd.n7267 vdd.n7266 0.019
R62339 vdd.n7294 vdd.n7293 0.019
R62340 vdd.n7198 vdd.n7197 0.019
R62341 vdd.n7236 vdd.n7235 0.019
R62342 vdd.n7095 vdd.n7094 0.019
R62343 vdd.n7097 vdd.n7096 0.019
R62344 vdd.n7129 vdd.n7127 0.019
R62345 vdd.n7039 vdd.n7038 0.019
R62346 vdd.n7041 vdd.n7040 0.019
R62347 vdd.n6985 vdd.n6984 0.019
R62348 vdd.n6927 vdd.n6926 0.019
R62349 vdd.n6929 vdd.n6928 0.019
R62350 vdd.n6958 vdd.n6957 0.019
R62351 vdd.n6871 vdd.n6870 0.019
R62352 vdd.n6873 vdd.n6872 0.019
R62353 vdd.n6817 vdd.n6816 0.019
R62354 vdd.n6756 vdd.n6755 0.019
R62355 vdd.n6758 vdd.n6757 0.019
R62356 vdd.n6790 vdd.n6789 0.019
R62357 vdd.n6703 vdd.n6702 0.019
R62358 vdd.n6648 vdd.n6647 0.019
R62359 vdd.n6677 vdd.n6676 0.019
R62360 vdd.n6587 vdd.n6586 0.019
R62361 vdd.n6589 vdd.n6588 0.019
R62362 vdd.n6617 vdd.n6616 0.019
R62363 vdd.n6532 vdd.n6531 0.019
R62364 vdd.n6534 vdd.n6533 0.019
R62365 vdd.n6477 vdd.n6476 0.019
R62366 vdd.n6417 vdd.n6416 0.019
R62367 vdd.n6419 vdd.n6418 0.019
R62368 vdd.n6451 vdd.n6450 0.019
R62369 vdd.n7913 vdd.n7912 0.019
R62370 vdd.n7856 vdd.n7855 0.019
R62371 vdd.n7858 vdd.n7857 0.019
R62372 vdd.n7800 vdd.n7799 0.019
R62373 vdd.n7802 vdd.n7801 0.019
R62374 vdd.n7742 vdd.n7741 0.019
R62375 vdd.n7772 vdd.n7771 0.019
R62376 vdd.n7685 vdd.n7684 0.019
R62377 vdd.n7687 vdd.n7686 0.019
R62378 vdd.n7628 vdd.n7627 0.019
R62379 vdd.n7630 vdd.n7629 0.019
R62380 vdd.n7570 vdd.n7569 0.019
R62381 vdd.n7572 vdd.n7571 0.019
R62382 vdd.n7514 vdd.n7513 0.019
R62383 vdd.n7516 vdd.n7515 0.019
R62384 vdd.n7459 vdd.n7458 0.019
R62385 vdd.n7484 vdd.n7483 0.019
R62386 vdd.n7402 vdd.n7401 0.019
R62387 vdd.n7433 vdd.n7432 0.019
R62388 vdd.n7344 vdd.n7343 0.019
R62389 vdd.n7346 vdd.n7345 0.019
R62390 vdd.n7290 vdd.n7289 0.019
R62391 vdd.n7292 vdd.n7291 0.019
R62392 vdd.n7232 vdd.n7231 0.019
R62393 vdd.n7234 vdd.n7233 0.019
R62394 vdd.n7123 vdd.n7122 0.019
R62395 vdd.n7126 vdd.n7125 0.019
R62396 vdd.n7066 vdd.n7065 0.019
R62397 vdd.n7093 vdd.n7092 0.019
R62398 vdd.n7012 vdd.n7011 0.019
R62399 vdd.n7014 vdd.n7013 0.019
R62400 vdd.n6955 vdd.n6954 0.019
R62401 vdd.n6982 vdd.n6981 0.019
R62402 vdd.n6898 vdd.n6897 0.019
R62403 vdd.n6900 vdd.n6899 0.019
R62404 vdd.n6843 vdd.n6842 0.019
R62405 vdd.n6869 vdd.n6868 0.019
R62406 vdd.n6787 vdd.n6786 0.019
R62407 vdd.n6814 vdd.n6813 0.019
R62408 vdd.n6726 vdd.n6725 0.019
R62409 vdd.n6754 vdd.n6753 0.019
R62410 vdd.n6673 vdd.n6672 0.019
R62411 vdd.n6675 vdd.n6674 0.019
R62412 vdd.n6613 vdd.n6612 0.019
R62413 vdd.n6615 vdd.n6614 0.019
R62414 vdd.n6561 vdd.n6560 0.019
R62415 vdd.n6585 vdd.n6584 0.019
R62416 vdd.n6504 vdd.n6503 0.019
R62417 vdd.n6530 vdd.n6529 0.019
R62418 vdd.n6447 vdd.n6446 0.019
R62419 vdd.n6449 vdd.n6448 0.019
R62420 vdd.n6383 vdd.n6382 0.019
R62421 vdd.n6415 vdd.n6414 0.019
R62422 vdd.n6380 vdd.n6379 0.019
R62423 vdd.n7943 vdd.n7942 0.019
R62424 vdd.n7945 vdd.n7944 0.019
R62425 vdd.n7941 vdd.n7940 0.019
R62426 vdd.n7886 vdd.n7884 0.019
R62427 vdd.n7911 vdd.n7910 0.019
R62428 vdd.n7939 vdd.n7938 0.019
R62429 vdd.n7830 vdd.n7828 0.019
R62430 vdd.n7854 vdd.n7853 0.019
R62431 vdd.n7770 vdd.n7768 0.019
R62432 vdd.n7798 vdd.n7797 0.019
R62433 vdd.n7715 vdd.n7713 0.019
R62434 vdd.n7740 vdd.n7739 0.019
R62435 vdd.n7658 vdd.n7656 0.019
R62436 vdd.n7683 vdd.n7682 0.019
R62437 vdd.n7601 vdd.n7599 0.019
R62438 vdd.n7626 vdd.n7625 0.019
R62439 vdd.n7543 vdd.n7541 0.019
R62440 vdd.n7568 vdd.n7567 0.019
R62441 vdd.n7482 vdd.n7480 0.019
R62442 vdd.n7512 vdd.n7511 0.019
R62443 vdd.n7431 vdd.n7429 0.019
R62444 vdd.n7457 vdd.n7456 0.019
R62445 vdd.n7375 vdd.n7373 0.019
R62446 vdd.n7400 vdd.n7399 0.019
R62447 vdd.n7318 vdd.n7316 0.019
R62448 vdd.n7342 vdd.n7341 0.019
R62449 vdd.n7263 vdd.n7261 0.019
R62450 vdd.n7288 vdd.n7287 0.019
R62451 vdd.n7192 vdd.n7190 0.019
R62452 vdd.n7230 vdd.n7229 0.019
R62453 vdd.n7091 vdd.n7089 0.019
R62454 vdd.n7121 vdd.n7119 0.019
R62455 vdd.n7036 vdd.n7034 0.019
R62456 vdd.n7064 vdd.n7063 0.019
R62457 vdd.n6980 vdd.n6978 0.019
R62458 vdd.n7010 vdd.n7009 0.019
R62459 vdd.n6920 vdd.n6919 0.019
R62460 vdd.n6924 vdd.n6922 0.019
R62461 vdd.n6953 vdd.n6952 0.019
R62462 vdd.n6894 vdd.n6893 0.019
R62463 vdd.n6838 vdd.n6837 0.019
R62464 vdd.n6841 vdd.n6840 0.019
R62465 vdd.n6781 vdd.n6780 0.019
R62466 vdd.n6784 vdd.n6783 0.019
R62467 vdd.n6722 vdd.n6721 0.019
R62468 vdd.n6724 vdd.n6723 0.019
R62469 vdd.n6644 vdd.n6642 0.019
R62470 vdd.n6671 vdd.n6670 0.019
R62471 vdd.n6608 vdd.n6607 0.019
R62472 vdd.n6610 vdd.n6609 0.019
R62473 vdd.n6528 vdd.n6527 0.019
R62474 vdd.n6558 vdd.n6557 0.019
R62475 vdd.n6498 vdd.n6497 0.019
R62476 vdd.n6501 vdd.n6500 0.019
R62477 vdd.n6441 vdd.n6440 0.019
R62478 vdd.n6444 vdd.n6443 0.019
R62479 vdd.n6375 vdd.n6374 0.019
R62480 vdd.n6377 vdd.n6376 0.019
R62481 vdd.n7956 vdd.n7955 0.019
R62482 vdd.n7976 vdd.n7975 0.019
R62483 vdd.n7088 vdd.n7086 0.019
R62484 vdd.n7228 vdd.n7227 0.019
R62485 vdd.n7259 vdd.n7257 0.019
R62486 vdd.n7286 vdd.n7285 0.019
R62487 vdd.n7340 vdd.n7338 0.019
R62488 vdd.n7372 vdd.n7370 0.019
R62489 vdd.n7398 vdd.n7396 0.019
R62490 vdd.n7428 vdd.n7426 0.019
R62491 vdd.n7455 vdd.n7453 0.019
R62492 vdd.n7479 vdd.n7477 0.019
R62493 vdd.n7510 vdd.n7508 0.019
R62494 vdd.n7540 vdd.n7538 0.019
R62495 vdd.n7566 vdd.n7564 0.019
R62496 vdd.n7598 vdd.n7596 0.019
R62497 vdd.n7624 vdd.n7622 0.019
R62498 vdd.n7655 vdd.n7653 0.019
R62499 vdd.n7681 vdd.n7679 0.019
R62500 vdd.n7712 vdd.n7710 0.019
R62501 vdd.n7738 vdd.n7736 0.019
R62502 vdd.n7767 vdd.n7765 0.019
R62503 vdd.n7796 vdd.n7794 0.019
R62504 vdd.n7827 vdd.n7825 0.019
R62505 vdd.n6864 vdd.n6863 0.019
R62506 vdd.n6641 vdd.n6639 0.019
R62507 vdd.n6411 vdd.n6409 0.019
R62508 vdd.n687 vdd.n686 0.018
R62509 vdd.n1165 vdd.n1164 0.018
R62510 vdd.n5181 vdd.n5178 0.018
R62511 vdd.n29950 vdd.n29949 0.018
R62512 vdd.n30594 vdd.n30282 0.018
R62513 vdd.n34344 vdd.n34343 0.018
R62514 vdd.n27640 vdd.n27638 0.018
R62515 vdd.n4771 vdd.n4713 0.018
R62516 vdd.n11754 vdd.n11683 0.018
R62517 vdd.n21835 vdd.n21834 0.018
R62518 vdd.n34440 vdd.n34439 0.018
R62519 vdd.n25766 vdd.n25765 0.018
R62520 vdd.n776 vdd.n773 0.018
R62521 vdd.n4706 vdd.n4705 0.018
R62522 vdd.n32600 vdd.n32599 0.018
R62523 vdd.n29375 vdd.n29374 0.018
R62524 vdd.n26236 vdd.n26235 0.018
R62525 vdd.n27421 vdd.n27420 0.018
R62526 vdd.n33363 vdd.n33362 0.018
R62527 vdd.n573 vdd.n572 0.018
R62528 vdd.n1169 vdd.n1168 0.018
R62529 vdd.n586 vdd.n503 0.018
R62530 vdd.n27643 vdd.n27641 0.018
R62531 vdd.n27520 vdd.n27519 0.018
R62532 vdd.n27414 vdd.n27413 0.018
R62533 vdd.n27527 vdd.n27526 0.018
R62534 vdd.n27733 vdd.n27732 0.018
R62535 vdd.n31234 vdd.n31233 0.018
R62536 vdd.n26045 vdd.n26043 0.018
R62537 vdd.n25883 vdd.n25882 0.018
R62538 vdd.n27512 vdd.n27510 0.018
R62539 vdd.n33436 vdd.n33435 0.018
R62540 vdd.n33310 vdd.n33309 0.018
R62541 vdd.n33347 vdd.n33342 0.018
R62542 vdd.n33327 vdd.n33326 0.018
R62543 vdd.n33544 vdd.n33543 0.018
R62544 vdd.n33564 vdd.n33560 0.018
R62545 vdd.n33646 vdd.n33644 0.018
R62546 vdd.n33594 vdd.n33588 0.018
R62547 vdd.n33826 vdd.n33824 0.018
R62548 vdd.n33842 vdd.n33841 0.018
R62549 vdd.n34089 vdd.n34088 0.018
R62550 vdd.n34113 vdd.n34112 0.018
R62551 vdd.n34285 vdd.n34284 0.018
R62552 vdd.n34322 vdd.n34317 0.018
R62553 vdd.n34178 vdd.n34176 0.018
R62554 vdd.n34427 vdd.n34424 0.018
R62555 vdd.n33910 vdd.n33905 0.018
R62556 vdd.n34005 vdd.n34004 0.018
R62557 vdd.n35167 vdd.n35166 0.018
R62558 vdd.n35588 vdd.n35583 0.018
R62559 vdd.n35551 vdd.n35550 0.018
R62560 vdd.n35497 vdd.n35494 0.018
R62561 vdd.n35250 vdd.n35249 0.018
R62562 vdd.n35579 vdd.n35578 0.018
R62563 vdd.n35518 vdd.n35517 0.018
R62564 vdd.n35274 vdd.n35273 0.018
R62565 vdd.n35502 vdd.n35501 0.018
R62566 vdd.n35266 vdd.n35265 0.018
R62567 vdd.n35079 vdd.n35074 0.018
R62568 vdd.n35385 vdd.n35382 0.018
R62569 vdd.n35126 vdd.n35116 0.018
R62570 vdd.n35432 vdd.n35431 0.018
R62571 vdd.n35067 vdd.n35066 0.018
R62572 vdd.n35197 vdd.n35196 0.018
R62573 vdd.n35327 vdd.n35326 0.018
R62574 vdd.n35323 vdd.n35321 0.018
R62575 vdd.n34663 vdd.n34662 0.018
R62576 vdd.n34945 vdd.n34942 0.018
R62577 vdd.n34921 vdd.n34920 0.018
R62578 vdd.n34894 vdd.n34889 0.018
R62579 vdd.n34728 vdd.n34726 0.018
R62580 vdd.n34857 vdd.n34854 0.018
R62581 vdd.n34492 vdd.n34487 0.018
R62582 vdd.n34589 vdd.n34588 0.018
R62583 vdd.n639 vdd.n638 0.018
R62584 vdd.n613 vdd.n608 0.018
R62585 vdd.n1083 vdd.n1081 0.018
R62586 vdd.n840 vdd.n837 0.018
R62587 vdd.n518 vdd.n513 0.018
R62588 vdd.n537 vdd.n536 0.018
R62589 vdd.n551 vdd.n550 0.018
R62590 vdd.n32 vdd.n30 0.018
R62591 vdd.n21 vdd.n20 0.018
R62592 vdd.n52 vdd.n49 0.018
R62593 vdd.n441 vdd.n440 0.018
R62594 vdd.n243 vdd.n238 0.018
R62595 vdd.n244 vdd.n243 0.018
R62596 vdd.n254 vdd.n248 0.018
R62597 vdd.n262 vdd.n259 0.018
R62598 vdd.n101 vdd.n100 0.018
R62599 vdd.n150 vdd.n149 0.018
R62600 vdd.n294 vdd.n290 0.018
R62601 vdd.n6300 vdd.n6299 0.018
R62602 vdd.n5937 vdd.n5932 0.018
R62603 vdd.n5964 vdd.n5963 0.018
R62604 vdd.n5791 vdd.n5790 0.018
R62605 vdd.n6003 vdd.n5995 0.018
R62606 vdd.n5833 vdd.n5806 0.018
R62607 vdd.n6025 vdd.n6024 0.018
R62608 vdd.n6008 vdd.n6007 0.018
R62609 vdd.n5838 vdd.n5837 0.018
R62610 vdd.n6184 vdd.n6179 0.018
R62611 vdd.n6078 vdd.n6075 0.018
R62612 vdd.n6186 vdd.n6185 0.018
R62613 vdd.n6250 vdd.n6249 0.018
R62614 vdd.n6115 vdd.n6114 0.018
R62615 vdd.n6291 vdd.n6290 0.018
R62616 vdd.n5885 vdd.n5884 0.018
R62617 vdd.n5881 vdd.n5879 0.018
R62618 vdd.n5410 vdd.n5409 0.018
R62619 vdd.n5692 vdd.n5689 0.018
R62620 vdd.n5668 vdd.n5667 0.018
R62621 vdd.n5641 vdd.n5636 0.018
R62622 vdd.n5475 vdd.n5473 0.018
R62623 vdd.n5604 vdd.n5601 0.018
R62624 vdd.n5239 vdd.n5234 0.018
R62625 vdd.n5336 vdd.n5335 0.018
R62626 vdd.n4648 vdd.n4647 0.018
R62627 vdd.n5109 vdd.n5108 0.018
R62628 vdd.n4815 vdd.n4814 0.018
R62629 vdd.n5098 vdd.n5097 0.018
R62630 vdd.n5074 vdd.n5073 0.018
R62631 vdd.n4719 vdd.n4716 0.018
R62632 vdd.n4989 vdd.n4984 0.018
R62633 vdd.n4735 vdd.n4734 0.018
R62634 vdd.n5059 vdd.n5056 0.018
R62635 vdd.n4628 vdd.n4623 0.018
R62636 vdd.n4687 vdd.n4686 0.018
R62637 vdd.n4923 vdd.n4922 0.018
R62638 vdd.n4919 vdd.n4918 0.018
R62639 vdd.n4240 vdd.n4239 0.018
R62640 vdd.n4519 vdd.n4516 0.018
R62641 vdd.n4495 vdd.n4494 0.018
R62642 vdd.n4468 vdd.n4463 0.018
R62643 vdd.n4579 vdd.n4578 0.018
R62644 vdd.n4562 vdd.n4561 0.018
R62645 vdd.n4264 vdd.n4263 0.018
R62646 vdd.n4302 vdd.n4300 0.018
R62647 vdd.n4317 vdd.n4316 0.018
R62648 vdd.n4431 vdd.n4428 0.018
R62649 vdd.n4069 vdd.n4064 0.018
R62650 vdd.n4116 vdd.n4106 0.018
R62651 vdd.n4409 vdd.n4408 0.018
R62652 vdd.n4167 vdd.n4166 0.018
R62653 vdd.n28969 vdd.n28959 0.018
R62654 vdd.n27485 vdd.n27484 0.018
R62655 vdd.n27544 vdd.n27539 0.018
R62656 vdd.n27295 vdd.n27291 0.018
R62657 vdd.n27389 vdd.n27388 0.018
R62658 vdd.n27454 vdd.n27449 0.018
R62659 vdd.n27320 vdd.n27318 0.018
R62660 vdd.n25706 vdd.n25705 0.018
R62661 vdd.n25981 vdd.n25976 0.018
R62662 vdd.n25747 vdd.n25743 0.018
R62663 vdd.n25835 vdd.n25834 0.018
R62664 vdd.n25900 vdd.n25895 0.018
R62665 vdd.n25772 vdd.n25770 0.018
R62666 vdd.n25505 vdd.n25500 0.018
R62667 vdd.n25640 vdd.n25636 0.018
R62668 vdd.n31011 vdd.n31010 0.018
R62669 vdd.n3878 vdd.n3808 0.018
R62670 vdd.n2519 vdd.n2432 0.018
R62671 vdd.n1861 vdd.n1860 0.018
R62672 vdd.n26350 vdd.n26349 0.018
R62673 vdd.n31827 vdd.n31708 0.018
R62674 vdd.n32043 vdd.n32042 0.018
R62675 vdd.n32295 vdd.n32294 0.018
R62676 vdd.n32296 vdd.n32295 0.018
R62677 vdd.n32383 vdd.n32382 0.018
R62678 vdd.n12583 vdd.n12582 0.018
R62679 vdd.n12577 vdd.n10127 0.018
R62680 vdd.n10195 vdd.n10136 0.018
R62681 vdd.n10196 vdd.n10195 0.018
R62682 vdd.n10685 vdd.n10684 0.018
R62683 vdd.n12331 vdd.n12330 0.018
R62684 vdd.n11033 vdd.n11032 0.018
R62685 vdd.n12126 vdd.n11180 0.018
R62686 vdd.n12025 vdd.n12024 0.018
R62687 vdd.n11515 vdd.n11462 0.018
R62688 vdd.n11539 vdd.n11538 0.018
R62689 vdd.n11613 vdd.n11612 0.018
R62690 ldomc_0.otaldom_0.pdiffm_0.vdd vdd.n13740 0.018
R62691 vdd.n11490 vdd.n11489 0.018
R62692 vdd.n11908 ldomc_0.otaldom_0.pcascodeupm_0.vdd 0.018
R62693 vdd.n13126 vdd.n13124 0.018
R62694 vdd.n13194 vdd.n9218 0.018
R62695 vdd.n13192 vdd.n9219 0.018
R62696 vdd.n13181 vdd.n9207 0.018
R62697 vdd.n13212 vdd.n13210 0.018
R62698 vdd.n13252 vdd.n13251 0.018
R62699 vdd.n13271 vdd.n9162 0.018
R62700 vdd.n13273 vdd.n9147 0.018
R62701 vdd.n14320 vdd.n8339 0.018
R62702 vdd.n14353 vdd.n14351 0.018
R62703 vdd.n14400 vdd.n8300 0.018
R62704 vdd.n14425 vdd.n8279 0.018
R62705 vdd.n14423 vdd.n8280 0.018
R62706 vdd.n14458 vdd.n14457 0.018
R62707 vdd.n8257 vdd.n8250 0.018
R62708 vdd.n14492 vdd.n8219 0.018
R62709 vdd.n14650 vdd.n8152 0.018
R62710 vdd.n14666 vdd.n8137 0.018
R62711 vdd.n14668 vdd.n8132 0.018
R62712 vdd.n14691 vdd.n14679 0.018
R62713 vdd.n14689 vdd.n14680 0.018
R62714 vdd.n14709 vdd.n8110 0.018
R62715 vdd.n14736 vdd.n14720 0.018
R62716 vdd.n14734 vdd.n14721 0.018
R62717 vdd.n14753 vdd.n8097 0.018
R62718 vdd.n14755 vdd.n8091 0.018
R62719 vdd.n14768 vdd.n14766 0.018
R62720 vdd.n14793 vdd.n8068 0.018
R62721 vdd.n14796 vdd.n8062 0.018
R62722 vdd.n14824 vdd.n14807 0.018
R62723 vdd.n14822 vdd.n14808 0.018
R62724 vdd.n14838 vdd.n8047 0.018
R62725 vdd.n14840 vdd.n8042 0.018
R62726 vdd.n14865 vdd.n14851 0.018
R62727 vdd.n14863 vdd.n14852 0.018
R62728 vdd.n14901 vdd.n14882 0.018
R62729 vdd.n14899 vdd.n14883 0.018
R62730 vdd.n14888 vdd.n8013 0.018
R62731 vdd.n14921 vdd.n14920 0.018
R62732 vdd.n14936 vdd.n14935 0.018
R62733 vdd.n15049 vdd.n15048 0.018
R62734 vdd.n15063 vdd.n15056 0.018
R62735 vdd.n16721 vdd.n16720 0.018
R62736 vdd.n16722 vdd.n16721 0.018
R62737 vdd.n17128 vdd.n17127 0.018
R62738 vdd.n17400 vdd.n17399 0.018
R62739 vdd.n17658 vdd.n17657 0.018
R62740 vdd.n17929 vdd.n17928 0.018
R62741 vdd.n18201 vdd.n18200 0.018
R62742 vdd.n18357 vdd.n18356 0.018
R62743 vdd.n18377 vdd.n18376 0.018
R62744 vdd.n21677 vdd.n21676 0.018
R62745 vdd.n21093 bandgapmd_0.otam_1.pdiffm_0.vdd 0.018
R62746 vdd.n16809 vdd.n16808 0.018
R62747 vdd.n20678 vdd.n20676 0.018
R62748 vdd.n20662 vdd.n20660 0.018
R62749 vdd.n20646 vdd.n20644 0.018
R62750 vdd.n20627 vdd.n20615 0.018
R62751 vdd.n20611 vdd.n20599 0.018
R62752 vdd.n20595 vdd.n20583 0.018
R62753 vdd.n20579 vdd.n20567 0.018
R62754 vdd.n20563 vdd.n20551 0.018
R62755 vdd.n20465 vdd.n20464 0.018
R62756 vdd.n20456 vdd.n20454 0.018
R62757 vdd.n20441 vdd.n20439 0.018
R62758 vdd.n20425 vdd.n20423 0.018
R62759 vdd.n20409 vdd.n20407 0.018
R62760 vdd.n20384 vdd.n20369 0.018
R62761 vdd.n20365 vdd.n20353 0.018
R62762 vdd.n20349 vdd.n20337 0.018
R62763 vdd.n20333 vdd.n20321 0.018
R62764 vdd.n20317 vdd.n20305 0.018
R62765 vdd.n20301 vdd.n20289 0.018
R62766 vdd.n20285 vdd.n20273 0.018
R62767 vdd.n20269 vdd.n20267 0.018
R62768 vdd.n20253 vdd.n20251 0.018
R62769 vdd.n20237 vdd.n20235 0.018
R62770 vdd.n20221 vdd.n20219 0.018
R62771 vdd.n20205 vdd.n20203 0.018
R62772 vdd.n20189 vdd.n20187 0.018
R62773 vdd.n20173 vdd.n20171 0.018
R62774 vdd.n20148 vdd.n20133 0.018
R62775 vdd.n20129 vdd.n20117 0.018
R62776 vdd.n20113 vdd.n20101 0.018
R62777 vdd.n20097 vdd.n20085 0.018
R62778 vdd.n20081 vdd.n20069 0.018
R62779 vdd.n19354 vdd.n19342 0.018
R62780 vdd.n19370 vdd.n19358 0.018
R62781 vdd.n19386 vdd.n19374 0.018
R62782 vdd.n19402 vdd.n19390 0.018
R62783 vdd.n19421 vdd.n19406 0.018
R62784 vdd.n19437 vdd.n19435 0.018
R62785 vdd.n19453 vdd.n19451 0.018
R62786 vdd.n19469 vdd.n19467 0.018
R62787 vdd.n21998 vdd 0.018
R62788 vdd.n24952 vdd.n24951 0.018
R62789 vdd.n24722 vdd.n24721 0.018
R62790 vdd.n35607 vdd.n35606 0.018
R62791 vdd.n35019 vdd.n35018 0.018
R62792 vdd.n5766 vdd.n5765 0.018
R62793 vdd.n4596 vdd.n4595 0.018
R62794 vdd.n2484 vdd.n2454 0.018
R62795 vdd.n27518 vdd.n27516 0.018
R62796 vdd.n2602 vdd.n2593 0.018
R62797 vdd.n12600 vdd.n10092 0.018
R62798 vdd.n16743 vdd.n16740 0.018
R62799 vdd.n27428 vdd.n27427 0.018
R62800 vdd.n27308 vdd.n27307 0.018
R62801 vdd.n30141 vdd.n30140 0.018
R62802 vdd.n29355 vdd.n29354 0.018
R62803 vdd.n26565 vdd.n26564 0.018
R62804 vdd.n30196 vdd.n30195 0.018
R62805 vdd.n31436 vdd.n31435 0.018
R62806 vdd.n4437 vdd.n4436 0.018
R62807 vdd.n5610 vdd.n5609 0.018
R62808 vdd.n34863 vdd.n34862 0.018
R62809 vdd.n34433 vdd.n34432 0.018
R62810 vdd.n27633 vdd.n27631 0.018
R62811 vdd.n831 vdd.n830 0.018
R62812 vdd.n25973 vdd.n25972 0.018
R62813 vdd.n5060 vdd.n5059 0.018
R62814 vdd.n24902 vdd.n24896 0.018
R62815 vdd.n682 vdd.n681 0.017
R62816 vdd.n4939 vdd.n4936 0.017
R62817 vdd.n27624 vdd.n27622 0.017
R62818 vdd.n25475 vdd.n25473 0.017
R62819 vdd.n25640 vdd.n25634 0.017
R62820 vdd.n6135 vdd.n6134 0.017
R62821 vdd.n30990 vdd.n30989 0.017
R62822 vdd.n34072 vdd.n34071 0.017
R62823 vdd.n35234 vdd.n35233 0.017
R62824 vdd.n34647 vdd.n34646 0.017
R62825 vdd.n6357 vdd.n6356 0.017
R62826 vdd.n5394 vdd.n5393 0.017
R62827 vdd.n4224 vdd.n4223 0.017
R62828 vdd.n4948 vdd.n4947 0.017
R62829 vdd.n27437 vdd.n27436 0.017
R62830 vdd.n27314 vdd.n27313 0.017
R62831 vdd.n30240 vdd.n30239 0.017
R62832 vdd.n25775 vdd.n25774 0.017
R62833 vdd.n32552 vdd.n32551 0.017
R62834 vdd.n33473 vdd.n33472 0.017
R62835 vdd.n33660 vdd.n33659 0.017
R62836 vdd.n33614 vdd.n33613 0.017
R62837 vdd.n33942 vdd.n33941 0.017
R62838 vdd.n34496 vdd.n34495 0.017
R62839 vdd.n487 vdd.n486 0.017
R62840 vdd.n81 vdd.n80 0.017
R62841 vdd.n302 vdd.n301 0.017
R62842 vdd.n353 vdd.n352 0.017
R62843 vdd.n5243 vdd.n5242 0.017
R62844 vdd.n5090 vdd.n5089 0.017
R62845 vdd.n5136 vdd.n5135 0.017
R62846 vdd.n5029 vdd.n5028 0.017
R62847 vdd.n5021 vdd.n5020 0.017
R62848 vdd.n4546 vdd.n4515 0.017
R62849 vdd.n4259 vdd.n4255 0.017
R62850 vdd.n4073 vdd.n4072 0.017
R62851 vdd.n4057 vdd.n4056 0.017
R62852 vdd.n4158 vdd.n4157 0.017
R62853 vdd.n2675 vdd.n2673 0.017
R62854 vdd.n26424 vdd.n26423 0.017
R62855 vdd.n25374 vdd.n25373 0.017
R62856 vdd.n3943 vdd.n3782 0.017
R62857 vdd.n2656 vdd.n2579 0.017
R62858 vdd.n10214 vdd.n10076 0.017
R62859 vdd.n10225 vdd.n10133 0.017
R62860 vdd.n10592 vdd.n10589 0.017
R62861 vdd.n12477 vdd.n12476 0.017
R62862 vdd.n12377 vdd.n10746 0.017
R62863 vdd.n10785 vdd.n10752 0.017
R62864 vdd.n10944 vdd.n10926 0.017
R62865 vdd.n10949 vdd.n10948 0.017
R62866 vdd.n12184 vdd.n11089 0.017
R62867 vdd.n11124 vdd.n11111 0.017
R62868 vdd.n12079 vdd.n12078 0.017
R62869 vdd.n11294 vdd.n11293 0.017
R62870 vdd.n11489 vdd.n11468 0.017
R62871 vdd.n11512 vdd.n11456 0.017
R62872 vdd.n11952 vdd.n11541 0.017
R62873 vdd.n10182 vdd.n10143 0.017
R62874 vdd.n10182 vdd.n10181 0.017
R62875 vdd.n11698 vdd.n11696 0.017
R62876 vdd.n11707 vdd.n11700 0.017
R62877 vdd.n11858 vdd.n11810 0.017
R62878 vdd.n11851 vdd.n11850 0.017
R62879 vdd.n24164 vdd.n24162 0.017
R62880 vdd.n24012 vdd.n24010 0.017
R62881 vdd.n23932 vdd.n23930 0.017
R62882 vdd.n23780 vdd.n23778 0.017
R62883 vdd.n23700 vdd.n23698 0.017
R62884 vdd.n23092 vdd.n23090 0.017
R62885 vdd.n23244 vdd.n23242 0.017
R62886 vdd.n23324 vdd.n23322 0.017
R62887 vdd.n23476 vdd.n23474 0.017
R62888 vdd.n23556 vdd.n23554 0.017
R62889 vdd.n22513 vdd.n22511 0.017
R62890 vdd.n22665 vdd.n22663 0.017
R62891 vdd.n22745 vdd.n22743 0.017
R62892 vdd.n22897 vdd.n22895 0.017
R62893 vdd.n22977 vdd.n22975 0.017
R62894 vdd.n16689 vdd.n16685 0.017
R62895 vdd.n16678 vdd.n16677 0.017
R62896 vdd.n16980 vdd.n16969 0.017
R62897 vdd.n16997 vdd.n16996 0.017
R62898 vdd.n17252 vdd.n17241 0.017
R62899 vdd.n17269 vdd.n17268 0.017
R62900 vdd.n17524 vdd.n17513 0.017
R62901 vdd.n17541 vdd.n17540 0.017
R62902 vdd.n17782 vdd.n17771 0.017
R62903 vdd.n17799 vdd.n17798 0.017
R62904 vdd.n18053 vdd.n18042 0.017
R62905 vdd.n18070 vdd.n18069 0.017
R62906 vdd.n16809 vdd.n16797 0.017
R62907 vdd.n18419 vdd.n18418 0.017
R62908 vdd.n18423 vdd.n18422 0.017
R62909 vdd.n16707 vdd.n16706 0.017
R62910 vdd.n16708 vdd.n16707 0.017
R62911 vdd.n21796 vdd.n21793 0.017
R62912 vdd.n21783 vdd.n21781 0.017
R62913 vdd.n21949 vdd.n21901 0.017
R62914 vdd.n21942 vdd.n21941 0.017
R62915 vdd.n24910 vdd.n24909 0.017
R62916 vdd.n24861 vdd.n24860 0.017
R62917 vdd.n24872 vdd.n24871 0.017
R62918 vdd.n24853 vdd.n24852 0.017
R62919 vdd.n24859 vdd.n24858 0.017
R62920 vdd.n24875 vdd.n24874 0.017
R62921 vdd.n34224 vdd.n34221 0.017
R62922 vdd.n33800 vdd.n33799 0.017
R62923 vdd.n25858 vdd.n25856 0.017
R62924 vdd.n33959 vdd.n33887 0.017
R62925 vdd.n34511 vdd.n34446 0.017
R62926 vdd.n5258 vdd.n5193 0.017
R62927 vdd.n4088 vdd.n4023 0.017
R62928 vdd.n33860 vdd.n33856 0.017
R62929 vdd.n961 vdd.n956 0.017
R62930 vdd.n26429 vdd.n26425 0.017
R62931 vdd.n27536 vdd.n27535 0.017
R62932 vdd.n30967 vdd.n30966 0.017
R62933 vdd.n31315 vdd.n31314 0.017
R62934 vdd.n31417 vdd.n31416 0.017
R62935 vdd.n22043 vdd.n22042 0.016
R62936 vdd.n31380 vdd.n31375 0.016
R62937 vdd.n30949 vdd.n30948 0.016
R62938 vdd.n25942 vdd.n25940 0.016
R62939 vdd.n25850 vdd.n25848 0.016
R62940 vdd.n33689 vdd.n33686 0.016
R62941 vdd.n24965 vdd.n24959 0.016
R62942 vdd.n11795 vdd.n11793 0.016
R62943 vdd.n21886 vdd.n21884 0.016
R62944 vdd.n13138 vdd.n9253 0.016
R62945 vdd.n21688 vdd.n21628 0.016
R62946 vdd.n30207 vdd.n30203 0.016
R62947 vdd.n27940 vdd.n27936 0.016
R62948 vdd.n27412 vdd.n27410 0.016
R62949 vdd.n27976 vdd.n27975 0.016
R62950 vdd.n30194 vdd.n30183 0.016
R62951 vdd.n29829 vdd.n29828 0.016
R62952 vdd.n27917 vdd.n27905 0.016
R62953 vdd.n27823 vdd.n27822 0.016
R62954 vdd.n28067 vdd.n28055 0.016
R62955 vdd.n28806 vdd.n28805 0.016
R62956 vdd.n27323 vdd.n27322 0.016
R62957 vdd.n2866 vdd.n2859 0.016
R62958 vdd.n2922 vdd.n2920 0.016
R62959 vdd.n3047 vdd.n3040 0.016
R62960 vdd.n3103 vdd.n3101 0.016
R62961 vdd.n3228 vdd.n3221 0.016
R62962 vdd.n3284 vdd.n3282 0.016
R62963 vdd.n3409 vdd.n3402 0.016
R62964 vdd.n3465 vdd.n3463 0.016
R62965 vdd.n3590 vdd.n3583 0.016
R62966 vdd.n33757 vdd.n33756 0.016
R62967 vdd.n34125 vdd.n34124 0.016
R62968 vdd.n34144 vdd.n34140 0.016
R62969 vdd.n34144 vdd.n34143 0.016
R62970 vdd.n33912 vdd.n33911 0.016
R62971 vdd.n33937 vdd.n33936 0.016
R62972 vdd.n34416 vdd.n34415 0.016
R62973 vdd.n34033 vdd.n34032 0.016
R62974 vdd.n34043 vdd.n34042 0.016
R62975 vdd.n34035 vdd.n34034 0.016
R62976 vdd.n35083 vdd.n35082 0.016
R62977 vdd.n34969 vdd.n34941 0.016
R62978 vdd.n34685 vdd.n34678 0.016
R62979 vdd.n34969 vdd.n34968 0.016
R62980 vdd.n34685 vdd.n34684 0.016
R62981 vdd.n34471 vdd.n34470 0.016
R62982 vdd.n34846 vdd.n34845 0.016
R62983 vdd.n34480 vdd.n34479 0.016
R62984 vdd.n34580 vdd.n34579 0.016
R62985 vdd.n34615 vdd.n34614 0.016
R62986 vdd.n34620 vdd.n34619 0.016
R62987 vdd.n786 vdd.n706 0.016
R62988 vdd.n786 vdd.n785 0.016
R62989 vdd.n643 vdd.n642 0.016
R62990 vdd.n652 vdd.n651 0.016
R62991 vdd.n1067 vdd.n1066 0.016
R62992 vdd.n1101 vdd.n1100 0.016
R62993 vdd.n1141 vdd.n1140 0.016
R62994 vdd.n1136 vdd.n1135 0.016
R62995 vdd.n1124 vdd.n1123 0.016
R62996 vdd.n6226 vdd.n6225 0.016
R62997 vdd.n5716 vdd.n5688 0.016
R62998 vdd.n5432 vdd.n5425 0.016
R62999 vdd.n5716 vdd.n5715 0.016
R63000 vdd.n5432 vdd.n5431 0.016
R63001 vdd.n5218 vdd.n5217 0.016
R63002 vdd.n5593 vdd.n5592 0.016
R63003 vdd.n5227 vdd.n5226 0.016
R63004 vdd.n5327 vdd.n5326 0.016
R63005 vdd.n5362 vdd.n5361 0.016
R63006 vdd.n5367 vdd.n5366 0.016
R63007 vdd.n2068 vdd.n2063 0.016
R63008 vdd.n36005 vdd.n35995 0.016
R63009 vdd.n36077 vdd.n36075 0.016
R63010 vdd.n36236 vdd.n36226 0.016
R63011 vdd.n36308 vdd.n36306 0.016
R63012 vdd.n36467 vdd.n36457 0.016
R63013 vdd.n36539 vdd.n36537 0.016
R63014 vdd.n36698 vdd.n36688 0.016
R63015 vdd.n36770 vdd.n36768 0.016
R63016 vdd.n36929 vdd.n36919 0.016
R63017 vdd.n38056 vdd.n38054 0.016
R63018 vdd.n37984 vdd.n37974 0.016
R63019 vdd.n37825 vdd.n37823 0.016
R63020 vdd.n37753 vdd.n37743 0.016
R63021 vdd.n28195 vdd.n28185 0.016
R63022 vdd.n28267 vdd.n28265 0.016
R63023 vdd.n28426 vdd.n28416 0.016
R63024 vdd.n28498 vdd.n28496 0.016
R63025 vdd.n28657 vdd.n28647 0.016
R63026 vdd.n28729 vdd.n28727 0.016
R63027 vdd.n1684 vdd.n1682 0.016
R63028 vdd.n1628 vdd.n1621 0.016
R63029 vdd.n1503 vdd.n1501 0.016
R63030 vdd.n1447 vdd.n1440 0.016
R63031 vdd.n1322 vdd.n1320 0.016
R63032 vdd.n26788 vdd.n26786 0.016
R63033 vdd.n26913 vdd.n26906 0.016
R63034 vdd.n26969 vdd.n26967 0.016
R63035 vdd.n27094 vdd.n27087 0.016
R63036 vdd.n27150 vdd.n27148 0.016
R63037 vdd.n28991 vdd.n28981 0.016
R63038 vdd.n28928 vdd.n28927 0.016
R63039 vdd.n27927 vdd.n27926 0.016
R63040 vdd.n29782 vdd.n29781 0.016
R63041 vdd.n3865 vdd.n3822 0.016
R63042 vdd.n31929 vdd.n31925 0.016
R63043 vdd.n26179 vdd.n26178 0.016
R63044 vdd.n26350 vdd.n26337 0.016
R63045 vdd.n31950 vdd.n31949 0.016
R63046 vdd.n32368 vdd.n32367 0.016
R63047 vdd.n32468 vdd.n32467 0.016
R63048 vdd.n10209 vdd.n10091 0.016
R63049 vdd.n12435 vdd.n10659 0.016
R63050 vdd.n10696 vdd.n10695 0.016
R63051 vdd.n10850 vdd.n10830 0.016
R63052 vdd.n10855 vdd.n10852 0.016
R63053 vdd.n11025 vdd.n11024 0.016
R63054 vdd.n12228 vdd.n12227 0.016
R63055 vdd.n12128 vdd.n11175 0.016
R63056 vdd.n11206 vdd.n11205 0.016
R63057 vdd.n11359 vdd.n11339 0.016
R63058 vdd.n11364 vdd.n11361 0.016
R63059 vdd.n11603 vdd.n11585 0.016
R63060 vdd.n13140 vdd.n9250 0.016
R63061 vdd.n13139 vdd.n9252 0.016
R63062 vdd.n11514 vdd.n11513 0.016
R63063 vdd.n11540 vdd.n11452 0.016
R63064 vdd.n12574 vdd.n10260 0.016
R63065 vdd.n10174 vdd.n10173 0.016
R63066 vdd.n11760 vdd.n11759 0.016
R63067 vdd.n11916 vdd.n11909 0.016
R63068 vdd.n22255 vdd.n22242 0.016
R63069 vdd.n22131 vdd.n22118 0.016
R63070 vdd.n24132 vdd.n24122 0.016
R63071 vdd.n24052 vdd.n24050 0.016
R63072 vdd.n23900 vdd.n23890 0.016
R63073 vdd.n23820 vdd.n23818 0.016
R63074 vdd.n23668 vdd.n23658 0.016
R63075 vdd.n23132 vdd.n23130 0.016
R63076 vdd.n23212 vdd.n23202 0.016
R63077 vdd.n23364 vdd.n23362 0.016
R63078 vdd.n23444 vdd.n23434 0.016
R63079 vdd.n23596 vdd.n23594 0.016
R63080 vdd.n22553 vdd.n22551 0.016
R63081 vdd.n22633 vdd.n22623 0.016
R63082 vdd.n22785 vdd.n22783 0.016
R63083 vdd.n22865 vdd.n22855 0.016
R63084 vdd.n23017 vdd.n23015 0.016
R63085 vdd.n16738 vdd.n16737 0.016
R63086 vdd.n17108 vdd.n17094 0.016
R63087 vdd.n17144 vdd.n17143 0.016
R63088 vdd.n17380 vdd.n17366 0.016
R63089 vdd.n17416 vdd.n17415 0.016
R63090 vdd.n17638 vdd.n17624 0.016
R63091 vdd.n17674 vdd.n17673 0.016
R63092 vdd.n17909 vdd.n17895 0.016
R63093 vdd.n17945 vdd.n17944 0.016
R63094 vdd.n18181 vdd.n18167 0.016
R63095 vdd.n18217 vdd.n18216 0.016
R63096 vdd.n21701 vdd.n21700 0.016
R63097 vdd.n21682 vdd.n21678 0.016
R63098 vdd.n21690 vdd.n21689 0.016
R63099 vdd.n18417 vdd.n18416 0.016
R63100 vdd.n18421 vdd.n18420 0.016
R63101 vdd.n16796 vdd.n16795 0.016
R63102 vdd.n16762 vdd.n16757 0.016
R63103 vdd.n21840 vdd.n21839 0.016
R63104 vdd.n25044 vdd.n25042 0.016
R63105 vdd.n25008 vdd.n25005 0.016
R63106 vdd.n24619 vdd.n24617 0.016
R63107 vdd.n24584 vdd.n24581 0.016
R63108 vdd.n25140 vdd.n25139 0.016
R63109 vdd.n35345 vdd.n35342 0.016
R63110 vdd.n34761 vdd.n34758 0.016
R63111 vdd.n5508 vdd.n5505 0.016
R63112 vdd.n4335 vdd.n4332 0.016
R63113 vdd.n2241 vdd.n2207 0.016
R63114 vdd.n31380 vdd.n31379 0.016
R63115 vdd.n304 vdd.n303 0.016
R63116 vdd.n29453 vdd.n29452 0.016
R63117 vdd.n27505 vdd.n27503 0.016
R63118 vdd.n27404 vdd.n27402 0.016
R63119 vdd.n29966 vdd.n29965 0.016
R63120 vdd.n29892 vdd.n29891 0.016
R63121 vdd.n388 vdd.n387 0.016
R63122 vdd.n25661 vdd.n25659 0.016
R63123 vdd.n1155 vdd.n1152 0.015
R63124 vdd.n29878 vdd.n29877 0.015
R63125 vdd.n28977 vdd.n28976 0.015
R63126 vdd.n25892 vdd.n25891 0.015
R63127 vdd.n33852 vdd.n33794 0.015
R63128 vdd.n28892 vdd.n28106 0.015
R63129 vdd.n26369 vdd.n26368 0.015
R63130 vdd.n34016 vdd.n34015 0.015
R63131 vdd.n35178 vdd.n35172 0.015
R63132 vdd.n34603 vdd.n34602 0.015
R63133 vdd.n6314 vdd.n6308 0.015
R63134 vdd.n5350 vdd.n5349 0.015
R63135 vdd.n4181 vdd.n4180 0.015
R63136 vdd.n1771 vdd.n1288 0.015
R63137 vdd.n27252 vdd.n27251 0.015
R63138 vdd.n25817 vdd.n25815 0.015
R63139 vdd.n2645 vdd.n2582 0.015
R63140 vdd.n3982 vdd.n3761 0.015
R63141 vdd.n33457 vdd.n33454 0.015
R63142 vdd.n33465 vdd.n33462 0.015
R63143 vdd.n33473 vdd.n33466 0.015
R63144 vdd.n33675 vdd.n33674 0.015
R63145 vdd.n33651 vdd.n33650 0.015
R63146 vdd.n33608 vdd.n33607 0.015
R63147 vdd.n34066 vdd.n34063 0.015
R63148 vdd.n35502 vdd.n35493 0.015
R63149 vdd.n35266 vdd.n35262 0.015
R63150 vdd.n35058 vdd.n35057 0.015
R63151 vdd.n35443 vdd.n35442 0.015
R63152 vdd.n35195 vdd.n35194 0.015
R63153 vdd.n35205 vdd.n35204 0.015
R63154 vdd.n487 vdd.n480 0.015
R63155 vdd.n479 vdd.n476 0.015
R63156 vdd.n471 vdd.n468 0.015
R63157 vdd.n81 vdd.n77 0.015
R63158 vdd.n201 vdd.n198 0.015
R63159 vdd.n300 vdd.n299 0.015
R63160 vdd.n113 vdd.n112 0.015
R63161 vdd.n369 vdd.n368 0.015
R63162 vdd.n344 vdd.n343 0.015
R63163 vdd.n6003 vdd.n6002 0.015
R63164 vdd.n5833 vdd.n5832 0.015
R63165 vdd.n6042 vdd.n6041 0.015
R63166 vdd.n6221 vdd.n6220 0.015
R63167 vdd.n6120 vdd.n6119 0.015
R63168 vdd.n6356 vdd.n6355 0.015
R63169 vdd.n6326 vdd.n6325 0.015
R63170 vdd.n6331 vdd.n6330 0.015
R63171 vdd.n5152 vdd.n5151 0.015
R63172 vdd.n5128 vdd.n5127 0.015
R63173 vdd.n4756 vdd.n4755 0.015
R63174 vdd.n5019 vdd.n5018 0.015
R63175 vdd.n4546 vdd.n4545 0.015
R63176 vdd.n4259 vdd.n4258 0.015
R63177 vdd.n4048 vdd.n4047 0.015
R63178 vdd.n4420 vdd.n4419 0.015
R63179 vdd.n4193 vdd.n4192 0.015
R63180 vdd.n4198 vdd.n4197 0.015
R63181 vdd.n29849 vdd.n29848 0.015
R63182 vdd.n29035 vdd.n29034 0.015
R63183 vdd.n29017 vdd.n27756 0.015
R63184 vdd.n28832 vdd.n28826 0.015
R63185 vdd.n28938 vdd.n28935 0.015
R63186 vdd.n28023 vdd.n28022 0.015
R63187 vdd.n30627 vdd.n30626 0.015
R63188 vdd.n30620 vdd.n30619 0.015
R63189 vdd.n30709 vdd.n30708 0.015
R63190 vdd.n30159 vdd.n30158 0.015
R63191 vdd.n30022 vdd.n30021 0.015
R63192 vdd.n29475 vdd.n29474 0.015
R63193 vdd.n26542 vdd.n26541 0.015
R63194 vdd.n31296 vdd.n31293 0.015
R63195 vdd.n2265 vdd.n2148 0.015
R63196 vdd.n2356 vdd.n2106 0.015
R63197 vdd.n12581 vdd.n12580 0.015
R63198 vdd.n10219 vdd.n10070 0.015
R63199 vdd.n10202 vdd.n10079 0.015
R63200 vdd.n12494 vdd.n10567 0.015
R63201 vdd.n12466 vdd.n12465 0.015
R63202 vdd.n12389 vdd.n12388 0.015
R63203 vdd.n10792 vdd.n10791 0.015
R63204 vdd.n10933 vdd.n10932 0.015
R63205 vdd.n10972 vdd.n10971 0.015
R63206 vdd.n12186 vdd.n11083 0.015
R63207 vdd.n12168 vdd.n12167 0.015
R63208 vdd.n11265 vdd.n11246 0.015
R63209 vdd.n11301 vdd.n11300 0.015
R63210 vdd.n11477 vdd.n11476 0.015
R63211 vdd.n11493 vdd.n11492 0.015
R63212 vdd.n11509 vdd.n11460 0.015
R63213 vdd.n11496 vdd.n11495 0.015
R63214 vdd.n11604 vdd.n11584 0.015
R63215 vdd.n10175 vdd.n10144 0.015
R63216 vdd.n11755 vdd.n11684 0.015
R63217 vdd.n11703 vdd.n11702 0.015
R63218 vdd.n11866 vdd.n11812 0.015
R63219 vdd.n11845 vdd.n11842 0.015
R63220 vdd.n11880 vdd.n11879 0.015
R63221 vdd.n13372 vdd.n13371 0.015
R63222 vdd.n13372 vdd.n9050 0.015
R63223 vdd.n13504 vdd.n8954 0.015
R63224 vdd.n13664 vdd.n13663 0.015
R63225 vdd.n13664 vdd.n8829 0.015
R63226 vdd.n8662 vdd.n8627 0.015
R63227 vdd.n8627 vdd.n8608 0.015
R63228 vdd.n14113 vdd.n14112 0.015
R63229 vdd.n8441 vdd.n8405 0.015
R63230 vdd.n8405 vdd.n8386 0.015
R63231 vdd.n24320 vdd.n24319 0.015
R63232 vdd.n24319 vdd.n24311 0.015
R63233 vdd.n22375 vdd.n22374 0.015
R63234 vdd.n22374 vdd.n22366 0.015
R63235 vdd.n15055 vdd.n15054 0.015
R63236 vdd.n16595 vdd.n16591 0.015
R63237 vdd.n16702 vdd.n16695 0.015
R63238 vdd.n16967 vdd.n16953 0.015
R63239 vdd.n17013 vdd.n17012 0.015
R63240 vdd.n17239 vdd.n17225 0.015
R63241 vdd.n17285 vdd.n17284 0.015
R63242 vdd.n17511 vdd.n17497 0.015
R63243 vdd.n17557 vdd.n17556 0.015
R63244 vdd.n17769 vdd.n17755 0.015
R63245 vdd.n17815 vdd.n17814 0.015
R63246 vdd.n18040 vdd.n18026 0.015
R63247 vdd.n18086 vdd.n18085 0.015
R63248 vdd.n18306 vdd.n18293 0.015
R63249 vdd.n18313 vdd.n18312 0.015
R63250 vdd.n18348 vdd.n18335 0.015
R63251 vdd.n16805 vdd.n16804 0.015
R63252 vdd.n21699 vdd.n21698 0.015
R63253 vdd.n16771 vdd.n16770 0.015
R63254 vdd.n19526 vdd.n19520 0.015
R63255 vdd.n19527 vdd.n19526 0.015
R63256 vdd.n19626 vdd.n19625 0.015
R63257 vdd.n19727 vdd.n19721 0.015
R63258 vdd.n19728 vdd.n19727 0.015
R63259 vdd.n20925 vdd.n20924 0.015
R63260 vdd.n20924 vdd.n20918 0.015
R63261 vdd.n20831 vdd.n20830 0.015
R63262 vdd.n20736 vdd.n20735 0.015
R63263 vdd.n20735 vdd.n20729 0.015
R63264 vdd.n21769 vdd.n21766 0.015
R63265 vdd.n21776 vdd.n21774 0.015
R63266 vdd.n21957 vdd.n21903 0.015
R63267 vdd.n21936 vdd.n21933 0.015
R63268 vdd.n21971 vdd.n21970 0.015
R63269 bandgapmd_0.bg_pmosm_0.vdd vdd.n25248 0.015
R63270 vdd.n25786 vdd.n25785 0.015
R63271 vdd.n32689 vdd.n32687 0.015
R63272 vdd.n29053 vdd.n29051 0.015
R63273 vdd.n25984 vdd.n25983 0.015
R63274 vdd.n27446 vdd.n27445 0.015
R63275 vdd.n30790 vdd.n30789 0.014
R63276 vdd.n29751 vdd.n29750 0.014
R63277 vdd.n35354 vdd.n35353 0.014
R63278 vdd.n34770 vdd.n34769 0.014
R63279 vdd.n5517 vdd.n5516 0.014
R63280 vdd.n4344 vdd.n4343 0.014
R63281 vdd.n31319 vdd.n31307 0.014
R63282 vdd.n1928 vdd.n1927 0.014
R63283 vdd.n28981 vdd.n28978 0.014
R63284 vdd.n27365 vdd.n27363 0.014
R63285 vdd.n26125 vdd.n26124 0.014
R63286 vdd.n29323 vdd.n29321 0.014
R63287 vdd.n24549 vdd.n24537 0.014
R63288 vdd.n31071 vdd.n31044 0.014
R63289 vdd.n27334 vdd.n27333 0.014
R63290 vdd.n2219 vdd.n2210 0.014
R63291 vdd.n27252 vdd.n27246 0.014
R63292 vdd.n33400 vdd.n33395 0.014
R63293 vdd.n33410 vdd.n33407 0.014
R63294 vdd.n33417 vdd.n33416 0.014
R63295 vdd.n33428 vdd.n33427 0.014
R63296 vdd.n33375 vdd.n33374 0.014
R63297 vdd.n33491 vdd.n33490 0.014
R63298 vdd.n33558 vdd.n33555 0.014
R63299 vdd.n33320 vdd.n33317 0.014
R63300 vdd.n33342 vdd.n33341 0.014
R63301 vdd.n33351 vdd.n33350 0.014
R63302 vdd.n33725 vdd.n33720 0.014
R63303 vdd.n33727 vdd.n33726 0.014
R63304 vdd.n33736 vdd.n33730 0.014
R63305 vdd.n33737 vdd.n33736 0.014
R63306 vdd.n33744 vdd.n33741 0.014
R63307 vdd.n33729 vdd.n33728 0.014
R63308 vdd.n33601 vdd.n33598 0.014
R63309 vdd.n33633 vdd.n33630 0.014
R63310 vdd.n33757 vdd.n33753 0.014
R63311 vdd.n33586 vdd.n33585 0.014
R63312 vdd.n33772 vdd.n33771 0.014
R63313 vdd.n33828 vdd.n33827 0.014
R63314 vdd.n34098 vdd.n34097 0.014
R63315 vdd.n34257 vdd.n34256 0.014
R63316 vdd.n34270 vdd.n34269 0.014
R63317 vdd.n34284 vdd.n34281 0.014
R63318 vdd.n34182 vdd.n34179 0.014
R63319 vdd.n34201 vdd.n34200 0.014
R63320 vdd.n34383 vdd.n34382 0.014
R63321 vdd.n34388 vdd.n34383 0.014
R63322 vdd.n34396 vdd.n34393 0.014
R63323 vdd.n33917 vdd.n33914 0.014
R63324 vdd.n34352 vdd.n34351 0.014
R63325 vdd.n33982 vdd.n33977 0.014
R63326 vdd.n34003 vdd.n34000 0.014
R63327 vdd.n35165 vdd.n35162 0.014
R63328 vdd.n35550 vdd.n35547 0.014
R63329 vdd.n35536 vdd.n35535 0.014
R63330 vdd.n35523 vdd.n35522 0.014
R63331 vdd.n35259 vdd.n35258 0.014
R63332 vdd.n35565 vdd.n35564 0.014
R63333 vdd.n35063 vdd.n35060 0.014
R63334 vdd.n35412 vdd.n35409 0.014
R63335 vdd.n35402 vdd.n35401 0.014
R63336 vdd.n35407 vdd.n35402 0.014
R63337 vdd.n35370 vdd.n35369 0.014
R63338 vdd.n35458 vdd.n35457 0.014
R63339 vdd.n35144 vdd.n35139 0.014
R63340 vdd.n35285 vdd.n35284 0.014
R63341 vdd.n35325 vdd.n35324 0.014
R63342 vdd.n34675 vdd.n34674 0.014
R63343 vdd.n34938 vdd.n34937 0.014
R63344 vdd.n34925 vdd.n34924 0.014
R63345 vdd.n34920 vdd.n34917 0.014
R63346 vdd.n34741 vdd.n34729 0.014
R63347 vdd.n34701 vdd.n34700 0.014
R63348 vdd.n34806 vdd.n34805 0.014
R63349 vdd.n34811 vdd.n34806 0.014
R63350 vdd.n34816 vdd.n34813 0.014
R63351 vdd.n34476 vdd.n34473 0.014
R63352 vdd.n34780 vdd.n34779 0.014
R63353 vdd.n34557 vdd.n34552 0.014
R63354 vdd.n34585 vdd.n34582 0.014
R63355 vdd.n719 vdd.n714 0.014
R63356 vdd.n734 vdd.n731 0.014
R63357 vdd.n743 vdd.n742 0.014
R63358 vdd.n978 vdd.n977 0.014
R63359 vdd.n1040 vdd.n996 0.014
R63360 vdd.n630 vdd.n627 0.014
R63361 vdd.n608 vdd.n607 0.014
R63362 vdd.n670 vdd.n669 0.014
R63363 vdd.n889 vdd.n884 0.014
R63364 vdd.n891 vdd.n890 0.014
R63365 vdd.n938 vdd.n937 0.014
R63366 vdd.n937 vdd.n931 0.014
R63367 vdd.n921 vdd.n918 0.014
R63368 vdd.n940 vdd.n939 0.014
R63369 vdd.n1112 vdd.n1109 0.014
R63370 vdd.n1090 vdd.n1087 0.014
R63371 vdd.n513 vdd.n512 0.014
R63372 vdd.n530 vdd.n527 0.014
R63373 vdd.n561 vdd.n560 0.014
R63374 vdd.n585 vdd.n584 0.014
R63375 vdd.n75 vdd.n72 0.014
R63376 vdd.n415 vdd.n414 0.014
R63377 vdd.n425 vdd.n422 0.014
R63378 vdd.n450 vdd.n445 0.014
R63379 vdd.n67 vdd.n66 0.014
R63380 vdd.n429 vdd.n428 0.014
R63381 vdd.n400 vdd.n399 0.014
R63382 vdd.n132 vdd.n129 0.014
R63383 vdd.n145 vdd.n143 0.014
R63384 vdd.n165 vdd.n164 0.014
R63385 vdd.n189 vdd.n186 0.014
R63386 vdd.n107 vdd.n106 0.014
R63387 vdd.n276 vdd.n275 0.014
R63388 vdd.n288 vdd.n287 0.014
R63389 vdd.n351 vdd.n349 0.014
R63390 vdd.n6296 vdd.n6293 0.014
R63391 vdd.n5963 vdd.n5960 0.014
R63392 vdd.n5968 vdd.n5967 0.014
R63393 vdd.n5981 vdd.n5980 0.014
R63394 vdd.n5803 vdd.n5802 0.014
R63395 vdd.n5949 vdd.n5948 0.014
R63396 vdd.n6191 vdd.n6188 0.014
R63397 vdd.n6109 vdd.n6106 0.014
R63398 vdd.n6096 vdd.n6095 0.014
R63399 vdd.n6101 vdd.n6096 0.014
R63400 vdd.n6058 vdd.n6057 0.014
R63401 vdd.n6131 vdd.n6073 0.014
R63402 vdd.n6267 vdd.n6262 0.014
R63403 vdd.n5902 vdd.n5901 0.014
R63404 vdd.n5883 vdd.n5882 0.014
R63405 vdd.n5422 vdd.n5421 0.014
R63406 vdd.n5685 vdd.n5684 0.014
R63407 vdd.n5672 vdd.n5671 0.014
R63408 vdd.n5667 vdd.n5664 0.014
R63409 vdd.n5488 vdd.n5476 0.014
R63410 vdd.n5448 vdd.n5447 0.014
R63411 vdd.n5553 vdd.n5552 0.014
R63412 vdd.n5558 vdd.n5553 0.014
R63413 vdd.n5563 vdd.n5560 0.014
R63414 vdd.n5223 vdd.n5220 0.014
R63415 vdd.n5527 vdd.n5526 0.014
R63416 vdd.n5304 vdd.n5299 0.014
R63417 vdd.n5332 vdd.n5329 0.014
R63418 vdd.n4650 vdd.n4649 0.014
R63419 vdd.n4647 vdd.n4644 0.014
R63420 vdd.n5161 vdd.n5156 0.014
R63421 vdd.n5123 vdd.n5120 0.014
R63422 vdd.n5083 vdd.n5082 0.014
R63423 vdd.n4862 vdd.n4859 0.014
R63424 vdd.n4816 vdd.n4815 0.014
R63425 vdd.n4862 vdd.n4861 0.014
R63426 vdd.n4796 vdd.n4795 0.014
R63427 vdd.n4752 vdd.n4747 0.014
R63428 vdd.n4747 vdd.n4746 0.014
R63429 vdd.n4739 vdd.n4736 0.014
R63430 vdd.n4994 vdd.n4991 0.014
R63431 vdd.n4787 vdd.n4786 0.014
R63432 vdd.n4679 vdd.n4678 0.014
R63433 vdd.n4900 vdd.n4899 0.014
R63434 vdd.n4917 vdd.n4915 0.014
R63435 vdd.n4252 vdd.n4251 0.014
R63436 vdd.n4512 vdd.n4511 0.014
R63437 vdd.n4499 vdd.n4498 0.014
R63438 vdd.n4494 vdd.n4491 0.014
R63439 vdd.n4480 vdd.n4479 0.014
R63440 vdd.n4315 vdd.n4303 0.014
R63441 vdd.n4275 vdd.n4274 0.014
R63442 vdd.n4379 vdd.n4378 0.014
R63443 vdd.n4384 vdd.n4379 0.014
R63444 vdd.n4389 vdd.n4386 0.014
R63445 vdd.n4053 vdd.n4050 0.014
R63446 vdd.n4354 vdd.n4353 0.014
R63447 vdd.n4443 vdd.n4442 0.014
R63448 vdd.n4134 vdd.n4129 0.014
R63449 vdd.n4163 vdd.n4160 0.014
R63450 vdd.n30690 vdd.n30686 0.014
R63451 vdd.n29887 vdd.n29882 0.014
R63452 vdd.n27957 vdd.n27894 0.014
R63453 vdd.n27988 vdd.n27863 0.014
R63454 vdd.n28005 vdd.n27853 0.014
R63455 vdd.n29038 vdd.n29037 0.014
R63456 vdd.n28919 vdd.n28918 0.014
R63457 vdd.n28833 vdd.n28832 0.014
R63458 vdd.n28950 vdd.n28947 0.014
R63459 vdd.n29908 vdd.n29905 0.014
R63460 vdd.n30611 vdd.n30610 0.014
R63461 vdd.n27637 vdd.n27636 0.014
R63462 vdd.n27501 vdd.n27500 0.014
R63463 vdd.n27500 vdd.n27499 0.014
R63464 vdd.n27509 vdd.n27508 0.014
R63465 vdd.n27531 vdd.n27528 0.014
R63466 vdd.n27372 vdd.n27367 0.014
R63467 vdd.n27409 vdd.n27408 0.014
R63468 vdd.n27425 vdd.n27422 0.014
R63469 vdd.n27337 vdd.n27336 0.014
R63470 vdd.n26029 vdd.n26028 0.014
R63471 vdd.n26058 vdd.n26057 0.014
R63472 vdd.n25938 vdd.n25937 0.014
R63473 vdd.n25937 vdd.n25936 0.014
R63474 vdd.n25946 vdd.n25945 0.014
R63475 vdd.n25968 vdd.n25965 0.014
R63476 vdd.n25740 vdd.n25735 0.014
R63477 vdd.n25855 vdd.n25854 0.014
R63478 vdd.n25871 vdd.n25868 0.014
R63479 vdd.n25789 vdd.n25788 0.014
R63480 vdd.n25404 vdd.n25403 0.014
R63481 vdd.n25622 vdd.n25621 0.014
R63482 vdd.n30843 vdd.n30842 0.014
R63483 vdd.n26407 vdd.n26370 0.014
R63484 vdd.n26520 vdd.n26508 0.014
R63485 vdd.n29093 vdd.n29083 0.014
R63486 vdd.n29101 vdd.n29056 0.014
R63487 vdd.n29336 vdd.n29327 0.014
R63488 vdd.n29464 vdd.n29454 0.014
R63489 vdd.n32664 vdd.n32659 0.014
R63490 vdd.n32703 vdd.n32694 0.014
R63491 vdd.n29671 vdd.n29661 0.014
R63492 vdd.n29995 vdd.n29986 0.014
R63493 vdd.n32563 vdd.n32553 0.014
R63494 vdd.n30860 vdd.n30850 0.014
R63495 vdd.n30767 vdd.n30751 0.014
R63496 vdd.n31225 vdd.n31223 0.014
R63497 vdd.n31010 vdd.n31009 0.014
R63498 vdd.n31011 vdd.n31008 0.014
R63499 vdd.n30767 vdd.n30752 0.014
R63500 vdd.n31207 vdd.n31206 0.014
R63501 vdd.n26217 vdd.n26108 0.014
R63502 vdd.n26673 vdd.n26654 0.014
R63503 vdd.n26524 vdd.n26489 0.014
R63504 vdd.n26524 vdd.n26491 0.014
R63505 vdd.n29311 vdd.n29301 0.014
R63506 vdd.n29552 vdd.n29542 0.014
R63507 vdd.n30104 vdd.n30094 0.014
R63508 vdd.n38216 vdd.n35620 0.014
R63509 vdd.n3855 vdd.n3847 0.014
R63510 vdd.n2506 vdd.n2439 0.014
R63511 vdd.n1845 vdd.n1844 0.014
R63512 vdd.n1774 vdd.n1773 0.014
R63513 vdd.n31933 vdd.n31929 0.014
R63514 vdd.n26156 vdd.n26155 0.014
R63515 vdd.n26318 vdd.n26317 0.014
R63516 vdd.n31699 vdd.n31698 0.014
R63517 vdd.n32024 vdd.n32023 0.014
R63518 vdd.n32138 vdd.n32137 0.014
R63519 vdd.n32356 vdd.n32355 0.014
R63520 vdd.n26711 vdd.n26641 0.014
R63521 vdd.n26673 vdd.n26643 0.014
R63522 vdd.n26407 vdd.n26379 0.014
R63523 vdd.n26524 vdd.n26503 0.014
R63524 vdd.n26472 vdd.n26443 0.014
R63525 vdd.n29206 vdd.n29205 0.014
R63526 vdd.n29336 vdd.n29335 0.014
R63527 vdd.n29311 vdd.n29310 0.014
R63528 vdd.n29464 vdd.n29463 0.014
R63529 vdd.n7173 vdd.n7172 0.014
R63530 vdd.n29552 vdd.n29551 0.014
R63531 vdd.n29530 vdd.n29529 0.014
R63532 vdd.n32703 vdd.n32702 0.014
R63533 vdd.n29671 vdd.n29670 0.014
R63534 vdd.n30125 vdd.n30124 0.014
R63535 vdd.n30104 vdd.n30103 0.014
R63536 vdd.n32563 vdd.n32562 0.014
R63537 vdd.n30860 vdd.n30859 0.014
R63538 vdd.n30831 vdd.n30830 0.014
R63539 vdd.n30767 vdd.n30766 0.014
R63540 vdd.n10196 vdd.n10087 0.014
R63541 vdd.n10541 vdd.n10539 0.014
R63542 vdd.n12437 vdd.n10653 0.014
R63543 vdd.n12419 vdd.n12418 0.014
R63544 vdd.n10840 vdd.n10839 0.014
R63545 vdd.n10881 vdd.n10880 0.014
R63546 vdd.n12245 vdd.n10997 0.014
R63547 vdd.n12217 vdd.n12216 0.014
R63548 vdd.n12140 vdd.n12139 0.014
R63549 vdd.n11217 vdd.n11216 0.014
R63550 vdd.n11349 vdd.n11348 0.014
R63551 vdd.n11390 vdd.n11389 0.014
R63552 vdd.n11488 vdd.n11487 0.014
R63553 vdd.n11494 vdd.n11464 0.014
R63554 vdd.n11950 vdd.n11544 0.014
R63555 vdd.n13949 vdd.n13948 0.014
R63556 vdd.n13999 vdd.n8598 0.014
R63557 vdd.n14239 vdd.n14238 0.014
R63558 vdd.n14290 vdd.n8376 0.014
R63559 vdd.n14607 vdd.n14606 0.014
R63560 vdd.n14609 vdd.n14608 0.014
R63561 vdd.n13384 vdd.n13383 0.014
R63562 vdd.n13385 vdd.n9026 0.014
R63563 vdd.n13676 vdd.n13675 0.014
R63564 vdd.n13677 vdd.n8806 0.014
R63565 vdd.n11491 vdd.n11465 0.014
R63566 vdd.n11511 vdd.n11510 0.014
R63567 vdd.n11594 vdd.n11593 0.014
R63568 vdd.n10349 vdd.n10348 0.014
R63569 vdd.n10374 vdd.n10350 0.014
R63570 vdd.n9447 vdd.n9446 0.014
R63571 vdd.n9450 vdd.n9448 0.014
R63572 vdd.n12894 vdd.n9603 0.014
R63573 vdd.n9639 vdd.n9634 0.014
R63574 vdd.n9806 vdd.n9805 0.014
R63575 vdd.n9809 vdd.n9807 0.014
R63576 vdd.n12686 vdd.n9963 0.014
R63577 vdd.n9999 vdd.n9994 0.014
R63578 vdd.n11750 vdd.n11749 0.014
R63579 vdd.n11769 vdd.n11669 0.014
R63580 vdd.n22363 vdd.n22349 0.014
R63581 vdd.n24308 vdd.n22065 0.014
R63582 vdd.n22328 vdd.n22327 0.014
R63583 vdd.n22327 vdd.n22326 0.014
R63584 vdd.n24321 vdd.n24320 0.014
R63585 vdd.n24311 vdd.n24310 0.014
R63586 vdd.n24300 vdd.n24299 0.014
R63587 vdd.n24299 vdd.n24298 0.014
R63588 vdd.n24150 vdd.n24148 0.014
R63589 vdd.n24026 vdd.n24024 0.014
R63590 vdd.n23918 vdd.n23916 0.014
R63591 vdd.n23794 vdd.n23792 0.014
R63592 vdd.n23686 vdd.n23684 0.014
R63593 vdd.n23106 vdd.n23104 0.014
R63594 vdd.n23230 vdd.n23228 0.014
R63595 vdd.n23338 vdd.n23336 0.014
R63596 vdd.n23462 vdd.n23460 0.014
R63597 vdd.n23570 vdd.n23568 0.014
R63598 vdd.n22527 vdd.n22525 0.014
R63599 vdd.n22651 vdd.n22649 0.014
R63600 vdd.n22759 vdd.n22757 0.014
R63601 vdd.n22883 vdd.n22881 0.014
R63602 vdd.n22991 vdd.n22989 0.014
R63603 vdd.n22376 vdd.n22375 0.014
R63604 vdd.n22366 vdd.n22365 0.014
R63605 vdd.n22006 vdd.n22005 0.014
R63606 vdd.n22007 vdd.n22006 0.014
R63607 vdd.n22008 vdd.n22007 0.014
R63608 vdd.n22009 vdd.n22008 0.014
R63609 vdd.n22010 vdd.n22009 0.014
R63610 vdd.n22011 vdd.n22010 0.014
R63611 vdd.n22012 vdd.n22011 0.014
R63612 vdd.n22013 vdd.n22012 0.014
R63613 vdd.n22014 vdd.n22013 0.014
R63614 vdd.n22015 vdd.n22014 0.014
R63615 vdd.n22016 vdd.n22015 0.014
R63616 vdd.n22017 vdd.n22016 0.014
R63617 vdd.n22018 vdd.n22017 0.014
R63618 vdd.n22019 vdd.n22018 0.014
R63619 vdd.n22020 vdd.n22019 0.014
R63620 vdd.n22021 vdd.n22020 0.014
R63621 vdd.n22022 vdd.n22021 0.014
R63622 vdd.n22023 vdd.n22022 0.014
R63623 vdd.n22024 vdd.n22023 0.014
R63624 vdd.n22025 vdd.n22024 0.014
R63625 vdd.n22026 vdd.n22025 0.014
R63626 vdd.n22027 vdd.n22026 0.014
R63627 vdd.n22028 vdd.n22027 0.014
R63628 vdd.n22029 vdd.n22028 0.014
R63629 vdd.n22031 vdd.n22030 0.014
R63630 vdd.n22032 vdd.n22031 0.014
R63631 vdd.n22034 vdd.n22033 0.014
R63632 vdd.n22035 vdd.n22034 0.014
R63633 vdd.n22036 vdd.n22035 0.014
R63634 vdd.n22037 vdd.n22036 0.014
R63635 vdd.n22038 vdd.n22037 0.014
R63636 vdd.n22039 vdd.n22038 0.014
R63637 vdd.n22040 vdd.n22039 0.014
R63638 vdd.n22041 vdd.n22040 0.014
R63639 vdd.n22042 vdd.n22041 0.014
R63640 vdd.n24370 vdd.n24369 0.014
R63641 vdd.n24371 vdd.n24370 0.014
R63642 vdd.n24372 vdd.n24371 0.014
R63643 vdd.n24373 vdd.n24372 0.014
R63644 vdd.n24374 vdd.n24373 0.014
R63645 vdd.n24375 vdd.n24374 0.014
R63646 vdd.n24376 vdd.n24375 0.014
R63647 vdd.n24377 vdd.n24376 0.014
R63648 vdd.n24378 vdd.n24377 0.014
R63649 vdd.n24379 vdd.n24378 0.014
R63650 vdd.n24380 vdd.n24379 0.014
R63651 vdd.n24381 vdd.n24380 0.014
R63652 vdd.n24382 vdd.n24381 0.014
R63653 vdd.n24383 vdd.n24382 0.014
R63654 vdd.n24384 vdd.n24383 0.014
R63655 vdd.n24385 vdd.n24384 0.014
R63656 vdd.n24386 vdd.n24385 0.014
R63657 vdd.n24388 vdd.n24387 0.014
R63658 vdd.n24389 vdd.n24388 0.014
R63659 vdd.n24391 vdd.n24390 0.014
R63660 vdd.n24392 vdd.n24391 0.014
R63661 vdd.n24393 vdd.n24392 0.014
R63662 vdd.n24394 vdd.n24393 0.014
R63663 vdd.n24395 vdd.n24394 0.014
R63664 vdd.n24396 vdd.n24395 0.014
R63665 vdd.n24397 vdd.n24396 0.014
R63666 vdd.n24398 vdd.n24397 0.014
R63667 vdd.n24399 vdd.n24398 0.014
R63668 vdd.n24400 vdd.n24399 0.014
R63669 vdd.n24401 vdd.n24400 0.014
R63670 vdd.n24402 vdd.n24401 0.014
R63671 vdd.n24403 vdd.n24402 0.014
R63672 vdd.n24404 vdd.n24403 0.014
R63673 vdd.n24405 vdd.n24404 0.014
R63674 vdd.n24406 vdd.n24405 0.014
R63675 vdd.n24407 vdd.n24406 0.014
R63676 vdd.n16730 vdd.n16722 0.014
R63677 vdd.n16888 vdd.n16887 0.014
R63678 vdd.n17092 vdd.n17078 0.014
R63679 vdd.n17160 vdd.n17159 0.014
R63680 vdd.n17364 vdd.n17350 0.014
R63681 vdd.n17432 vdd.n17431 0.014
R63682 vdd.n17622 vdd.n17608 0.014
R63683 vdd.n17690 vdd.n17689 0.014
R63684 vdd.n17893 vdd.n17879 0.014
R63685 vdd.n17961 vdd.n17960 0.014
R63686 vdd.n18165 vdd.n18151 0.014
R63687 vdd.n18232 vdd.n18231 0.014
R63688 vdd.n18310 vdd.n18309 0.014
R63689 vdd.n18315 vdd.n18314 0.014
R63690 vdd.n18389 vdd.n18388 0.014
R63691 vdd.n19035 vdd.n19020 0.014
R63692 vdd.n19019 vdd.n19018 0.014
R63693 vdd.n18776 vdd.n18761 0.014
R63694 vdd.n18760 vdd.n18759 0.014
R63695 vdd.n18517 vdd.n18502 0.014
R63696 vdd.n18501 vdd.n18500 0.014
R63697 vdd.n21401 vdd.n21386 0.014
R63698 vdd.n21385 vdd.n21384 0.014
R63699 vdd.n21142 vdd.n21127 0.014
R63700 vdd.n21126 vdd.n21125 0.014
R63701 vdd.n16807 vdd.n16806 0.014
R63702 vdd.n16799 vdd.n16798 0.014
R63703 vdd.n18431 vdd.n18430 0.014
R63704 vdd.n15417 vdd.n15416 0.014
R63705 vdd.n15419 vdd.n15418 0.014
R63706 vdd.n15667 vdd.n15666 0.014
R63707 vdd.n15669 vdd.n15668 0.014
R63708 vdd.n15923 vdd.n15922 0.014
R63709 vdd.n15925 vdd.n15924 0.014
R63710 vdd.n16179 vdd.n16178 0.014
R63711 vdd.n16181 vdd.n16180 0.014
R63712 vdd.n16435 vdd.n16434 0.014
R63713 vdd.n16437 vdd.n16436 0.014
R63714 vdd.n21823 vdd.n21822 0.014
R63715 vdd.n21857 vdd.n21856 0.014
R63716 vdd.n325 vdd.n324 0.014
R63717 vdd.n27547 vdd.n27546 0.014
R63718 vdd.n33701 vdd.n33700 0.014
R63719 vdd.n29847 vdd.n29846 0.014
R63720 vdd.n27785 vdd.n27784 0.014
R63721 vdd.n26034 vdd.n26032 0.014
R63722 vdd.n25931 vdd.n25929 0.014
R63723 vdd.n25839 vdd.n25837 0.014
R63724 vdd.n28120 vdd.n28119 0.014
R63725 vdd.n25422 vdd.n25417 0.014
R63726 vdd.n26568 vdd.n26567 0.014
R63727 vdd.n29359 vdd.n29357 0.014
R63728 vdd.n30145 vdd.n30143 0.014
R63729 vdd.n35424 vdd.n35423 0.014
R63730 vdd.n6214 vdd.n6213 0.014
R63731 vdd.n30250 vdd.n30249 0.013
R63732 vdd.n5010 vdd.n5008 0.013
R63733 vdd.n4401 vdd.n4400 0.013
R63734 vdd.n24941 vdd.n24940 0.013
R63735 vdd.n34828 vdd.n34827 0.013
R63736 vdd.n5575 vdd.n5574 0.013
R63737 vdd.n24899 vdd.n24898 0.013
R63738 vdd.n32691 vdd.n32690 0.013
R63739 vdd.n6370 vdd.n6369 0.013
R63740 vdd.n208 vdd.n207 0.013
R63741 vdd.n2631 vdd.n2588 0.013
R63742 vdd.n3924 vdd.n3796 0.013
R63743 vdd.n3967 vdd.n3767 0.013
R63744 vdd.n31216 vdd.n31197 0.013
R63745 vdd.n25536 vdd.n25535 0.013
R63746 vdd.n2776 vdd.n2774 0.013
R63747 vdd.n2826 vdd.n2824 0.013
R63748 vdd.n2957 vdd.n2955 0.013
R63749 vdd.n3007 vdd.n3005 0.013
R63750 vdd.n3138 vdd.n3136 0.013
R63751 vdd.n3188 vdd.n3186 0.013
R63752 vdd.n3319 vdd.n3317 0.013
R63753 vdd.n3369 vdd.n3367 0.013
R63754 vdd.n3500 vdd.n3498 0.013
R63755 vdd.n3550 vdd.n3548 0.013
R63756 vdd.n1763 vdd.n1761 0.013
R63757 vdd.n34290 vdd.n34289 0.013
R63758 vdd.n34263 vdd.n34262 0.013
R63759 vdd.n34299 vdd.n34298 0.013
R63760 vdd.n34211 vdd.n34210 0.013
R63761 vdd.n34436 vdd.n34367 0.013
R63762 vdd.n34436 vdd.n34435 0.013
R63763 vdd.n34906 vdd.n34905 0.013
R63764 vdd.n34997 vdd.n34996 0.013
R63765 vdd.n34988 vdd.n34987 0.013
R63766 vdd.n34748 vdd.n34747 0.013
R63767 vdd.n34869 vdd.n34865 0.013
R63768 vdd.n34869 vdd.n34868 0.013
R63769 vdd.n738 vdd.n737 0.013
R63770 vdd.n751 vdd.n750 0.013
R63771 vdd.n759 vdd.n758 0.013
R63772 vdd.n689 vdd.n590 0.013
R63773 vdd.n689 vdd.n688 0.013
R63774 vdd.n1023 vdd.n1022 0.013
R63775 vdd.n947 vdd.n928 0.013
R63776 vdd.n876 vdd.n875 0.013
R63777 vdd.n947 vdd.n946 0.013
R63778 vdd.n878 vdd.n877 0.013
R63779 vdd.n585 vdd.n578 0.013
R63780 vdd.n454 vdd.n453 0.013
R63781 vdd.n420 vdd.n419 0.013
R63782 vdd.n392 vdd.n391 0.013
R63783 vdd.n174 vdd.n173 0.013
R63784 vdd.n288 vdd.n284 0.013
R63785 vdd.n5830 vdd.n5819 0.013
R63786 vdd.n5653 vdd.n5652 0.013
R63787 vdd.n5744 vdd.n5743 0.013
R63788 vdd.n5735 vdd.n5734 0.013
R63789 vdd.n5495 vdd.n5494 0.013
R63790 vdd.n5616 vdd.n5612 0.013
R63791 vdd.n5616 vdd.n5615 0.013
R63792 vdd.n4862 vdd.n4858 0.013
R63793 vdd.n4787 vdd.n4773 0.013
R63794 vdd.n4663 vdd.n4662 0.013
R63795 vdd.n4677 vdd.n4676 0.013
R63796 vdd.n4910 vdd.n4909 0.013
R63797 vdd.n2673 vdd.n2669 0.013
R63798 vdd.n2000 vdd.n1999 0.013
R63799 vdd.n2005 vdd.n2004 0.013
R63800 vdd.n35890 vdd.n35888 0.013
R63801 vdd.n35953 vdd.n35951 0.013
R63802 vdd.n36121 vdd.n36119 0.013
R63803 vdd.n36184 vdd.n36182 0.013
R63804 vdd.n36352 vdd.n36350 0.013
R63805 vdd.n36415 vdd.n36413 0.013
R63806 vdd.n36583 vdd.n36581 0.013
R63807 vdd.n36646 vdd.n36644 0.013
R63808 vdd.n36814 vdd.n36812 0.013
R63809 vdd.n36877 vdd.n36875 0.013
R63810 vdd.n38100 vdd.n38098 0.013
R63811 vdd.n37932 vdd.n37930 0.013
R63812 vdd.n37869 vdd.n37867 0.013
R63813 vdd.n37701 vdd.n37699 0.013
R63814 vdd.n37638 vdd.n37636 0.013
R63815 vdd.n28311 vdd.n28309 0.013
R63816 vdd.n28374 vdd.n28372 0.013
R63817 vdd.n28542 vdd.n28540 0.013
R63818 vdd.n28605 vdd.n28603 0.013
R63819 vdd.n28773 vdd.n28771 0.013
R63820 vdd.n1719 vdd.n1717 0.013
R63821 vdd.n1588 vdd.n1586 0.013
R63822 vdd.n1538 vdd.n1536 0.013
R63823 vdd.n1407 vdd.n1405 0.013
R63824 vdd.n1357 vdd.n1355 0.013
R63825 vdd.n26823 vdd.n26821 0.013
R63826 vdd.n26873 vdd.n26871 0.013
R63827 vdd.n27004 vdd.n27002 0.013
R63828 vdd.n27054 vdd.n27052 0.013
R63829 vdd.n27185 vdd.n27183 0.013
R63830 vdd.n29767 vdd.n29755 0.013
R63831 vdd.n29842 vdd.n29841 0.013
R63832 vdd.n28027 vdd.n27785 0.013
R63833 vdd.n28865 vdd.n28130 0.013
R63834 vdd.n28843 vdd.n28838 0.013
R63835 vdd.n28995 vdd.n28992 0.013
R63836 vdd.n29008 vdd.n29005 0.013
R63837 vdd.n28027 vdd.n28026 0.013
R63838 vdd.n29921 vdd.n29918 0.013
R63839 vdd.n29942 vdd.n29941 0.013
R63840 vdd.n30602 vdd.n30601 0.013
R63841 vdd.n30757 vdd.n30756 0.013
R63842 vdd.n29070 vdd.n29069 0.013
R63843 vdd.n32670 vdd.n32669 0.013
R63844 vdd.n31374 vdd.n31373 0.013
R63845 vdd.n26083 vdd.n26082 0.013
R63846 vdd.n26092 vdd.n25360 0.013
R63847 vdd.n25354 vdd.n25339 0.013
R63848 vdd.n26226 vdd.n26094 0.013
R63849 vdd.n26718 vdd.n26584 0.013
R63850 vdd.n26578 vdd.n26561 0.013
R63851 vdd.n26250 vdd.n26231 0.013
R63852 vdd.n26267 vdd.n26252 0.013
R63853 vdd.n26415 vdd.n26270 0.013
R63854 vdd.n26557 vdd.n26540 0.013
R63855 vdd.n26438 vdd.n26419 0.013
R63856 vdd.n26534 vdd.n26442 0.013
R63857 vdd.n27681 vdd.n27664 0.013
R63858 vdd.n27704 vdd.n27685 0.013
R63859 vdd.n27723 vdd.n27708 0.013
R63860 vdd.n27743 vdd.n27727 0.013
R63861 vdd.n29110 vdd.n29042 0.013
R63862 vdd.n29144 vdd.n29116 0.013
R63863 vdd.n29172 vdd.n29147 0.013
R63864 vdd.n29248 vdd.n29219 0.013
R63865 vdd.n29214 vdd.n29179 0.013
R63866 vdd.n29266 vdd.n29253 0.013
R63867 vdd.n29346 vdd.n29270 0.013
R63868 vdd.n29367 vdd.n29351 0.013
R63869 vdd.n29389 vdd.n29371 0.013
R63870 vdd.n29405 vdd.n29392 0.013
R63871 vdd.n29464 vdd.n29439 0.013
R63872 vdd.n29472 vdd.n29410 0.013
R63873 vdd.n29481 vdd.n29480 0.013
R63874 vdd.n7218 vdd.n7213 0.013
R63875 vdd.n29561 vdd.n29497 0.013
R63876 vdd.n29588 vdd.n29569 0.013
R63877 vdd.n29610 vdd.n29592 0.013
R63878 vdd.n29628 vdd.n29614 0.013
R63879 vdd.n32731 vdd.n32714 0.013
R63880 vdd.n32711 vdd.n32638 0.013
R63881 vdd.n32634 vdd.n32620 0.013
R63882 vdd.n29679 vdd.n29630 0.013
R63883 vdd.n30035 vdd.n30017 0.013
R63884 vdd.n30004 vdd.n29956 0.013
R63885 vdd.n30068 vdd.n30039 0.013
R63886 vdd.n30133 vdd.n30072 0.013
R63887 vdd.n30155 vdd.n30137 0.013
R63888 vdd.n32613 vdd.n32596 0.013
R63889 vdd.n32593 vdd.n32575 0.013
R63890 vdd.n32571 vdd.n31407 0.013
R63891 vdd.n30173 vdd.n30157 0.013
R63892 vdd.n30869 vdd.n30724 0.013
R63893 vdd.n30720 vdd.n30702 0.013
R63894 vdd.n30892 vdd.n30873 0.013
R63895 vdd.n30915 vdd.n30895 0.013
R63896 vdd.n30927 vdd.n30926 0.013
R63897 vdd.n30936 vdd.n30919 0.013
R63898 vdd.n31400 vdd.n31367 0.013
R63899 vdd.n31364 vdd.n31351 0.013
R63900 vdd.n31347 vdd.n31331 0.013
R63901 vdd.n30984 vdd.n30938 0.013
R63902 vdd.n27660 vdd.n25357 0.013
R63903 vdd.n26092 vdd.n26091 0.013
R63904 vdd.n27660 vdd.n25337 0.013
R63905 vdd.n25354 vdd.n25353 0.013
R63906 vdd.n27660 vdd.n26227 0.013
R63907 vdd.n26226 vdd.n26225 0.013
R63908 vdd.n27660 vdd.n26719 0.013
R63909 vdd.n27660 vdd.n26580 0.013
R63910 vdd.n26578 vdd.n26577 0.013
R63911 vdd.n27660 vdd.n26229 0.013
R63912 vdd.n26250 vdd.n26249 0.013
R63913 vdd.n27660 vdd.n26268 0.013
R63914 vdd.n26267 vdd.n26266 0.013
R63915 vdd.n27660 vdd.n26416 0.013
R63916 vdd.n26415 vdd.n26414 0.013
R63917 vdd.n27660 vdd.n26538 0.013
R63918 vdd.n27660 vdd.n26440 0.013
R63919 vdd.n26438 vdd.n26437 0.013
R63920 vdd.n27660 vdd.n26535 0.013
R63921 vdd.n26534 vdd.n26533 0.013
R63922 vdd.n32737 vdd.n27662 0.013
R63923 vdd.n27681 vdd.n27680 0.013
R63924 vdd.n32737 vdd.n27705 0.013
R63925 vdd.n27704 vdd.n27703 0.013
R63926 vdd.n32737 vdd.n27706 0.013
R63927 vdd.n32737 vdd.n27745 0.013
R63928 vdd.n32737 vdd.n29112 0.013
R63929 vdd.n32737 vdd.n29114 0.013
R63930 vdd.n32737 vdd.n29174 0.013
R63931 vdd.n32737 vdd.n29217 0.013
R63932 vdd.n32737 vdd.n29177 0.013
R63933 vdd.n32737 vdd.n29251 0.013
R63934 vdd.n32737 vdd.n29348 0.013
R63935 vdd.n29346 vdd.n29345 0.013
R63936 vdd.n32737 vdd.n29349 0.013
R63937 vdd.n29367 vdd.n29366 0.013
R63938 vdd.n32737 vdd.n29390 0.013
R63939 vdd.n32737 vdd.n29407 0.013
R63940 vdd.n32737 vdd.n29409 0.013
R63941 vdd.n32737 vdd.n29493 0.013
R63942 vdd.n7218 vdd.n7217 0.013
R63943 vdd.n32737 vdd.n29495 0.013
R63944 vdd.n29561 vdd.n29560 0.013
R63945 vdd.n32737 vdd.n29567 0.013
R63946 vdd.n29588 vdd.n29587 0.013
R63947 vdd.n32737 vdd.n29590 0.013
R63948 vdd.n29610 vdd.n29609 0.013
R63949 vdd.n32737 vdd.n29612 0.013
R63950 vdd.n32737 vdd.n32733 0.013
R63951 vdd.n32731 vdd.n32730 0.013
R63952 vdd.n32737 vdd.n32636 0.013
R63953 vdd.n32711 vdd.n32710 0.013
R63954 vdd.n32737 vdd.n32618 0.013
R63955 vdd.n32634 vdd.n32633 0.013
R63956 vdd.n32737 vdd.n29680 0.013
R63957 vdd.n29679 vdd.n29678 0.013
R63958 vdd.n32737 vdd.n30015 0.013
R63959 vdd.n30035 vdd.n30034 0.013
R63960 vdd.n32737 vdd.n29954 0.013
R63961 vdd.n30004 vdd.n30003 0.013
R63962 vdd.n32737 vdd.n30037 0.013
R63963 vdd.n30068 vdd.n30067 0.013
R63964 vdd.n32737 vdd.n30070 0.013
R63965 vdd.n30133 vdd.n30132 0.013
R63966 vdd.n32737 vdd.n30135 0.013
R63967 vdd.n30155 vdd.n30154 0.013
R63968 vdd.n32737 vdd.n32614 0.013
R63969 vdd.n32613 vdd.n32612 0.013
R63970 vdd.n32737 vdd.n32573 0.013
R63971 vdd.n32593 vdd.n32592 0.013
R63972 vdd.n32737 vdd.n31405 0.013
R63973 vdd.n32571 vdd.n32570 0.013
R63974 vdd.n32737 vdd.n30174 0.013
R63975 vdd.n30173 vdd.n30172 0.013
R63976 vdd.n32737 vdd.n30722 0.013
R63977 vdd.n30869 vdd.n30868 0.013
R63978 vdd.n32737 vdd.n30700 0.013
R63979 vdd.n30720 vdd.n30719 0.013
R63980 vdd.n32737 vdd.n30871 0.013
R63981 vdd.n30892 vdd.n30891 0.013
R63982 vdd.n32737 vdd.n30894 0.013
R63983 vdd.n30915 vdd.n30914 0.013
R63984 vdd.n32737 vdd.n30917 0.013
R63985 vdd.n30936 vdd.n30935 0.013
R63986 vdd.n32737 vdd.n31401 0.013
R63987 vdd.n31400 vdd.n31399 0.013
R63988 vdd.n32737 vdd.n31349 0.013
R63989 vdd.n31364 vdd.n31363 0.013
R63990 vdd.n32737 vdd.n31329 0.013
R63991 vdd.n31347 vdd.n31346 0.013
R63992 vdd.n32737 vdd.n30985 0.013
R63993 vdd.n30984 vdd.n30983 0.013
R63994 vdd.n32737 vdd.n31306 0.013
R63995 vdd.n3930 vdd.n3790 0.013
R63996 vdd.n2268 vdd.n2146 0.013
R63997 vdd.n1927 vdd.n1926 0.013
R63998 vdd.n31881 vdd.n31693 0.013
R63999 vdd.n31304 vdd.n31303 0.013
R64000 vdd.n12496 vdd.n10561 0.013
R64001 vdd.n10634 vdd.n10608 0.013
R64002 vdd.n10744 vdd.n10725 0.013
R64003 vdd.n10803 vdd.n10779 0.013
R64004 vdd.n12298 vdd.n10899 0.013
R64005 vdd.n10979 vdd.n10978 0.013
R64006 vdd.n12198 vdd.n12197 0.013
R64007 vdd.n12157 vdd.n12156 0.013
R64008 vdd.n11254 vdd.n11253 0.013
R64009 vdd.n11312 vdd.n11287 0.013
R64010 vdd.n11992 vdd.n11408 0.013
R64011 vdd.n13875 vdd.n8704 0.013
R64012 vdd.n14102 vdd.n14101 0.013
R64013 vdd.n14164 vdd.n8481 0.013
R64014 vdd.n14390 vdd.n8292 0.013
R64015 vdd.n14444 vdd.n8266 0.013
R64016 vdd.n13815 vdd.n13814 0.013
R64017 vdd.n11623 vdd.n11580 0.013
R64018 vdd.n11618 vdd.n11583 0.013
R64019 vdd.n9198 vdd.n9197 0.013
R64020 vdd.n13282 vdd.n13281 0.013
R64021 vdd.n8976 vdd.n8975 0.013
R64022 vdd.n13574 vdd.n13573 0.013
R64023 vdd.n11608 vdd.n11605 0.013
R64024 vdd.n11620 vdd.n11619 0.013
R64025 vdd.n11951 vdd.n11542 0.013
R64026 vdd.n10181 vdd.n10082 0.013
R64027 vdd.n10449 vdd.n10287 0.013
R64028 vdd.n10303 vdd.n10302 0.013
R64029 vdd.n9339 vdd.n9334 0.013
R64030 vdd.n13037 vdd.n13036 0.013
R64031 vdd.n12942 vdd.n12941 0.013
R64032 vdd.n9534 vdd.n9530 0.013
R64033 vdd.n9699 vdd.n9694 0.013
R64034 vdd.n12829 vdd.n12828 0.013
R64035 vdd.n12734 vdd.n12733 0.013
R64036 vdd.n9895 vdd.n9891 0.013
R64037 vdd.n11893 vdd.n11797 0.013
R64038 vdd.n11918 vdd.n11663 0.013
R64039 vdd.n14331 vdd.n8354 0.013
R64040 vdd.n22324 vdd.n22323 0.013
R64041 vdd.n22309 vdd.n22308 0.013
R64042 vdd.n24324 vdd.n24323 0.013
R64043 vdd.n24296 vdd.n24295 0.013
R64044 vdd.n24281 vdd.n24280 0.013
R64045 vdd.n24207 vdd.n24206 0.013
R64046 vdd.n24146 vdd.n24136 0.013
R64047 vdd.n24038 vdd.n24036 0.013
R64048 vdd.n23914 vdd.n23904 0.013
R64049 vdd.n23806 vdd.n23804 0.013
R64050 vdd.n23682 vdd.n23672 0.013
R64051 vdd.n23118 vdd.n23116 0.013
R64052 vdd.n23226 vdd.n23216 0.013
R64053 vdd.n23350 vdd.n23348 0.013
R64054 vdd.n23458 vdd.n23448 0.013
R64055 vdd.n23582 vdd.n23580 0.013
R64056 vdd.n22539 vdd.n22537 0.013
R64057 vdd.n22647 vdd.n22637 0.013
R64058 vdd.n22771 vdd.n22769 0.013
R64059 vdd.n22879 vdd.n22869 0.013
R64060 vdd.n23003 vdd.n23001 0.013
R64061 vdd.n22468 vdd.n22467 0.013
R64062 vdd.n22453 vdd.n22452 0.013
R64063 vdd.n22379 vdd.n22378 0.013
R64064 vdd.n16951 vdd.n16937 0.013
R64065 vdd.n17029 vdd.n17028 0.013
R64066 vdd.n17223 vdd.n17209 0.013
R64067 vdd.n17301 vdd.n17300 0.013
R64068 vdd.n17495 vdd.n17481 0.013
R64069 vdd.n17573 vdd.n17572 0.013
R64070 vdd.n17753 vdd.n17739 0.013
R64071 vdd.n17831 vdd.n17830 0.013
R64072 vdd.n18024 vdd.n18010 0.013
R64073 vdd.n18102 vdd.n18101 0.013
R64074 vdd.n18291 vdd.n18278 0.013
R64075 vdd.n19134 vdd.n19132 0.013
R64076 vdd.n18910 vdd.n18908 0.013
R64077 vdd.n18876 vdd.n18874 0.013
R64078 vdd.n18651 vdd.n18649 0.013
R64079 vdd.n18617 vdd.n18615 0.013
R64080 vdd.n21019 vdd.n21017 0.013
R64081 vdd.n21647 vdd.n21646 0.013
R64082 vdd.n21651 vdd.n21649 0.013
R64083 vdd.n21535 vdd.n21533 0.013
R64084 vdd.n21501 vdd.n21499 0.013
R64085 vdd.n21276 vdd.n21274 0.013
R64086 vdd.n21242 vdd.n21240 0.013
R64087 vdd.n21697 vdd.n21696 0.013
R64088 vdd.n21693 vdd.n21692 0.013
R64089 vdd.n18425 vdd.n18424 0.013
R64090 vdd.n16717 vdd.n16708 0.013
R64091 vdd.n15308 vdd.n15294 0.013
R64092 vdd.n15329 vdd.n15328 0.013
R64093 vdd.n15536 vdd.n15519 0.013
R64094 vdd.n15563 vdd.n15562 0.013
R64095 vdd.n15792 vdd.n15775 0.013
R64096 vdd.n15819 vdd.n15818 0.013
R64097 vdd.n16048 vdd.n16031 0.013
R64098 vdd.n16075 vdd.n16074 0.013
R64099 vdd.n16304 vdd.n16287 0.013
R64100 vdd.n16331 vdd.n16330 0.013
R64101 vdd.n20694 vdd.n20692 0.013
R64102 vdd.n21984 vdd.n21888 0.013
R64103 vdd.n22004 vdd.n21755 0.013
R64104 vdd.n24956 vdd.n24955 0.013
R64105 vdd.n69 vdd.n39 0.013
R64106 vdd.n5846 vdd.n5845 0.013
R64107 vdd.n24953 vdd.n24952 0.013
R64108 vdd.n24953 vdd.n24886 0.013
R64109 vdd.n403 vdd.n402 0.013
R64110 vdd.n31382 vdd.n31381 0.013
R64111 vdd.n25452 vdd.n25451 0.013
R64112 vdd.n28005 vdd.n27850 0.013
R64113 vdd.n30841 vdd.n30840 0.013
R64114 vdd.n25365 vdd.n25364 0.013
R64115 vdd.n30849 vdd.n30848 0.013
R64116 vdd.n29660 vdd.n29659 0.013
R64117 vdd.n29198 vdd.n29197 0.013
R64118 vdd.n30758 vdd.n30757 0.013
R64119 vdd.n30802 vdd.n30798 0.013
R64120 vdd.n26728 vdd.n26727 0.013
R64121 vdd.n26142 vdd.n26137 0.013
R64122 vdd.n30765 vdd.n30764 0.013
R64123 vdd.n30812 vdd.n30811 0.013
R64124 vdd.n30829 vdd.n30828 0.013
R64125 vdd.n30102 vdd.n30101 0.013
R64126 vdd.n30058 vdd.n30057 0.013
R64127 vdd.n29550 vdd.n29549 0.013
R64128 vdd.n29309 vdd.n29308 0.013
R64129 vdd.n29222 vdd.n29221 0.013
R64130 vdd.n29135 vdd.n29134 0.013
R64131 vdd.n26502 vdd.n26501 0.013
R64132 vdd.n26646 vdd.n26645 0.013
R64133 vdd.n26097 vdd.n26096 0.013
R64134 vdd.n26130 vdd.n26127 0.013
R64135 vdd.n26726 vdd.n26725 0.013
R64136 vdd.n29228 vdd.n29227 0.013
R64137 vdd.n26632 vdd.n26631 0.013
R64138 vdd.n26366 vdd.n26365 0.013
R64139 vdd.n29156 vdd.n29155 0.013
R64140 vdd.n29195 vdd.n29194 0.013
R64141 vdd.n29450 vdd.n29449 0.013
R64142 vdd.n29657 vdd.n29656 0.013
R64143 vdd.n29984 vdd.n29983 0.013
R64144 vdd.n30115 vdd.n30114 0.013
R64145 vdd.n32549 vdd.n32548 0.013
R64146 vdd.n30846 vdd.n30845 0.013
R64147 vdd.n26361 vdd.n26360 0.013
R64148 vdd.n26358 vdd.n26357 0.013
R64149 vdd.n26428 vdd.n26427 0.013
R64150 vdd.n26484 vdd.n26483 0.013
R64151 vdd.n29445 vdd.n29444 0.013
R64152 vdd.n29442 vdd.n29441 0.013
R64153 vdd.n29651 vdd.n29650 0.013
R64154 vdd.n29979 vdd.n29978 0.013
R64155 vdd.n32544 vdd.n32543 0.013
R64156 vdd.n32541 vdd.n32540 0.013
R64157 vdd.n30837 vdd.n30836 0.013
R64158 vdd.n30973 vdd.n30972 0.013
R64159 vdd.n29273 vdd.n29271 0.013
R64160 vdd.n29417 vdd.n29415 0.013
R64161 vdd.n29413 vdd.n29411 0.013
R64162 vdd.n32651 vdd.n32649 0.013
R64163 vdd.n32648 vdd.n32646 0.013
R64164 vdd.n32641 vdd.n32639 0.013
R64165 vdd.n29633 vdd.n29631 0.013
R64166 vdd.n29959 vdd.n29957 0.013
R64167 vdd.n30041 vdd.n30040 0.013
R64168 vdd.n30075 vdd.n30073 0.013
R64169 vdd.n31413 vdd.n31411 0.013
R64170 vdd.n31410 vdd.n31408 0.013
R64171 vdd.n30727 vdd.n30725 0.013
R64172 vdd.n29182 vdd.n29180 0.013
R64173 vdd.n29162 vdd.n29161 0.013
R64174 vdd.n29121 vdd.n29120 0.013
R64175 vdd.n29047 vdd.n29046 0.013
R64176 vdd.n29066 vdd.n29065 0.013
R64177 vdd.n29090 vdd.n29089 0.013
R64178 vdd.n26479 vdd.n26478 0.013
R64179 vdd.n26516 vdd.n26515 0.013
R64180 vdd.n26355 vdd.n26354 0.013
R64181 vdd.n26273 vdd.n26272 0.013
R64182 vdd.n26625 vdd.n26624 0.013
R64183 vdd.n26115 vdd.n26114 0.013
R64184 vdd.n26118 vdd.n26117 0.013
R64185 vdd.n30733 vdd.n30732 0.013
R64186 vdd.n29965 vdd.n29964 0.013
R64187 vdd.n24930 vdd.n24929 0.013
R64188 vdd.n25650 vdd.n25649 0.013
R64189 vdd.n25344 vdd.n25341 0.013
R64190 vdd.n27613 vdd.n27611 0.013
R64191 vdd.n27494 vdd.n27492 0.013
R64192 vdd.n27393 vdd.n27391 0.013
R64193 vdd.n25585 vdd.n25584 0.013
R64194 vdd.n34164 vdd.n34163 0.013
R64195 vdd.n34737 vdd.n34736 0.013
R64196 vdd.n5484 vdd.n5483 0.013
R64197 vdd.n4311 vdd.n4310 0.013
R64198 vdd.n1958 vdd.n1957 0.013
R64199 vdd.n2368 vdd.n2105 0.013
R64200 vdd.n24840 vdd.n24839 0.013
R64201 vdd.n24843 vdd.n24840 0.013
R64202 vdd.n24855 vdd.n24854 0.013
R64203 vdd.n24857 vdd.n24856 0.013
R64204 vdd.n24856 vdd.n24855 0.013
R64205 vdd.n24845 vdd.n24844 0.013
R64206 vdd.n24846 vdd.n24845 0.013
R64207 vdd.n24867 vdd.n24866 0.013
R64208 vdd.n24868 vdd.n24867 0.013
R64209 vdd.n24870 vdd.n24869 0.013
R64210 vdd.n24869 vdd.n24868 0.013
R64211 vdd.n24851 vdd.n24850 0.013
R64212 vdd.n24850 vdd.n24849 0.013
R64213 vdd.n24842 vdd.n24841 0.013
R64214 vdd.n24849 vdd.n24848 0.013
R64215 vdd.n24848 vdd.n24847 0.013
R64216 vdd.n22280 vdd.n22043 0.012
R64217 vdd.n26705 vdd.n26703 0.012
R64218 vdd.n31617 vdd.n31615 0.012
R64219 vdd.n30963 vdd.n30962 0.012
R64220 vdd.n26425 vdd.n26424 0.012
R64221 vdd.n33299 vdd.n33298 0.012
R64222 vdd.n33717 vdd.n33716 0.012
R64223 vdd.n913 vdd.n912 0.012
R64224 vdd.n655 vdd.n654 0.012
R64225 vdd.n35465 vdd.n35464 0.012
R64226 vdd.n32624 vdd.n32623 0.012
R64227 vdd.n31356 vdd.n31355 0.012
R64228 vdd.n31236 vdd.n31230 0.012
R64229 vdd.n33426 vdd.n33425 0.012
R64230 vdd.n33441 vdd.n33440 0.012
R64231 vdd.n33375 vdd.n33368 0.012
R64232 vdd.n33550 vdd.n33549 0.012
R64233 vdd.n33558 vdd.n33557 0.012
R64234 vdd.n33586 vdd.n33583 0.012
R64235 vdd.n33770 vdd.n33769 0.012
R64236 vdd.n33819 vdd.n33818 0.012
R64237 vdd.n34138 vdd.n34137 0.012
R64238 vdd.n35556 vdd.n35555 0.012
R64239 vdd.n35529 vdd.n35528 0.012
R64240 vdd.n35458 vdd.n35454 0.012
R64241 vdd.n35332 vdd.n35331 0.012
R64242 vdd.n1040 vdd.n995 0.012
R64243 vdd.n6020 vdd.n6019 0.012
R64244 vdd.n6011 vdd.n6010 0.012
R64245 vdd.n6131 vdd.n6130 0.012
R64246 vdd.n5912 vdd.n5911 0.012
R64247 vdd.n4574 vdd.n4573 0.012
R64248 vdd.n4565 vdd.n4564 0.012
R64249 vdd.n4322 vdd.n4321 0.012
R64250 vdd.n4443 vdd.n4439 0.012
R64251 vdd.n32474 vdd.n32421 0.012
R64252 vdd.n32138 vdd.n32136 0.012
R64253 vdd.n32166 vdd.n31575 0.012
R64254 vdd.n29713 vdd.n29711 0.012
R64255 vdd.n28870 vdd.n28865 0.012
R64256 vdd.n28005 vdd.n28004 0.012
R64257 vdd.n27988 vdd.n27973 0.012
R64258 vdd.n29790 vdd.n29787 0.012
R64259 vdd.n29767 vdd.n29741 0.012
R64260 vdd.n31006 vdd.n31005 0.012
R64261 vdd.n30955 vdd.n30954 0.012
R64262 vdd.n2497 vdd.n2491 0.012
R64263 vdd.n31827 vdd.n31709 0.012
R64264 vdd.n31686 vdd.n31685 0.012
R64265 vdd.n31690 vdd.n31686 0.012
R64266 vdd.n31852 vdd.n31695 0.012
R64267 vdd.n10142 vdd.n10088 0.012
R64268 vdd.n10206 vdd.n10093 0.012
R64269 vdd.n10233 vdd.n10073 0.012
R64270 vdd.n10549 vdd.n10548 0.012
R64271 vdd.n12449 vdd.n12448 0.012
R64272 vdd.n12408 vdd.n12407 0.012
R64273 vdd.n12346 vdd.n10810 0.012
R64274 vdd.n10892 vdd.n10891 0.012
R64275 vdd.n12247 vdd.n10991 0.012
R64276 vdd.n11042 vdd.n11039 0.012
R64277 vdd.n11153 vdd.n11151 0.012
R64278 vdd.n12109 vdd.n12108 0.012
R64279 vdd.n12040 vdd.n11319 0.012
R64280 vdd.n11401 vdd.n11400 0.012
R64281 vdd.n11507 vdd.n11503 0.012
R64282 vdd.n11591 vdd.n11590 0.012
R64283 vdd.n13957 vdd.n13956 0.012
R64284 vdd.n14015 vdd.n8585 0.012
R64285 vdd.n14247 vdd.n14246 0.012
R64286 vdd.n14305 vdd.n8365 0.012
R64287 vdd.n14543 vdd.n14537 0.012
R64288 vdd.n9084 vdd.n9083 0.012
R64289 vdd.n13432 vdd.n13431 0.012
R64290 vdd.n8864 vdd.n8863 0.012
R64291 vdd.n13724 vdd.n13723 0.012
R64292 vdd.n10399 vdd.n10332 0.012
R64293 vdd.n10361 vdd.n10352 0.012
R64294 vdd.n9428 vdd.n9404 0.012
R64295 vdd.n12979 vdd.n12978 0.012
R64296 vdd.n9602 vdd.n9601 0.012
R64297 vdd.n9642 vdd.n9641 0.012
R64298 vdd.n9788 vdd.n9764 0.012
R64299 vdd.n12771 vdd.n12770 0.012
R64300 vdd.n9962 vdd.n9961 0.012
R64301 vdd.n10002 vdd.n10001 0.012
R64302 vdd.n22294 vdd.n22293 0.012
R64303 vdd.n24339 vdd.n24338 0.012
R64304 vdd.n24266 vdd.n24265 0.012
R64305 vdd.n24222 vdd.n24221 0.012
R64306 vdd.n22438 vdd.n22437 0.012
R64307 vdd.n22394 vdd.n22393 0.012
R64308 vdd.n16705 vdd.n16703 0.012
R64309 vdd.n16734 vdd.n16733 0.012
R64310 vdd.n16588 vdd.n16587 0.012
R64311 vdd.n16904 vdd.n16903 0.012
R64312 vdd.n17076 vdd.n17062 0.012
R64313 vdd.n17176 vdd.n17175 0.012
R64314 vdd.n17348 vdd.n17334 0.012
R64315 vdd.n17448 vdd.n17447 0.012
R64316 vdd.n17606 vdd.n16819 0.012
R64317 vdd.n17706 vdd.n17705 0.012
R64318 vdd.n17877 vdd.n17864 0.012
R64319 vdd.n17977 vdd.n17976 0.012
R64320 vdd.n18149 vdd.n18135 0.012
R64321 vdd.n18247 vdd.n18246 0.012
R64322 vdd.n18333 vdd.n18331 0.012
R64323 vdd.n18406 vdd.n18405 0.012
R64324 vdd.n19051 vdd.n19039 0.012
R64325 vdd.n19004 vdd.n19002 0.012
R64326 vdd.n18792 vdd.n18780 0.012
R64327 vdd.n18745 vdd.n18743 0.012
R64328 vdd.n18533 vdd.n18521 0.012
R64329 vdd.n21417 vdd.n21405 0.012
R64330 vdd.n21370 vdd.n21368 0.012
R64331 vdd.n21158 vdd.n21146 0.012
R64332 vdd.n21111 vdd.n21109 0.012
R64333 vdd.n15414 vdd.n15401 0.012
R64334 vdd.n15433 vdd.n15432 0.012
R64335 vdd.n15664 vdd.n15649 0.012
R64336 vdd.n15686 vdd.n15685 0.012
R64337 vdd.n15920 vdd.n15905 0.012
R64338 vdd.n15942 vdd.n15941 0.012
R64339 vdd.n16176 vdd.n16161 0.012
R64340 vdd.n16198 vdd.n16197 0.012
R64341 vdd.n16432 vdd.n16417 0.012
R64342 vdd.n16454 vdd.n16453 0.012
R64343 vdd.n24553 vdd.n24551 0.012
R64344 vdd.n25051 vdd.n25050 0.012
R64345 vdd.n25258 vdd.n14975 0.012
R64346 vdd.n31386 vdd.n31385 0.012
R64347 vdd.n35313 vdd.n35312 0.012
R64348 vdd.n5865 vdd.n5864 0.012
R64349 vdd.n30006 vdd.n30005 0.012
R64350 vdd.n28129 vdd.n28128 0.012
R64351 vdd.n35179 vdd.n35178 0.012
R64352 vdd.n6315 vdd.n6314 0.012
R64353 vdd.n5100 vdd.n5099 0.012
R64354 vdd.n4182 vdd.n4181 0.012
R64355 vdd.n34017 vdd.n34016 0.012
R64356 vdd.n34604 vdd.n34603 0.012
R64357 vdd.n5351 vdd.n5350 0.012
R64358 vdd.n31243 vdd.n31242 0.012
R64359 vdd.n35180 vdd.n35179 0.012
R64360 vdd.n6316 vdd.n6315 0.012
R64361 vdd.n25999 vdd.n25998 0.012
R64362 vdd.n5101 vdd.n5100 0.012
R64363 vdd.n4183 vdd.n4182 0.012
R64364 vdd.n25916 vdd.n25914 0.012
R64365 vdd.n25814 vdd.n25812 0.012
R64366 vdd.n34018 vdd.n34017 0.012
R64367 vdd.n34605 vdd.n34604 0.012
R64368 vdd.n5352 vdd.n5351 0.012
R64369 vdd.n27660 vdd.n27659 0.011
R64370 vdd.n29086 vdd.n29084 0.011
R64371 vdd.n29743 vdd.n29742 0.011
R64372 vdd.n30946 vdd.n30945 0.011
R64373 vdd.n6128 vdd.n6127 0.011
R64374 vdd.n35452 vdd.n35451 0.011
R64375 vdd.n32812 vdd.n6386 0.011
R64376 vdd.n4661 vdd.n4655 0.011
R64377 vdd.n25631 vdd.n25630 0.011
R64378 vdd.n3955 vdd.n3775 0.011
R64379 vdd.n3938 vdd.n3788 0.011
R64380 vdd.n2558 vdd.n2408 0.011
R64381 vdd.n33298 vdd.n33297 0.011
R64382 vdd.n27583 vdd.n27582 0.011
R64383 vdd.n27660 vdd.n25356 0.011
R64384 vdd.n27660 vdd.n26228 0.011
R64385 vdd.n27660 vdd.n26582 0.011
R64386 vdd.n27660 vdd.n26720 0.011
R64387 vdd.n27660 vdd.n26581 0.011
R64388 vdd.n27660 vdd.n26559 0.011
R64389 vdd.n27660 vdd.n26417 0.011
R64390 vdd.n27660 vdd.n26558 0.011
R64391 vdd.n27660 vdd.n26537 0.011
R64392 vdd.n27660 vdd.n26536 0.011
R64393 vdd.n32737 vdd.n27683 0.011
R64394 vdd.n32737 vdd.n27724 0.011
R64395 vdd.n32737 vdd.n27725 0.011
R64396 vdd.n32737 vdd.n29040 0.011
R64397 vdd.n32737 vdd.n29145 0.011
R64398 vdd.n32737 vdd.n29175 0.011
R64399 vdd.n32737 vdd.n29215 0.011
R64400 vdd.n32737 vdd.n29249 0.011
R64401 vdd.n32737 vdd.n29267 0.011
R64402 vdd.n32737 vdd.n29268 0.011
R64403 vdd.n32737 vdd.n29368 0.011
R64404 vdd.n32737 vdd.n29369 0.011
R64405 vdd.n32737 vdd.n29391 0.011
R64406 vdd.n32737 vdd.n29473 0.011
R64407 vdd.n32737 vdd.n29494 0.011
R64408 vdd.n32737 vdd.n32736 0.011
R64409 vdd.n32737 vdd.n29562 0.011
R64410 vdd.n32737 vdd.n29589 0.011
R64411 vdd.n32737 vdd.n29611 0.011
R64412 vdd.n32737 vdd.n32735 0.011
R64413 vdd.n32737 vdd.n32712 0.011
R64414 vdd.n32737 vdd.n32734 0.011
R64415 vdd.n32737 vdd.n32635 0.011
R64416 vdd.n32737 vdd.n32617 0.011
R64417 vdd.n32737 vdd.n30014 0.011
R64418 vdd.n32737 vdd.n30036 0.011
R64419 vdd.n32737 vdd.n30069 0.011
R64420 vdd.n32737 vdd.n30134 0.011
R64421 vdd.n32737 vdd.n32616 0.011
R64422 vdd.n32737 vdd.n32594 0.011
R64423 vdd.n32737 vdd.n32615 0.011
R64424 vdd.n32737 vdd.n32572 0.011
R64425 vdd.n32737 vdd.n31404 0.011
R64426 vdd.n32737 vdd.n30870 0.011
R64427 vdd.n32737 vdd.n30721 0.011
R64428 vdd.n32737 vdd.n30893 0.011
R64429 vdd.n32737 vdd.n30916 0.011
R64430 vdd.n32737 vdd.n31403 0.011
R64431 vdd.n32737 vdd.n31365 0.011
R64432 vdd.n32737 vdd.n31402 0.011
R64433 vdd.n32737 vdd.n31348 0.011
R64434 vdd.n32737 vdd.n31328 0.011
R64435 vdd.n32737 vdd.n31327 0.011
R64436 vdd.n654 vdd.n653 0.011
R64437 vdd.n33507 vdd.n33504 0.011
R64438 vdd.n33508 vdd.n33507 0.011
R64439 vdd.n33497 vdd.n33496 0.011
R64440 vdd.n33322 vdd.n33320 0.011
R64441 vdd.n33361 vdd.n33360 0.011
R64442 vdd.n33558 vdd.n33554 0.011
R64443 vdd.n33324 vdd.n33323 0.011
R64444 vdd.n33709 vdd.n33708 0.011
R64445 vdd.n33773 vdd.n33710 0.011
R64446 vdd.n33658 vdd.n33656 0.011
R64447 vdd.n33685 vdd.n33684 0.011
R64448 vdd.n33751 vdd.n33748 0.011
R64449 vdd.n33625 vdd.n33624 0.011
R64450 vdd.n33851 vdd.n33850 0.011
R64451 vdd.n34082 vdd.n34081 0.011
R64452 vdd.n34092 vdd.n34091 0.011
R64453 vdd.n34297 vdd.n34295 0.011
R64454 vdd.n34326 vdd.n34325 0.011
R64455 vdd.n34138 vdd.n34133 0.011
R64456 vdd.n33927 vdd.n33926 0.011
R64457 vdd.n33898 vdd.n33893 0.011
R64458 vdd.n33881 vdd.n33880 0.011
R64459 vdd.n33952 vdd.n33950 0.011
R64460 vdd.n33950 vdd.n33947 0.011
R64461 vdd.n33871 vdd.n33870 0.011
R64462 vdd.n34351 vdd.n34350 0.011
R64463 vdd.n33945 vdd.n33944 0.011
R64464 vdd.n35563 vdd.n35561 0.011
R64465 vdd.n35253 vdd.n35252 0.011
R64466 vdd.n35241 vdd.n35240 0.011
R64467 vdd.n35592 vdd.n35591 0.011
R64468 vdd.n35476 vdd.n35475 0.011
R64469 vdd.n35491 vdd.n35490 0.011
R64470 vdd.n35122 vdd.n35121 0.011
R64471 vdd.n35106 vdd.n35105 0.011
R64472 vdd.n35038 vdd.n35036 0.011
R64473 vdd.n35036 vdd.n35033 0.011
R64474 vdd.n35092 vdd.n35087 0.011
R64475 vdd.n35053 vdd.n35052 0.011
R64476 vdd.n35369 vdd.n35368 0.011
R64477 vdd.n35096 vdd.n35095 0.011
R64478 vdd.n35114 vdd.n35113 0.011
R64479 vdd.n35429 vdd.n35428 0.011
R64480 vdd.n35305 vdd.n35304 0.011
R64481 vdd.n34654 vdd.n34653 0.011
R64482 vdd.n34669 vdd.n34668 0.011
R64483 vdd.n34913 vdd.n34911 0.011
R64484 vdd.n35005 vdd.n35004 0.011
R64485 vdd.n34466 vdd.n34465 0.011
R64486 vdd.n34505 vdd.n34500 0.011
R64487 vdd.n34519 vdd.n34518 0.011
R64488 vdd.n34454 vdd.n34452 0.011
R64489 vdd.n34452 vdd.n34449 0.011
R64490 vdd.n34535 vdd.n34534 0.011
R64491 vdd.n34779 vdd.n34778 0.011
R64492 vdd.n34509 vdd.n34508 0.011
R64493 vdd.n1031 vdd.n1028 0.011
R64494 vdd.n1032 vdd.n1031 0.011
R64495 vdd.n987 vdd.n986 0.011
R64496 vdd.n632 vdd.n630 0.011
R64497 vdd.n1040 vdd.n1039 0.011
R64498 vdd.n792 vdd.n788 0.011
R64499 vdd.n879 vdd.n874 0.011
R64500 vdd.n1074 vdd.n1072 0.011
R64501 vdd.n944 vdd.n943 0.011
R64502 vdd.n532 vdd.n530 0.011
R64503 vdd.n571 vdd.n570 0.011
R64504 vdd.n5 vdd.n4 0.011
R64505 vdd.n14 vdd.n13 0.011
R64506 vdd.n47 vdd.n42 0.011
R64507 vdd.n226 vdd.n225 0.011
R64508 vdd.n255 vdd.n254 0.011
R64509 vdd.n247 vdd.n246 0.011
R64510 vdd.n248 vdd.n247 0.011
R64511 vdd.n100 vdd.n97 0.011
R64512 vdd.n118 vdd.n117 0.011
R64513 vdd.n5956 vdd.n5954 0.011
R64514 vdd.n5797 vdd.n5796 0.011
R64515 vdd.n5784 vdd.n5783 0.011
R64516 vdd.n6028 vdd.n6027 0.011
R64517 vdd.n5830 vdd.n5829 0.011
R64518 vdd.n6145 vdd.n6144 0.011
R64519 vdd.n6155 vdd.n6154 0.011
R64520 vdd.n6236 vdd.n6234 0.011
R64521 vdd.n6234 vdd.n6231 0.011
R64522 vdd.n6172 vdd.n6167 0.011
R64523 vdd.n6201 vdd.n6200 0.011
R64524 vdd.n6057 vdd.n6056 0.011
R64525 vdd.n6247 vdd.n6149 0.011
R64526 vdd.n6205 vdd.n6204 0.011
R64527 vdd.n6229 vdd.n6228 0.011
R64528 vdd.n5874 vdd.n5873 0.011
R64529 vdd.n5401 vdd.n5400 0.011
R64530 vdd.n5416 vdd.n5415 0.011
R64531 vdd.n5660 vdd.n5658 0.011
R64532 vdd.n5752 vdd.n5751 0.011
R64533 vdd.n5213 vdd.n5212 0.011
R64534 vdd.n5252 vdd.n5247 0.011
R64535 vdd.n5266 vdd.n5265 0.011
R64536 vdd.n5201 vdd.n5199 0.011
R64537 vdd.n5199 vdd.n5196 0.011
R64538 vdd.n5282 vdd.n5281 0.011
R64539 vdd.n5526 vdd.n5525 0.011
R64540 vdd.n5256 vdd.n5255 0.011
R64541 vdd.n4642 vdd.n4640 0.011
R64542 vdd.n5095 vdd.n5094 0.011
R64543 vdd.n5082 vdd.n5081 0.011
R64544 vdd.n4818 vdd.n4817 0.011
R64545 vdd.n4826 vdd.n4825 0.011
R64546 vdd.n4849 vdd.n4848 0.011
R64547 vdd.n4795 vdd.n4794 0.011
R64548 vdd.n5002 vdd.n5001 0.011
R64549 vdd.n4980 vdd.n4975 0.011
R64550 vdd.n5040 vdd.n5037 0.011
R64551 vdd.n5042 vdd.n5040 0.011
R64552 vdd.n4964 vdd.n4963 0.011
R64553 vdd.n4957 vdd.n4956 0.011
R64554 vdd.n5035 vdd.n5034 0.011
R64555 vdd.n4692 vdd.n4691 0.011
R64556 vdd.n4231 vdd.n4230 0.011
R64557 vdd.n4246 vdd.n4245 0.011
R64558 vdd.n4487 vdd.n4485 0.011
R64559 vdd.n4543 vdd.n4527 0.011
R64560 vdd.n4582 vdd.n4581 0.011
R64561 vdd.n4540 vdd.n4539 0.011
R64562 vdd.n4295 vdd.n4294 0.011
R64563 vdd.n4043 vdd.n4042 0.011
R64564 vdd.n4082 vdd.n4077 0.011
R64565 vdd.n4096 vdd.n4095 0.011
R64566 vdd.n4031 vdd.n4029 0.011
R64567 vdd.n4029 vdd.n4026 0.011
R64568 vdd.n4112 vdd.n4111 0.011
R64569 vdd.n4353 vdd.n4352 0.011
R64570 vdd.n4086 vdd.n4085 0.011
R64571 vdd.n4104 vdd.n4103 0.011
R64572 vdd.n4406 vdd.n4405 0.011
R64573 vdd.n27226 vdd.n27225 0.011
R64574 vdd.n29946 vdd.n29943 0.011
R64575 vdd.n27753 vdd.n27749 0.011
R64576 vdd.n28972 vdd.n28971 0.011
R64577 vdd.n28838 vdd.n28806 0.011
R64578 vdd.n28882 vdd.n28877 0.011
R64579 vdd.n28897 vdd.n28892 0.011
R64580 vdd.n28910 vdd.n28905 0.011
R64581 vdd.n29017 vdd.n28048 0.011
R64582 vdd.n28029 vdd.n28028 0.011
R64583 vdd.n28026 vdd.n28023 0.011
R64584 vdd.n28014 vdd.n28013 0.011
R64585 vdd.n27996 vdd.n27995 0.011
R64586 vdd.n27966 vdd.n27964 0.011
R64587 vdd.n27957 vdd.n27956 0.011
R64588 vdd.n29802 vdd.n29799 0.011
R64589 vdd.n29783 vdd.n29782 0.011
R64590 vdd.n29781 vdd.n29778 0.011
R64591 vdd.n29774 vdd.n29773 0.011
R64592 vdd.n29733 vdd.n29732 0.011
R64593 vdd.n30670 vdd.n30665 0.011
R64594 vdd.n30690 vdd.n30652 0.011
R64595 vdd.n30644 vdd.n30643 0.011
R64596 vdd.n27278 vdd.n27274 0.011
R64597 vdd.n27555 vdd.n27550 0.011
R64598 vdd.n27576 vdd.n27575 0.011
R64599 vdd.n27563 vdd.n27561 0.011
R64600 vdd.n27561 vdd.n27559 0.011
R64601 vdd.n27589 vdd.n27588 0.011
R64602 vdd.n27301 vdd.n27297 0.011
R64603 vdd.n27374 vdd.n27373 0.011
R64604 vdd.n27434 vdd.n27432 0.011
R64605 vdd.n25724 vdd.n25720 0.011
R64606 vdd.n25992 vdd.n25987 0.011
R64607 vdd.n25689 vdd.n25688 0.011
R64608 vdd.n25699 vdd.n25697 0.011
R64609 vdd.n25697 vdd.n25695 0.011
R64610 vdd.n26005 vdd.n26004 0.011
R64611 vdd.n25753 vdd.n25749 0.011
R64612 vdd.n25742 vdd.n25741 0.011
R64613 vdd.n25880 vdd.n25878 0.011
R64614 vdd.n25657 vdd.n25654 0.011
R64615 vdd.n25579 vdd.n25574 0.011
R64616 vdd.n25472 vdd.n25471 0.011
R64617 vdd.n30881 vdd.n30879 0.011
R64618 vdd.n29576 vdd.n29574 0.011
R64619 vdd.n29477 vdd.n29476 0.011
R64620 vdd.n29479 vdd.n29478 0.011
R64621 vdd.n27671 vdd.n27669 0.011
R64622 vdd.n26424 vdd.n26422 0.011
R64623 vdd.n26513 vdd.n26512 0.011
R64624 vdd.n25372 vdd.n25371 0.011
R64625 vdd.n29086 vdd.n29085 0.011
R64626 vdd.n32658 vdd.n32657 0.011
R64627 vdd.n30749 vdd.n30748 0.011
R64628 vdd.n4021 vdd.n4020 0.011
R64629 vdd.n3914 vdd.n3911 0.011
R64630 vdd.n2660 vdd.n2577 0.011
R64631 vdd.n3680 vdd.n3679 0.011
R64632 vdd.n4015 vdd.n4013 0.011
R64633 vdd.n3858 vdd.n3855 0.011
R64634 vdd.n2241 vdd.n2233 0.011
R64635 vdd.n2257 vdd.n2256 0.011
R64636 vdd.n2298 vdd.n2297 0.011
R64637 vdd.n2514 vdd.n2511 0.011
R64638 vdd.n2500 vdd.n2497 0.011
R64639 vdd.n2483 vdd.n2480 0.011
R64640 vdd.n2624 vdd.n2616 0.011
R64641 vdd.n2656 vdd.n2648 0.011
R64642 vdd.n1993 vdd.n1991 0.011
R64643 vdd.n1802 vdd.n1799 0.011
R64644 vdd.n1784 vdd.n1783 0.011
R64645 vdd.n2082 vdd.n2081 0.011
R64646 vdd.n26403 vdd.n26402 0.011
R64647 vdd.n31808 vdd.n31718 0.011
R64648 vdd.n26620 vdd.n26612 0.011
R64649 vdd.n26706 vdd.n26686 0.011
R64650 vdd.n31872 vdd.n31869 0.011
R64651 vdd.n31942 vdd.n31939 0.011
R64652 vdd.n31972 vdd.n31967 0.011
R64653 vdd.n31986 vdd.n31981 0.011
R64654 vdd.n32034 vdd.n32031 0.011
R64655 vdd.n32236 vdd.n32233 0.011
R64656 vdd.n32303 vdd.n32300 0.011
R64657 vdd.n31124 vdd.n31121 0.011
R64658 vdd.n32013 vdd.n32012 0.011
R64659 vdd.n32185 vdd.n32184 0.011
R64660 vdd.n32245 vdd.n32244 0.011
R64661 vdd.n32277 vdd.n32276 0.011
R64662 vdd.n32300 vdd.n32299 0.011
R64663 vdd.n12508 vdd.n12507 0.011
R64664 vdd.n10641 vdd.n10640 0.011
R64665 vdd.n10733 vdd.n10732 0.011
R64666 vdd.n12359 vdd.n12358 0.011
R64667 vdd.n12300 vdd.n10893 0.011
R64668 vdd.n10990 vdd.n10965 0.011
R64669 vdd.n11081 vdd.n11062 0.011
R64670 vdd.n11157 vdd.n11131 0.011
R64671 vdd.n12096 vdd.n11224 0.011
R64672 vdd.n12053 vdd.n12052 0.011
R64673 vdd.n11994 vdd.n11402 0.011
R64674 vdd.n11499 vdd.n11498 0.011
R64675 vdd.n11499 vdd.n11435 0.011
R64676 vdd.n11595 vdd.n11587 0.011
R64677 vdd.n13883 vdd.n8700 0.011
R64678 vdd.n8547 vdd.n8529 0.011
R64679 vdd.n14172 vdd.n8477 0.011
R64680 vdd.n14387 vdd.n14386 0.011
R64681 vdd.n14447 vdd.n14446 0.011
R64682 vdd.n8760 vdd.n8742 0.011
R64683 vdd.n13224 vdd.n13223 0.011
R64684 vdd.n13309 vdd.n9136 0.011
R64685 vdd.n13516 vdd.n13515 0.011
R64686 vdd.n13601 vdd.n8914 0.011
R64687 vdd.n11589 vdd.n11588 0.011
R64688 vdd.n10180 vdd.n10177 0.011
R64689 vdd.n10461 vdd.n10460 0.011
R64690 vdd.n10435 vdd.n10434 0.011
R64691 vdd.n13053 vdd.n9311 0.011
R64692 vdd.n9377 vdd.n9372 0.011
R64693 vdd.n9512 vdd.n9506 0.011
R64694 vdd.n12925 vdd.n9547 0.011
R64695 vdd.n12845 vdd.n9672 0.011
R64696 vdd.n9737 vdd.n9732 0.011
R64697 vdd.n9872 vdd.n9866 0.011
R64698 vdd.n12717 vdd.n9907 0.011
R64699 vdd.n12637 vdd.n10032 0.011
R64700 vdd.n11916 vdd.n11915 0.011
R64701 vdd.n13298 vdd.n13293 0.011
R64702 vdd.n13296 vdd.n9100 0.011
R64703 vdd.n13343 vdd.n13342 0.011
R64704 vdd.n13370 vdd.n9066 0.011
R64705 vdd.n13398 vdd.n13397 0.011
R64706 vdd.n13396 vdd.n9039 0.011
R64707 vdd.n13419 vdd.n13416 0.011
R64708 vdd.n13488 vdd.n8998 0.011
R64709 vdd.n13486 vdd.n8999 0.011
R64710 vdd.n13502 vdd.n8985 0.011
R64711 vdd.n13505 vdd.n13503 0.011
R64712 vdd.n13543 vdd.n13542 0.011
R64713 vdd.n13563 vdd.n8941 0.011
R64714 vdd.n13565 vdd.n8926 0.011
R64715 vdd.n13590 vdd.n13585 0.011
R64716 vdd.n13588 vdd.n8879 0.011
R64717 vdd.n13635 vdd.n13634 0.011
R64718 vdd.n13662 vdd.n8846 0.011
R64719 vdd.n13688 vdd.n8818 0.011
R64720 vdd.n13712 vdd.n13710 0.011
R64721 vdd.n13768 vdd.n8781 0.011
R64722 vdd.n13766 vdd.n8782 0.011
R64723 vdd.n13782 vdd.n8770 0.011
R64724 vdd.n13786 vdd.n13783 0.011
R64725 vdd.n13828 vdd.n13827 0.011
R64726 vdd.n13845 vdd.n8725 0.011
R64727 vdd.n13853 vdd.n13852 0.011
R64728 vdd.n13894 vdd.n8687 0.011
R64729 vdd.n13892 vdd.n8688 0.011
R64730 vdd.n13910 vdd.n13909 0.011
R64731 vdd.n13983 vdd.n13982 0.011
R64732 vdd.n13986 vdd.n13984 0.011
R64733 vdd.n14058 vdd.n8570 0.011
R64734 vdd.n14056 vdd.n8571 0.011
R64735 vdd.n14045 vdd.n14044 0.011
R64736 vdd.n14075 vdd.n14074 0.011
R64737 vdd.n14114 vdd.n8517 0.011
R64738 vdd.n14111 vdd.n8520 0.011
R64739 vdd.n14134 vdd.n8504 0.011
R64740 vdd.n14142 vdd.n14141 0.011
R64741 vdd.n14183 vdd.n8463 0.011
R64742 vdd.n14181 vdd.n8465 0.011
R64743 vdd.n14200 vdd.n14199 0.011
R64744 vdd.n8447 vdd.n8446 0.011
R64745 vdd.n14273 vdd.n14272 0.011
R64746 vdd.n14276 vdd.n14274 0.011
R64747 vdd.n14333 vdd.n8353 0.011
R64748 vdd.n24354 vdd.n24353 0.011
R64749 vdd.n24251 vdd.n24250 0.011
R64750 vdd.n24237 vdd.n24236 0.011
R64751 vdd.n24136 vdd.n24134 0.011
R64752 vdd.n24040 vdd.n24038 0.011
R64753 vdd.n23904 vdd.n23902 0.011
R64754 vdd.n23808 vdd.n23806 0.011
R64755 vdd.n23672 vdd.n23670 0.011
R64756 vdd.n23120 vdd.n23118 0.011
R64757 vdd.n23216 vdd.n23214 0.011
R64758 vdd.n23352 vdd.n23350 0.011
R64759 vdd.n23448 vdd.n23446 0.011
R64760 vdd.n23584 vdd.n23582 0.011
R64761 vdd.n22541 vdd.n22539 0.011
R64762 vdd.n22637 vdd.n22635 0.011
R64763 vdd.n22773 vdd.n22771 0.011
R64764 vdd.n22869 vdd.n22867 0.011
R64765 vdd.n23005 vdd.n23003 0.011
R64766 vdd.n22423 vdd.n22422 0.011
R64767 vdd.n22409 vdd.n22408 0.011
R64768 vdd.n24369 vdd.n24368 0.011
R64769 vdd.n16935 vdd.n16921 0.011
R64770 vdd.n17045 vdd.n17044 0.011
R64771 vdd.n17207 vdd.n17193 0.011
R64772 vdd.n17317 vdd.n17316 0.011
R64773 vdd.n17479 vdd.n17465 0.011
R64774 vdd.n17589 vdd.n17588 0.011
R64775 vdd.n17737 vdd.n17723 0.011
R64776 vdd.n17847 vdd.n17846 0.011
R64777 vdd.n18008 vdd.n17994 0.011
R64778 vdd.n18118 vdd.n18117 0.011
R64779 vdd.n18276 vdd.n18263 0.011
R64780 vdd.n18318 vdd.n18317 0.011
R64781 vdd.n18330 vdd.n18318 0.011
R64782 vdd.n18414 vdd.n18408 0.011
R64783 vdd.n19119 vdd.n19117 0.011
R64784 vdd.n18926 vdd.n18924 0.011
R64785 vdd.n18860 vdd.n18858 0.011
R64786 vdd.n18667 vdd.n18665 0.011
R64787 vdd.n18601 vdd.n18599 0.011
R64788 vdd.n21033 vdd.n21031 0.011
R64789 vdd.n21551 vdd.n21549 0.011
R64790 vdd.n21485 vdd.n21483 0.011
R64791 vdd.n21292 vdd.n21290 0.011
R64792 vdd.n21226 vdd.n21224 0.011
R64793 vdd.n18429 vdd.n18428 0.011
R64794 vdd.n16774 vdd.n16773 0.011
R64795 vdd.n15292 vdd.n15280 0.011
R64796 vdd.n15343 vdd.n15342 0.011
R64797 vdd.n15517 vdd.n15502 0.011
R64798 vdd.n15580 vdd.n15579 0.011
R64799 vdd.n15773 vdd.n15758 0.011
R64800 vdd.n15836 vdd.n15835 0.011
R64801 vdd.n16029 vdd.n16014 0.011
R64802 vdd.n16092 vdd.n16091 0.011
R64803 vdd.n16285 vdd.n16270 0.011
R64804 vdd.n16348 vdd.n16347 0.011
R64805 vdd.n16541 vdd.n16526 0.011
R64806 vdd.n19485 vdd.n19483 0.011
R64807 vdd.n19500 vdd.n19499 0.011
R64808 vdd.n19516 vdd.n19514 0.011
R64809 vdd.n19519 vdd.n19517 0.011
R64810 vdd.n19530 vdd.n19529 0.011
R64811 vdd.n19544 vdd.n19532 0.011
R64812 vdd.n19560 vdd.n19548 0.011
R64813 vdd.n19576 vdd.n19564 0.011
R64814 vdd.n19592 vdd.n19580 0.011
R64815 vdd.n19608 vdd.n19596 0.011
R64816 vdd.n19624 vdd.n19609 0.011
R64817 vdd.n19639 vdd.n19638 0.011
R64818 vdd.n19653 vdd.n19651 0.011
R64819 vdd.n19669 vdd.n19667 0.011
R64820 vdd.n19685 vdd.n19683 0.011
R64821 vdd.n19701 vdd.n19699 0.011
R64822 vdd.n19717 vdd.n19715 0.011
R64823 vdd.n19720 vdd.n19718 0.011
R64824 vdd.n19746 vdd.n19734 0.011
R64825 vdd.n19762 vdd.n19750 0.011
R64826 vdd.n19778 vdd.n19766 0.011
R64827 vdd.n19794 vdd.n19782 0.011
R64828 vdd.n19810 vdd.n19798 0.011
R64829 vdd.n19826 vdd.n19811 0.011
R64830 vdd.n19831 vdd.n19830 0.011
R64831 vdd.n20996 vdd.n20995 0.011
R64832 vdd.n20991 vdd.n20979 0.011
R64833 vdd.n20975 vdd.n20963 0.011
R64834 vdd.n20959 vdd.n20947 0.011
R64835 vdd.n20943 vdd.n20931 0.011
R64836 vdd.n20917 vdd.n20915 0.011
R64837 vdd.n20914 vdd.n20912 0.011
R64838 vdd.n20898 vdd.n20896 0.011
R64839 vdd.n20882 vdd.n20880 0.011
R64840 vdd.n20866 vdd.n20864 0.011
R64841 vdd.n20861 vdd.n20859 0.011
R64842 vdd.n20847 vdd.n20846 0.011
R64843 vdd.n20829 vdd.n20817 0.011
R64844 vdd.n20816 vdd.n20804 0.011
R64845 vdd.n20800 vdd.n20788 0.011
R64846 vdd.n20784 vdd.n20772 0.011
R64847 vdd.n20769 vdd.n20757 0.011
R64848 vdd.n20753 vdd.n20741 0.011
R64849 vdd.n20739 vdd.n20738 0.011
R64850 vdd.n20728 vdd.n20726 0.011
R64851 vdd.n20725 vdd.n20723 0.011
R64852 vdd.n20709 vdd.n20708 0.011
R64853 vdd.n22002 vdd.n22001 0.011
R64854 vdd.n25048 vdd.n25047 0.011
R64855 vdd.n30975 vdd.n30956 0.011
R64856 vdd.n26241 vdd.n26239 0.011
R64857 vdd.n29380 vdd.n29378 0.011
R64858 vdd.n32605 vdd.n32603 0.011
R64859 vdd.n27470 vdd.n27468 0.011
R64860 vdd.n27362 vdd.n27360 0.011
R64861 vdd.n25553 vdd.n25552 0.011
R64862 vdd.n25467 vdd.n25466 0.011
R64863 vdd.n31247 vdd.n31241 0.011
R64864 vdd.n31337 vdd.n31336 0.011
R64865 vdd.n32738 vdd.n7152 0.011
R64866 vdd.n35464 vdd.n35463 0.011
R64867 vdd.n2098 vdd.n2097 0.011
R64868 vdd.n33708 vdd.n33704 0.011
R64869 vdd.n795 vdd.n792 0.011
R64870 vdd.n233 vdd.n232 0.011
R64871 vdd.n7116 vdd.n7115 0.011
R64872 vdd.n11905 vdd.n11789 0.011
R64873 vdd.n21996 vdd.n21880 0.011
R64874 vdd.n402 vdd.n401 0.01
R64875 vdd.n6892 vdd.n6891 0.01
R64876 vdd.n6862 vdd.n6861 0.01
R64877 vdd.n6808 vdd.n6807 0.01
R64878 vdd.n6748 vdd.n6747 0.01
R64879 vdd.n6695 vdd.n6694 0.01
R64880 vdd.n6638 vdd.n6637 0.01
R64881 vdd.n6580 vdd.n6579 0.01
R64882 vdd.n6524 vdd.n6523 0.01
R64883 vdd.n6470 vdd.n6469 0.01
R64884 vdd.n6408 vdd.n6407 0.01
R64885 vdd.n31222 vdd.n31221 0.01
R64886 vdd.n32468 vdd.n32425 0.01
R64887 vdd.n32185 vdd.n31564 0.01
R64888 vdd.n34232 vdd.n34231 0.01
R64889 vdd.n26511 vdd.n26510 0.01
R64890 vdd.n4907 vdd.n4906 0.01
R64891 vdd.n2877 vdd.n2870 0.01
R64892 vdd.n2911 vdd.n2909 0.01
R64893 vdd.n3058 vdd.n3051 0.01
R64894 vdd.n3092 vdd.n3090 0.01
R64895 vdd.n3239 vdd.n3232 0.01
R64896 vdd.n3273 vdd.n3271 0.01
R64897 vdd.n3420 vdd.n3413 0.01
R64898 vdd.n3454 vdd.n3452 0.01
R64899 vdd.n3601 vdd.n3594 0.01
R64900 vdd.n33459 vdd.n33457 0.01
R64901 vdd.n33364 vdd.n33363 0.01
R64902 vdd.n33699 vdd.n33698 0.01
R64903 vdd.n34341 vdd.n34340 0.01
R64904 vdd.n34338 vdd.n34337 0.01
R64905 vdd.n34131 vdd.n34130 0.01
R64906 vdd.n34220 vdd.n34219 0.01
R64907 vdd.n34171 vdd.n34170 0.01
R64908 vdd.n34181 vdd.n34180 0.01
R64909 vdd.n33962 vdd.n33875 0.01
R64910 vdd.n34404 vdd.n34403 0.01
R64911 vdd.n33962 vdd.n33961 0.01
R64912 vdd.n34408 vdd.n34407 0.01
R64913 vdd.n34419 vdd.n34418 0.01
R64914 vdd.n34068 vdd.n34066 0.01
R64915 vdd.n34019 vdd.n34018 0.01
R64916 vdd.n34048 vdd.n34047 0.01
R64917 vdd.n35608 vdd.n35607 0.01
R64918 vdd.n35229 vdd.n35227 0.01
R64919 vdd.n35020 vdd.n35019 0.01
R64920 vdd.n34966 vdd.n34953 0.01
R64921 vdd.n34966 vdd.n34965 0.01
R64922 vdd.n34721 vdd.n34720 0.01
R64923 vdd.n34740 vdd.n34739 0.01
R64924 vdd.n34527 vdd.n34513 0.01
R64925 vdd.n34831 vdd.n34830 0.01
R64926 vdd.n34852 vdd.n34851 0.01
R64927 vdd.n34527 vdd.n34526 0.01
R64928 vdd.n34833 vdd.n34832 0.01
R64929 vdd.n34642 vdd.n34640 0.01
R64930 vdd.n34606 vdd.n34605 0.01
R64931 vdd.n34623 vdd.n34622 0.01
R64932 vdd.n778 vdd.n776 0.01
R64933 vdd.n683 vdd.n682 0.01
R64934 vdd.n625 vdd.n624 0.01
R64935 vdd.n662 vdd.n661 0.01
R64936 vdd.n1166 vdd.n1165 0.01
R64937 vdd.n1093 vdd.n1092 0.01
R64938 vdd.n1127 vdd.n1126 0.01
R64939 vdd.n546 vdd.n545 0.01
R64940 vdd.n548 vdd.n547 0.01
R64941 vdd.n574 vdd.n573 0.01
R64942 vdd.n473 vdd.n471 0.01
R64943 vdd.n75 vdd.n71 0.01
R64944 vdd.n75 vdd.n74 0.01
R64945 vdd.n204 vdd.n201 0.01
R64946 vdd.n138 vdd.n137 0.01
R64947 vdd.n282 vdd.n278 0.01
R64948 vdd.n147 vdd.n146 0.01
R64949 vdd.n6043 vdd.n6042 0.01
R64950 vdd.n6346 vdd.n6345 0.01
R64951 vdd.n6352 vdd.n6350 0.01
R64952 vdd.n5767 vdd.n5766 0.01
R64953 vdd.n5713 vdd.n5700 0.01
R64954 vdd.n5713 vdd.n5712 0.01
R64955 vdd.n5468 vdd.n5467 0.01
R64956 vdd.n5487 vdd.n5486 0.01
R64957 vdd.n5274 vdd.n5260 0.01
R64958 vdd.n5578 vdd.n5577 0.01
R64959 vdd.n5599 vdd.n5598 0.01
R64960 vdd.n5274 vdd.n5273 0.01
R64961 vdd.n5580 vdd.n5579 0.01
R64962 vdd.n5389 vdd.n5387 0.01
R64963 vdd.n5353 vdd.n5352 0.01
R64964 vdd.n5370 vdd.n5369 0.01
R64965 vdd.n5165 vdd.n5164 0.01
R64966 vdd.n5102 vdd.n5101 0.01
R64967 vdd.n4856 vdd.n4851 0.01
R64968 vdd.n4856 vdd.n4855 0.01
R64969 vdd.n5183 vdd.n5181 0.01
R64970 vdd.n4769 vdd.n4768 0.01
R64971 vdd.n5054 vdd.n5050 0.01
R64972 vdd.n5054 vdd.n5053 0.01
R64973 vdd.n4707 vdd.n4706 0.01
R64974 vdd.n4926 vdd.n4925 0.01
R64975 vdd.n4597 vdd.n4596 0.01
R64976 vdd.n4219 vdd.n4217 0.01
R64977 vdd.n36019 vdd.n36009 0.01
R64978 vdd.n36063 vdd.n36061 0.01
R64979 vdd.n36250 vdd.n36240 0.01
R64980 vdd.n36294 vdd.n36292 0.01
R64981 vdd.n36481 vdd.n36471 0.01
R64982 vdd.n36525 vdd.n36523 0.01
R64983 vdd.n36712 vdd.n36702 0.01
R64984 vdd.n36756 vdd.n36754 0.01
R64985 vdd.n36943 vdd.n36933 0.01
R64986 vdd.n38042 vdd.n38040 0.01
R64987 vdd.n37998 vdd.n37988 0.01
R64988 vdd.n37811 vdd.n37809 0.01
R64989 vdd.n37767 vdd.n37757 0.01
R64990 vdd.n28209 vdd.n28199 0.01
R64991 vdd.n28253 vdd.n28251 0.01
R64992 vdd.n28440 vdd.n28430 0.01
R64993 vdd.n28484 vdd.n28482 0.01
R64994 vdd.n28671 vdd.n28661 0.01
R64995 vdd.n28715 vdd.n28713 0.01
R64996 vdd.n1673 vdd.n1671 0.01
R64997 vdd.n1639 vdd.n1632 0.01
R64998 vdd.n1492 vdd.n1490 0.01
R64999 vdd.n1458 vdd.n1451 0.01
R65000 vdd.n1311 vdd.n1309 0.01
R65001 vdd.n26777 vdd.n26775 0.01
R65002 vdd.n26924 vdd.n26917 0.01
R65003 vdd.n26958 vdd.n26956 0.01
R65004 vdd.n27105 vdd.n27098 0.01
R65005 vdd.n27139 vdd.n27137 0.01
R65006 vdd.n31162 vdd.n31161 0.01
R65007 vdd.n31180 vdd.n31167 0.01
R65008 vdd.n28858 vdd.n28853 0.01
R65009 vdd.n28924 vdd.n28919 0.01
R65010 vdd.n28035 vdd.n28032 0.01
R65011 vdd.n28032 vdd.n28031 0.01
R65012 vdd.n27948 vdd.n27947 0.01
R65013 vdd.n29786 vdd.n29785 0.01
R65014 vdd.n30635 vdd.n30634 0.01
R65015 vdd.n27597 vdd.n27594 0.01
R65016 vdd.n27465 vdd.n27464 0.01
R65017 vdd.n26013 vdd.n26010 0.01
R65018 vdd.n25911 vdd.n25910 0.01
R65019 vdd.n25614 vdd.n25612 0.01
R65020 vdd.n25558 vdd.n25557 0.01
R65021 vdd.n25446 vdd.n25442 0.01
R65022 vdd.n25669 vdd.n25668 0.01
R65023 vdd.n30958 vdd.n30957 0.01
R65024 vdd.n30791 vdd.n30790 0.01
R65025 vdd.n30989 vdd.n30987 0.01
R65026 vdd.n31213 vdd.n31203 0.01
R65027 vdd.n31213 vdd.n31204 0.01
R65028 vdd.n30800 vdd.n30799 0.01
R65029 vdd.n25372 vdd.n25370 0.01
R65030 vdd.n30773 vdd.n30772 0.01
R65031 vdd.n26126 vdd.n26121 0.01
R65032 vdd.n26129 vdd.n26128 0.01
R65033 vdd.n27693 vdd.n27692 0.01
R65034 vdd.n27715 vdd.n27710 0.01
R65035 vdd.n7204 vdd.n7203 0.01
R65036 vdd.n29621 vdd.n29616 0.01
R65037 vdd.n30927 vdd.n30921 0.01
R65038 vdd.n3672 vdd.n3671 0.01
R65039 vdd.n3873 vdd.n3866 0.01
R65040 vdd.n1882 vdd.n1881 0.01
R65041 vdd.n1836 vdd.n1250 0.01
R65042 vdd.n1288 vdd.n1286 0.01
R65043 vdd.n27229 vdd.n27226 0.01
R65044 vdd.n32110 vdd.n31582 0.01
R65045 vdd.n26160 vdd.n26159 0.01
R65046 vdd.n10249 vdd.n10248 0.01
R65047 vdd.n10262 vdd.n10125 0.01
R65048 vdd.n12600 vdd.n10069 0.01
R65049 vdd.n10560 vdd.n10559 0.01
R65050 vdd.n10630 vdd.n10628 0.01
R65051 vdd.n10705 vdd.n10702 0.01
R65052 vdd.n12348 vdd.n10804 0.01
R65053 vdd.n12311 vdd.n12310 0.01
R65054 vdd.n12259 vdd.n12258 0.01
R65055 vdd.n11071 vdd.n11070 0.01
R65056 vdd.n11163 vdd.n11162 0.01
R65057 vdd.n12098 vdd.n12097 0.01
R65058 vdd.n12042 vdd.n11313 0.01
R65059 vdd.n12005 vdd.n12004 0.01
R65060 vdd.n13940 vdd.n8636 0.01
R65061 vdd.n14016 vdd.n8580 0.01
R65062 vdd.n14230 vdd.n8414 0.01
R65063 vdd.n14313 vdd.n8361 0.01
R65064 vdd.n14555 vdd.n14554 0.01
R65065 vdd.n11607 vdd.n11606 0.01
R65066 vdd.n11614 vdd.n11611 0.01
R65067 vdd.n9081 vdd.n9076 0.01
R65068 vdd.n13449 vdd.n9013 0.01
R65069 vdd.n8861 vdd.n8856 0.01
R65070 vdd.n13740 vdd.n8793 0.01
R65071 vdd.n11500 vdd.n11463 0.01
R65072 vdd.n11501 vdd.n11500 0.01
R65073 vdd.n11589 vdd.n11557 0.01
R65074 vdd.n12579 vdd.n10254 0.01
R65075 vdd.n10331 vdd.n10323 0.01
R65076 vdd.n10363 vdd.n10362 0.01
R65077 vdd.n13008 vdd.n13007 0.01
R65078 vdd.n12968 vdd.n12967 0.01
R65079 vdd.n9589 vdd.n9588 0.01
R65080 vdd.n9655 vdd.n9654 0.01
R65081 vdd.n12800 vdd.n12799 0.01
R65082 vdd.n12760 vdd.n12759 0.01
R65083 vdd.n9949 vdd.n9948 0.01
R65084 vdd.n10015 vdd.n10014 0.01
R65085 vdd.n10161 vdd.n10160 0.01
R65086 vdd.n10166 vdd.n10147 0.01
R65087 vdd.n11905 vdd.n11904 0.01
R65088 vdd.n11827 vdd.n11819 0.01
R65089 vdd.n22229 vdd.n22216 0.01
R65090 vdd.n22105 vdd.n22092 0.01
R65091 vdd.n22295 vdd.n22294 0.01
R65092 vdd.n24353 vdd.n24352 0.01
R65093 vdd.n24267 vdd.n24266 0.01
R65094 vdd.n24252 vdd.n24251 0.01
R65095 vdd.n24236 vdd.n24235 0.01
R65096 vdd.n24160 vdd.n24150 0.01
R65097 vdd.n24024 vdd.n24022 0.01
R65098 vdd.n23928 vdd.n23918 0.01
R65099 vdd.n23792 vdd.n23790 0.01
R65100 vdd.n23696 vdd.n23686 0.01
R65101 vdd.n23104 vdd.n23102 0.01
R65102 vdd.n23240 vdd.n23230 0.01
R65103 vdd.n23336 vdd.n23334 0.01
R65104 vdd.n23472 vdd.n23462 0.01
R65105 vdd.n23568 vdd.n23566 0.01
R65106 vdd.n22525 vdd.n22523 0.01
R65107 vdd.n22661 vdd.n22651 0.01
R65108 vdd.n22757 vdd.n22755 0.01
R65109 vdd.n22893 vdd.n22883 0.01
R65110 vdd.n22989 vdd.n22987 0.01
R65111 vdd.n22439 vdd.n22438 0.01
R65112 vdd.n22424 vdd.n22423 0.01
R65113 vdd.n22408 vdd.n22407 0.01
R65114 vdd.n16604 vdd.n16601 0.01
R65115 vdd.n15059 vdd.n15058 0.01
R65116 vdd.n16743 vdd.n16584 0.01
R65117 vdd.n16920 vdd.n16919 0.01
R65118 vdd.n17060 vdd.n17046 0.01
R65119 vdd.n17192 vdd.n17191 0.01
R65120 vdd.n17332 vdd.n17318 0.01
R65121 vdd.n17464 vdd.n17463 0.01
R65122 vdd.n17592 vdd.n17590 0.01
R65123 vdd.n17722 vdd.n17721 0.01
R65124 vdd.n17862 vdd.n17848 0.01
R65125 vdd.n17993 vdd.n17992 0.01
R65126 vdd.n18133 vdd.n18119 0.01
R65127 vdd.n18262 vdd.n18261 0.01
R65128 vdd.n19067 vdd.n19055 0.01
R65129 vdd.n18988 vdd.n18986 0.01
R65130 vdd.n18808 vdd.n18796 0.01
R65131 vdd.n18729 vdd.n18727 0.01
R65132 vdd.n18549 vdd.n18537 0.01
R65133 vdd.n21645 vdd.n21644 0.01
R65134 vdd.n21653 vdd.n21652 0.01
R65135 vdd.n21433 vdd.n21421 0.01
R65136 vdd.n21354 vdd.n21352 0.01
R65137 vdd.n21174 vdd.n21162 0.01
R65138 vdd.n21095 vdd.n21093 0.01
R65139 vdd.n16803 vdd.n16802 0.01
R65140 vdd.n16802 vdd.n16801 0.01
R65141 vdd.n18428 vdd.n18427 0.01
R65142 vdd.n16792 vdd.n16791 0.01
R65143 vdd.n15399 vdd.n15387 0.01
R65144 vdd.n15447 vdd.n15446 0.01
R65145 vdd.n15647 vdd.n15632 0.01
R65146 vdd.n15703 vdd.n15702 0.01
R65147 vdd.n15903 vdd.n15888 0.01
R65148 vdd.n15959 vdd.n15958 0.01
R65149 vdd.n16159 vdd.n16144 0.01
R65150 vdd.n16215 vdd.n16214 0.01
R65151 vdd.n16415 vdd.n16400 0.01
R65152 vdd.n16471 vdd.n16470 0.01
R65153 vdd.n16575 vdd.n16574 0.01
R65154 vdd.n16582 vdd.n16577 0.01
R65155 vdd.n21996 vdd.n21995 0.01
R65156 vdd.n21918 vdd.n21910 0.01
R65157 vdd.n24551 vdd.n24550 0.01
R65158 vdd.n24907 vdd.n24904 0.01
R65159 vdd.n25037 vdd.n25035 0.01
R65160 vdd.n25015 vdd.n25012 0.01
R65161 vdd.n24916 vdd.n24913 0.01
R65162 vdd.n24612 vdd.n24610 0.01
R65163 vdd.n24591 vdd.n24588 0.01
R65164 vdd.n24627 vdd.n24624 0.01
R65165 vdd.n25252 vdd.n25251 0.01
R65166 vdd.n11889 vdd.n11800 0.01
R65167 vdd.n21980 vdd.n21891 0.01
R65168 vdd.n35425 vdd.n35424 0.01
R65169 vdd.n6213 vdd.n6212 0.01
R65170 vdd.n30808 vdd.n30807 0.01
R65171 vdd.n5008 vdd.n5007 0.01
R65172 vdd.n4402 vdd.n4401 0.01
R65173 vdd.n31319 vdd.n31310 0.01
R65174 vdd.n34406 vdd.n34405 0.01
R65175 vdd.n34829 vdd.n34828 0.01
R65176 vdd.n5576 vdd.n5575 0.01
R65177 vdd.n1172 vdd.n1171 0.01
R65178 vdd.n29973 vdd.n29968 0.01
R65179 vdd.n31697 vdd.n31696 0.01
R65180 vdd.n210 vdd.n209 0.01
R65181 vdd.n30083 vdd.n30082 0.01
R65182 vdd.n29290 vdd.n29289 0.01
R65183 vdd.n26661 vdd.n26660 0.01
R65184 vdd.n4951 vdd.n4950 0.01
R65185 vdd.n31372 vdd.n31371 0.01
R65186 vdd.n31215 vdd.n31214 0.01
R65187 vdd.n12576 vdd.n10257 0.01
R65188 vdd.n15120 vdd.n15045 0.01
R65189 vdd.n33571 vdd.n33570 0.009
R65190 vdd.n11723 vdd.n11722 0.009
R65191 vdd.n21804 vdd.n21803 0.009
R65192 vdd.n27208 vdd.n26757 0.009
R65193 vdd.n25627 vdd.n25625 0.009
R65194 vdd.n25549 vdd.n25547 0.009
R65195 vdd.n25463 vdd.n25461 0.009
R65196 vdd.n32133 vdd.n31577 0.009
R65197 vdd.n2387 vdd.n2372 0.009
R65198 vdd.n1912 vdd.n1210 0.009
R65199 vdd.n26125 vdd.n26123 0.009
R65200 vdd.n305 vdd.n304 0.009
R65201 vdd.n29519 vdd.n29518 0.009
R65202 vdd.n30785 vdd.n30784 0.009
R65203 vdd.n33365 vdd.n33364 0.009
R65204 vdd.n33315 vdd.n33314 0.009
R65205 vdd.n33696 vdd.n33695 0.009
R65206 vdd.n33617 vdd.n33616 0.009
R65207 vdd.n33788 vdd.n33787 0.009
R65208 vdd.n35491 vdd.n35478 0.009
R65209 vdd.n35114 vdd.n35100 0.009
R65210 vdd.n35427 vdd.n35426 0.009
R65211 vdd.n35449 vdd.n35448 0.009
R65212 vdd.n35181 vdd.n35180 0.009
R65213 vdd.n35211 vdd.n35210 0.009
R65214 vdd.n35316 vdd.n35315 0.009
R65215 vdd.n575 vdd.n574 0.009
R65216 vdd.n192 vdd.n191 0.009
R65217 vdd.n215 vdd.n214 0.009
R65218 vdd.n5827 vdd.n5826 0.009
R65219 vdd.n6247 vdd.n6246 0.009
R65220 vdd.n6211 vdd.n6210 0.009
R65221 vdd.n6123 vdd.n6122 0.009
R65222 vdd.n6317 vdd.n6316 0.009
R65223 vdd.n6334 vdd.n6333 0.009
R65224 vdd.n5872 vdd.n5871 0.009
R65225 vdd.n4942 vdd.n4941 0.009
R65226 vdd.n4543 vdd.n4542 0.009
R65227 vdd.n4314 vdd.n4313 0.009
R65228 vdd.n4104 vdd.n4090 0.009
R65229 vdd.n4404 vdd.n4403 0.009
R65230 vdd.n4426 vdd.n4425 0.009
R65231 vdd.n4184 vdd.n4183 0.009
R65232 vdd.n4201 vdd.n4200 0.009
R65233 vdd.n30208 vdd.n30207 0.009
R65234 vdd.n29951 vdd.n29950 0.009
R65235 vdd.n27818 vdd.n27817 0.009
R65236 vdd.n30621 vdd.n30254 0.009
R65237 vdd.n30603 vdd.n30277 0.009
R65238 vdd.n28892 vdd.n28888 0.009
R65239 vdd.n28905 vdd.n28903 0.009
R65240 vdd.n28919 vdd.n28916 0.009
R65241 vdd.n28926 vdd.n28925 0.009
R65242 vdd.n28044 vdd.n28041 0.009
R65243 vdd.n27968 vdd.n27966 0.009
R65244 vdd.n27959 vdd.n27957 0.009
R65245 vdd.n27944 vdd.n27943 0.009
R65246 vdd.n29799 vdd.n29798 0.009
R65247 vdd.n30690 vdd.n30676 0.009
R65248 vdd.n25609 vdd.n25607 0.009
R65249 vdd.n31316 vdd.n31315 0.009
R65250 vdd.n25368 vdd.n25367 0.009
R65251 vdd.n30798 vdd.n30797 0.009
R65252 vdd.n26083 vdd.n25376 0.009
R65253 vdd.n26320 vdd.n26278 0.009
R65254 vdd.n29432 vdd.n29424 0.009
R65255 vdd.n7201 vdd.n7200 0.009
R65256 vdd.n31428 vdd.n31420 0.009
R65257 vdd.n30831 vdd.n30821 0.009
R65258 vdd.n30784 vdd.n30783 0.009
R65259 vdd.n26549 vdd.n26542 0.009
R65260 vdd.n29481 vdd.n29475 0.009
R65261 vdd.n30164 vdd.n30159 0.009
R65262 vdd.n7211 vdd.n7210 0.009
R65263 vdd.n2219 vdd.n2211 0.009
R65264 vdd.n2257 vdd.n2170 0.009
R65265 vdd.n2294 vdd.n2132 0.009
R65266 vdd.n2341 vdd.n2108 0.009
R65267 vdd.n2554 vdd.n2410 0.009
R65268 vdd.n1892 vdd.n1890 0.009
R65269 vdd.n1915 vdd.n1914 0.009
R65270 vdd.n26214 vdd.n26213 0.009
R65271 vdd.n26669 vdd.n26668 0.009
R65272 vdd.n31936 vdd.n31935 0.009
R65273 vdd.n32454 vdd.n32453 0.009
R65274 vdd.n10268 vdd.n10267 0.009
R65275 vdd.n12573 vdd.n10268 0.009
R65276 vdd.n11534 vdd.n11453 0.009
R65277 vdd.n11555 vdd.n11544 0.009
R65278 vdd.n11941 vdd.n11940 0.009
R65279 vdd.n11590 vdd.n11554 0.009
R65280 vdd.n13884 vdd.n8651 0.009
R65281 vdd.n14085 vdd.n14084 0.009
R65282 vdd.n14173 vdd.n8431 0.009
R65283 vdd.n8328 vdd.n8324 0.009
R65284 vdd.n14474 vdd.n14473 0.009
R65285 vdd.n13798 vdd.n13797 0.009
R65286 vdd.n11607 vdd.n11580 0.009
R65287 vdd.n11622 vdd.n11583 0.009
R65288 vdd.n13173 vdd.n13172 0.009
R65289 vdd.n13311 vdd.n13310 0.009
R65290 vdd.n13468 vdd.n13463 0.009
R65291 vdd.n13603 vdd.n13602 0.009
R65292 vdd.n11609 vdd.n11608 0.009
R65293 vdd.n11621 vdd.n11620 0.009
R65294 vdd.n10215 vdd.n10211 0.009
R65295 vdd.n10283 vdd.n10274 0.009
R65296 vdd.n10424 vdd.n10423 0.009
R65297 vdd.n13055 vdd.n9305 0.009
R65298 vdd.n9378 vdd.n9365 0.009
R65299 vdd.n9504 vdd.n9480 0.009
R65300 vdd.n9551 vdd.n9548 0.009
R65301 vdd.n12847 vdd.n9665 0.009
R65302 vdd.n9738 vdd.n9725 0.009
R65303 vdd.n9864 vdd.n9840 0.009
R65304 vdd.n9911 vdd.n9908 0.009
R65305 vdd.n12639 vdd.n10025 0.009
R65306 vdd.n11748 vdd.n11719 0.009
R65307 vdd.n11878 vdd.n11801 0.009
R65308 vdd.n13690 vdd.n13689 0.009
R65309 vdd.n8671 vdd.n8670 0.009
R65310 vdd.n22343 vdd.n22229 0.009
R65311 vdd.n22240 vdd.n22239 0.009
R65312 vdd.n24306 vdd.n22105 0.009
R65313 vdd.n22115 vdd.n22107 0.009
R65314 vdd.n22311 vdd.n22309 0.009
R65315 vdd.n24338 vdd.n24337 0.009
R65316 vdd.n24283 vdd.n24281 0.009
R65317 vdd.n24221 vdd.n24220 0.009
R65318 vdd.n22455 vdd.n22453 0.009
R65319 vdd.n22393 vdd.n22392 0.009
R65320 vdd.n15042 vdd.n15041 0.009
R65321 vdd.n15043 vdd.n15042 0.009
R65322 vdd.n18373 vdd.n18372 0.009
R65323 vdd.n18390 vdd.n18389 0.009
R65324 vdd.n18393 vdd.n18392 0.009
R65325 vdd.n18405 vdd.n18404 0.009
R65326 vdd.n19103 vdd.n19101 0.009
R65327 vdd.n18942 vdd.n18940 0.009
R65328 vdd.n18844 vdd.n18842 0.009
R65329 vdd.n18683 vdd.n18681 0.009
R65330 vdd.n18585 vdd.n18583 0.009
R65331 vdd.n21049 vdd.n21047 0.009
R65332 vdd.n21646 vdd.n21645 0.009
R65333 vdd.n21649 vdd.n21648 0.009
R65334 vdd.n21567 vdd.n21565 0.009
R65335 vdd.n21469 vdd.n21467 0.009
R65336 vdd.n21308 vdd.n21306 0.009
R65337 vdd.n21210 vdd.n21208 0.009
R65338 vdd.n21696 vdd.n21695 0.009
R65339 vdd.n21694 vdd.n21693 0.009
R65340 vdd.n16785 vdd.n16784 0.009
R65341 vdd.n15278 vdd.n15266 0.009
R65342 vdd.n15358 vdd.n15357 0.009
R65343 vdd.n15500 vdd.n15485 0.009
R65344 vdd.n15597 vdd.n15596 0.009
R65345 vdd.n15756 vdd.n15741 0.009
R65346 vdd.n15853 vdd.n15852 0.009
R65347 vdd.n16012 vdd.n15997 0.009
R65348 vdd.n16109 vdd.n16108 0.009
R65349 vdd.n16268 vdd.n16253 0.009
R65350 vdd.n16365 vdd.n16364 0.009
R65351 vdd.n16524 vdd.n16509 0.009
R65352 vdd.n19732 vdd.n19731 0.009
R65353 vdd.n20929 vdd.n20928 0.009
R65354 vdd.n21831 vdd.n21830 0.009
R65355 vdd.n21969 vdd.n21892 0.009
R65356 vdd.n24554 vdd.n24553 0.009
R65357 vdd.n24951 vdd.n24950 0.009
R65358 vdd.n25253 vdd.n25252 0.009
R65359 vdd.n11745 vdd.n11744 0.009
R65360 vdd.n21827 vdd.n21826 0.009
R65361 vdd.n25641 vdd.n25640 0.009
R65362 vdd.n31213 vdd.n31212 0.009
R65363 vdd.n4807 vdd.n4806 0.009
R65364 vdd.n32014 vdd.n32013 0.009
R65365 vdd.n32357 vdd.n32356 0.009
R65366 vdd.n1837 vdd.n1836 0.009
R65367 vdd.n32002 vdd.n31996 0.009
R65368 vdd.n32329 vdd.n32323 0.009
R65369 vdd.n32346 vdd.n32340 0.009
R65370 vdd.n30820 vdd.n30819 0.009
R65371 vdd.n11891 vdd.n11890 0.009
R65372 vdd.n21982 vdd.n21981 0.009
R65373 vdd.n1826 vdd.n1820 0.009
R65374 vdd.n24548 vdd.n24544 0.009
R65375 vdd.n26162 vdd.n26161 0.008
R65376 vdd.n31386 vdd.n31384 0.008
R65377 vdd.n30998 vdd.n30990 0.008
R65378 vdd.n26486 vdd.n26485 0.008
R65379 vdd.n30900 vdd.n30899 0.008
R65380 vdd.n234 vdd.n233 0.008
R65381 vdd.n30755 vdd.n30754 0.008
R65382 vdd.n7161 vdd.n7160 0.008
R65383 vdd.n33452 vdd.n33451 0.008
R65384 vdd.n466 vdd.n465 0.008
R65385 vdd.n184 vdd.n183 0.008
R65386 vdd.n380 vdd.n377 0.008
R65387 vdd.n2249 vdd.n2248 0.008
R65388 vdd.n5186 vdd.n5067 0.008
R65389 vdd.n29185 vdd.n29183 0.008
R65390 vdd.n30816 vdd.n30814 0.008
R65391 vdd.n26215 vdd.n26182 0.008
R65392 vdd.n2787 vdd.n2785 0.008
R65393 vdd.n2815 vdd.n2813 0.008
R65394 vdd.n2968 vdd.n2966 0.008
R65395 vdd.n2996 vdd.n2994 0.008
R65396 vdd.n3149 vdd.n3147 0.008
R65397 vdd.n3177 vdd.n3175 0.008
R65398 vdd.n3330 vdd.n3328 0.008
R65399 vdd.n3358 vdd.n3356 0.008
R65400 vdd.n3511 vdd.n3509 0.008
R65401 vdd.n3539 vdd.n3537 0.008
R65402 vdd.n1770 vdd.n1763 0.008
R65403 vdd.n1752 vdd.n1750 0.008
R65404 vdd.n33692 vdd.n33691 0.008
R65405 vdd.n33648 vdd.n33647 0.008
R65406 vdd.n34231 vdd.n34230 0.008
R65407 vdd.n34227 vdd.n34226 0.008
R65408 vdd.n34057 vdd.n34056 0.008
R65409 vdd.n35055 vdd.n35054 0.008
R65410 vdd.n35233 vdd.n35129 0.008
R65411 vdd.n35218 vdd.n35217 0.008
R65412 vdd.n35192 vdd.n35191 0.008
R65413 vdd.n35348 vdd.n35347 0.008
R65414 vdd.n34764 vdd.n34763 0.008
R65415 vdd.n34631 vdd.n34630 0.008
R65416 vdd.n1158 vdd.n1157 0.008
R65417 vdd.n869 vdd.n868 0.008
R65418 vdd.n312 vdd.n311 0.008
R65419 vdd.n6195 vdd.n6194 0.008
R65420 vdd.n6356 vdd.n6258 0.008
R65421 vdd.n6342 vdd.n6341 0.008
R65422 vdd.n6355 vdd.n6354 0.008
R65423 vdd.n6298 vdd.n6297 0.008
R65424 vdd.n5854 vdd.n5853 0.008
R65425 vdd.n5511 vdd.n5510 0.008
R65426 vdd.n5378 vdd.n5377 0.008
R65427 vdd.n5172 vdd.n5171 0.008
R65428 vdd.n4338 vdd.n4337 0.008
R65429 vdd.n4045 vdd.n4044 0.008
R65430 vdd.n4208 vdd.n4207 0.008
R65431 vdd.n4165 vdd.n4164 0.008
R65432 vdd.n38143 vdd.n38141 0.008
R65433 vdd.n35904 vdd.n35902 0.008
R65434 vdd.n35939 vdd.n35937 0.008
R65435 vdd.n36135 vdd.n36133 0.008
R65436 vdd.n36170 vdd.n36168 0.008
R65437 vdd.n36366 vdd.n36364 0.008
R65438 vdd.n36401 vdd.n36399 0.008
R65439 vdd.n36597 vdd.n36595 0.008
R65440 vdd.n36632 vdd.n36630 0.008
R65441 vdd.n36828 vdd.n36826 0.008
R65442 vdd.n36863 vdd.n36861 0.008
R65443 vdd.n38114 vdd.n38112 0.008
R65444 vdd.n37918 vdd.n37916 0.008
R65445 vdd.n37883 vdd.n37881 0.008
R65446 vdd.n37687 vdd.n37685 0.008
R65447 vdd.n37652 vdd.n37650 0.008
R65448 vdd.n28325 vdd.n28323 0.008
R65449 vdd.n28360 vdd.n28358 0.008
R65450 vdd.n28556 vdd.n28554 0.008
R65451 vdd.n28591 vdd.n28589 0.008
R65452 vdd.n28787 vdd.n28785 0.008
R65453 vdd.n1730 vdd.n1728 0.008
R65454 vdd.n1577 vdd.n1575 0.008
R65455 vdd.n1549 vdd.n1547 0.008
R65456 vdd.n1396 vdd.n1394 0.008
R65457 vdd.n1368 vdd.n1366 0.008
R65458 vdd.n26834 vdd.n26832 0.008
R65459 vdd.n26862 vdd.n26860 0.008
R65460 vdd.n27015 vdd.n27013 0.008
R65461 vdd.n27043 vdd.n27041 0.008
R65462 vdd.n27196 vdd.n27194 0.008
R65463 vdd.n29824 vdd.n29823 0.008
R65464 vdd.n27943 vdd.n27942 0.008
R65465 vdd.n28934 vdd.n28074 0.008
R65466 vdd.n28877 vdd.n28876 0.008
R65467 vdd.n29017 vdd.n29016 0.008
R65468 vdd.n27990 vdd.n27988 0.008
R65469 vdd.n27951 vdd.n27949 0.008
R65470 vdd.n30665 vdd.n30664 0.008
R65471 vdd.n30638 vdd.n30636 0.008
R65472 vdd.n30531 vdd.n30524 0.008
R65473 vdd.n30517 vdd.n30510 0.008
R65474 vdd.n27603 vdd.n27601 0.008
R65475 vdd.n27354 vdd.n27353 0.008
R65476 vdd.n26019 vdd.n26017 0.008
R65477 vdd.n25806 vdd.n25805 0.008
R65478 vdd.n25525 vdd.n25523 0.008
R65479 vdd.n25489 vdd.n25488 0.008
R65480 vdd.n30903 vdd.n30902 0.008
R65481 vdd.n32577 vdd.n32576 0.008
R65482 vdd.n29599 vdd.n29598 0.008
R65483 vdd.n29394 vdd.n29393 0.008
R65484 vdd.n27693 vdd.n27691 0.008
R65485 vdd.n26254 vdd.n26253 0.008
R65486 vdd.n30968 vdd.n30967 0.008
R65487 vdd.n30954 vdd.n30949 0.008
R65488 vdd.n26160 vdd.n26158 0.008
R65489 vdd.n30811 vdd.n30810 0.008
R65490 vdd.n7196 vdd.n7195 0.008
R65491 vdd.n26520 vdd.n26513 0.008
R65492 vdd.n29093 vdd.n29087 0.008
R65493 vdd.n32664 vdd.n32655 0.008
R65494 vdd.n30767 vdd.n30745 0.008
R65495 vdd.n27671 vdd.n27670 0.008
R65496 vdd.n27695 vdd.n27688 0.008
R65497 vdd.n29576 vdd.n29575 0.008
R65498 vdd.n29601 vdd.n29595 0.008
R65499 vdd.n30025 vdd.n30024 0.008
R65500 vdd.n30881 vdd.n30880 0.008
R65501 vdd.n30905 vdd.n30898 0.008
R65502 vdd.n7207 vdd.n7206 0.008
R65503 vdd.n7223 vdd.n7222 0.008
R65504 vdd.n29566 vdd.n29565 0.008
R65505 vdd.n3717 vdd.n3712 0.008
R65506 vdd.n3938 vdd.n3932 0.008
R65507 vdd.n3921 vdd.n3916 0.008
R65508 vdd.n2290 vdd.n2285 0.008
R65509 vdd.n2557 vdd.n2556 0.008
R65510 vdd.n1967 vdd.n1962 0.008
R65511 vdd.n2000 vdd.n1998 0.008
R65512 vdd.n1836 vdd.n1831 0.008
R65513 vdd.n31684 vdd.n31679 0.008
R65514 vdd.n27242 vdd.n27241 0.008
R65515 vdd.n31788 vdd.n31730 0.008
R65516 vdd.n26317 vdd.n26316 0.008
R65517 vdd.n31788 vdd.n31787 0.008
R65518 vdd.n31881 vdd.n31880 0.008
R65519 vdd.n31906 vdd.n31905 0.008
R65520 vdd.n32110 vdd.n32109 0.008
R65521 vdd.n32254 vdd.n32253 0.008
R65522 vdd.n32487 vdd.n32486 0.008
R65523 vdd.n31184 vdd.n31181 0.008
R65524 vdd.n31302 vdd.n31296 0.008
R65525 vdd.n10200 vdd.n10199 0.008
R65526 vdd.n10233 vdd.n10232 0.008
R65527 vdd.n10226 vdd.n10225 0.008
R65528 vdd.n10559 vdd.n10534 0.008
R65529 vdd.n10652 vdd.n10628 0.008
R65530 vdd.n12406 vdd.n10702 0.008
R65531 vdd.n12348 vdd.n12347 0.008
R65532 vdd.n12312 vdd.n12311 0.008
R65533 vdd.n12258 vdd.n12257 0.008
R65534 vdd.n11070 vdd.n11069 0.008
R65535 vdd.n11164 vdd.n11163 0.008
R65536 vdd.n12098 vdd.n11218 0.008
R65537 vdd.n12042 vdd.n12041 0.008
R65538 vdd.n12006 vdd.n12005 0.008
R65539 vdd.n11509 vdd.n11508 0.008
R65540 vdd.n13922 vdd.n13921 0.008
R65541 vdd.n8652 vdd.n8638 0.008
R65542 vdd.n14035 vdd.n14028 0.008
R65543 vdd.n14034 vdd.n14029 0.008
R65544 vdd.n14212 vdd.n14211 0.008
R65545 vdd.n8432 vdd.n8416 0.008
R65546 vdd.n14314 vdd.n8323 0.008
R65547 vdd.n14367 vdd.n14366 0.008
R65548 vdd.n14477 vdd.n14476 0.008
R65549 vdd.n8195 vdd.n8193 0.008
R65550 vdd.n13749 vdd.n8789 0.008
R65551 vdd.n13165 vdd.n9231 0.008
R65552 vdd.n13166 vdd.n9229 0.008
R65553 vdd.n9115 vdd.n9114 0.008
R65554 vdd.n9118 vdd.n9117 0.008
R65555 vdd.n13450 vdd.n9008 0.008
R65556 vdd.n13462 vdd.n13461 0.008
R65557 vdd.n8894 vdd.n8893 0.008
R65558 vdd.n8897 vdd.n8896 0.008
R65559 vdd.n11556 vdd.n11542 0.008
R65560 vdd.n10313 vdd.n10310 0.008
R65561 vdd.n10411 vdd.n10410 0.008
R65562 vdd.n9304 vdd.n9302 0.008
R65563 vdd.n13067 vdd.n13066 0.008
R65564 vdd.n13020 vdd.n9392 0.008
R65565 vdd.n13019 vdd.n9393 0.008
R65566 vdd.n9489 vdd.n9458 0.008
R65567 vdd.n9493 vdd.n9492 0.008
R65568 vdd.n12912 vdd.n12911 0.008
R65569 vdd.n9583 vdd.n9559 0.008
R65570 vdd.n9664 vdd.n9662 0.008
R65571 vdd.n12859 vdd.n12858 0.008
R65572 vdd.n12812 vdd.n9752 0.008
R65573 vdd.n12811 vdd.n9753 0.008
R65574 vdd.n9849 vdd.n9818 0.008
R65575 vdd.n9853 vdd.n9852 0.008
R65576 vdd.n12704 vdd.n12703 0.008
R65577 vdd.n9943 vdd.n9918 0.008
R65578 vdd.n10024 vdd.n10022 0.008
R65579 vdd.n12651 vdd.n12650 0.008
R65580 vdd.n10168 vdd.n10145 0.008
R65581 vdd.n10173 vdd.n10172 0.008
R65582 vdd.n12622 vdd.n12621 0.008
R65583 vdd.n11894 vdd.n11796 0.008
R65584 vdd.n22213 vdd.n22203 0.008
R65585 vdd.n22078 vdd.n22077 0.008
R65586 vdd.n22340 vdd.n22330 0.008
R65587 vdd.n22330 vdd.n22329 0.008
R65588 vdd.n22325 vdd.n22324 0.008
R65589 vdd.n24368 vdd.n24367 0.008
R65590 vdd.n24323 vdd.n24322 0.008
R65591 vdd.n24303 vdd.n24302 0.008
R65592 vdd.n24302 vdd.n24301 0.008
R65593 vdd.n24297 vdd.n24296 0.008
R65594 vdd.n24206 vdd.n24205 0.008
R65595 vdd.n24122 vdd.n24120 0.008
R65596 vdd.n24054 vdd.n24052 0.008
R65597 vdd.n23890 vdd.n23888 0.008
R65598 vdd.n23822 vdd.n23820 0.008
R65599 vdd.n23658 vdd.n23656 0.008
R65600 vdd.n23134 vdd.n23132 0.008
R65601 vdd.n23202 vdd.n23200 0.008
R65602 vdd.n23366 vdd.n23364 0.008
R65603 vdd.n23434 vdd.n23432 0.008
R65604 vdd.n23598 vdd.n23596 0.008
R65605 vdd.n22555 vdd.n22553 0.008
R65606 vdd.n22623 vdd.n22621 0.008
R65607 vdd.n22787 vdd.n22785 0.008
R65608 vdd.n22855 vdd.n22853 0.008
R65609 vdd.n23019 vdd.n23017 0.008
R65610 vdd.n22469 vdd.n22468 0.008
R65611 vdd.n22378 vdd.n22377 0.008
R65612 vdd.n16693 vdd.n16692 0.008
R65613 vdd.n16587 vdd.n16585 0.008
R65614 vdd.n16677 vdd.n16676 0.008
R65615 vdd.n16919 vdd.n16905 0.008
R65616 vdd.n17061 vdd.n17060 0.008
R65617 vdd.n17191 vdd.n17177 0.008
R65618 vdd.n17333 vdd.n17332 0.008
R65619 vdd.n17463 vdd.n17449 0.008
R65620 vdd.n17592 vdd.n17591 0.008
R65621 vdd.n17721 vdd.n17707 0.008
R65622 vdd.n17863 vdd.n17862 0.008
R65623 vdd.n17992 vdd.n17978 0.008
R65624 vdd.n18134 vdd.n18133 0.008
R65625 vdd.n18261 vdd.n18248 0.008
R65626 vdd.n18335 vdd.n18334 0.008
R65627 vdd.n19087 vdd.n19085 0.008
R65628 vdd.n19083 vdd.n19071 0.008
R65629 vdd.n18972 vdd.n18970 0.008
R65630 vdd.n18958 vdd.n18956 0.008
R65631 vdd.n18828 vdd.n18826 0.008
R65632 vdd.n18824 vdd.n18812 0.008
R65633 vdd.n18713 vdd.n18711 0.008
R65634 vdd.n18699 vdd.n18697 0.008
R65635 vdd.n18569 vdd.n18567 0.008
R65636 vdd.n18565 vdd.n18553 0.008
R65637 vdd.n21079 vdd.n21077 0.008
R65638 vdd.n21597 vdd.n21595 0.008
R65639 vdd.n21583 vdd.n21581 0.008
R65640 vdd.n21453 vdd.n21451 0.008
R65641 vdd.n21449 vdd.n21437 0.008
R65642 vdd.n21338 vdd.n21336 0.008
R65643 vdd.n21324 vdd.n21322 0.008
R65644 vdd.n21194 vdd.n21192 0.008
R65645 vdd.n21190 vdd.n21178 0.008
R65646 vdd.n18426 vdd.n18425 0.008
R65647 vdd.n15372 vdd.n15371 0.008
R65648 vdd.n15385 vdd.n15373 0.008
R65649 vdd.n15467 vdd.n15466 0.008
R65650 vdd.n15483 vdd.n15468 0.008
R65651 vdd.n15614 vdd.n15613 0.008
R65652 vdd.n15630 vdd.n15615 0.008
R65653 vdd.n15723 vdd.n15722 0.008
R65654 vdd.n15739 vdd.n15724 0.008
R65655 vdd.n15870 vdd.n15869 0.008
R65656 vdd.n15886 vdd.n15871 0.008
R65657 vdd.n15979 vdd.n15978 0.008
R65658 vdd.n15995 vdd.n15980 0.008
R65659 vdd.n16126 vdd.n16125 0.008
R65660 vdd.n16142 vdd.n16127 0.008
R65661 vdd.n16235 vdd.n16234 0.008
R65662 vdd.n16251 vdd.n16236 0.008
R65663 vdd.n16382 vdd.n16381 0.008
R65664 vdd.n16398 vdd.n16383 0.008
R65665 vdd.n16491 vdd.n16490 0.008
R65666 vdd.n16507 vdd.n16492 0.008
R65667 vdd.n16768 vdd.n16764 0.008
R65668 vdd.n16763 vdd.n16762 0.008
R65669 vdd.n16755 vdd.n16754 0.008
R65670 vdd.n21985 vdd.n21887 0.008
R65671 vdd.n24556 vdd.n24555 0.008
R65672 vdd.n24973 vdd.n24972 0.008
R65673 vdd.n24972 vdd.n24970 0.008
R65674 vdd.n25050 vdd.n25048 0.008
R65675 vdd.n24629 vdd.n24627 0.008
R65676 vdd.n26120 vdd.n26119 0.008
R65677 vdd.n31326 vdd.n31325 0.008
R65678 vdd.n25571 vdd.n25570 0.008
R65679 vdd.n25497 vdd.n25496 0.008
R65680 vdd.n30943 vdd.n30941 0.008
R65681 vdd.n2669 vdd.n2665 0.008
R65682 vdd.n31289 vdd.n31288 0.008
R65683 vdd.n30964 vdd.n30963 0.008
R65684 vdd.n32390 vdd.n32389 0.008
R65685 vdd.n31955 vdd.n31954 0.008
R65686 vdd.n25514 vdd.n25513 0.008
R65687 vdd.n30961 vdd.n30960 0.008
R65688 vdd.n27558 vdd.n27557 0.008
R65689 vdd.n31012 vdd.n31011 0.008
R65690 vdd.n31326 vdd.n31320 0.008
R65691 vdd.n34061 vdd.n34060 0.007
R65692 vdd.n6039 vdd.n6038 0.007
R65693 vdd.n5923 vdd.n5920 0.007
R65694 vdd.n25568 vdd.n25561 0.007
R65695 vdd.n30782 vdd.n30781 0.007
R65696 vdd.n31211 vdd.n31210 0.007
R65697 vdd.n25264 vdd.n7971 0.007
R65698 vdd.n30997 vdd.n30996 0.007
R65699 vdd.n30945 vdd.n30944 0.007
R65700 vdd.n32090 vdd.n32088 0.007
R65701 vdd.n25569 vdd.n25568 0.007
R65702 vdd.n32538 vdd.n32536 0.007
R65703 vdd.n33412 vdd.n33410 0.007
R65704 vdd.n33416 vdd.n33414 0.007
R65705 vdd.n33448 vdd.n33447 0.007
R65706 vdd.n33462 vdd.n33461 0.007
R65707 vdd.n33470 vdd.n33469 0.007
R65708 vdd.n33502 vdd.n33501 0.007
R65709 vdd.n33496 vdd.n33495 0.007
R65710 vdd.n33523 vdd.n33518 0.007
R65711 vdd.n33530 vdd.n33528 0.007
R65712 vdd.n33534 vdd.n33531 0.007
R65713 vdd.n33309 vdd.n33307 0.007
R65714 vdd.n33300 vdd.n33299 0.007
R65715 vdd.n33757 vdd.n33754 0.007
R65716 vdd.n33745 vdd.n33744 0.007
R65717 vdd.n33611 vdd.n33610 0.007
R65718 vdd.n33619 vdd.n33618 0.007
R65719 vdd.n33622 vdd.n33619 0.007
R65720 vdd.n33666 vdd.n33665 0.007
R65721 vdd.n33639 vdd.n33638 0.007
R65722 vdd.n34090 vdd.n34089 0.007
R65723 vdd.n34107 vdd.n34106 0.007
R65724 vdd.n34138 vdd.n34134 0.007
R65725 vdd.n34122 vdd.n34117 0.007
R65726 vdd.n34256 vdd.n34254 0.007
R65727 vdd.n34273 vdd.n34270 0.007
R65728 vdd.n34334 vdd.n34333 0.007
R65729 vdd.n34188 vdd.n34187 0.007
R65730 vdd.n34364 vdd.n34363 0.007
R65731 vdd.n34358 vdd.n34357 0.007
R65732 vdd.n34376 vdd.n34371 0.007
R65733 vdd.n34402 vdd.n34400 0.007
R65734 vdd.n33926 vdd.n33923 0.007
R65735 vdd.n33905 vdd.n33904 0.007
R65736 vdd.n33921 vdd.n33920 0.007
R65737 vdd.n33934 vdd.n33933 0.007
R65738 vdd.n34069 vdd.n34068 0.007
R65739 vdd.n33986 vdd.n33985 0.007
R65740 vdd.n33998 vdd.n33996 0.007
R65741 vdd.n34007 vdd.n34005 0.007
R65742 vdd.n34028 vdd.n34027 0.007
R65743 vdd.n34030 vdd.n34029 0.007
R65744 vdd.n35169 vdd.n35167 0.007
R65745 vdd.n35160 vdd.n35158 0.007
R65746 vdd.n35148 vdd.n35147 0.007
R65747 vdd.n35539 vdd.n35536 0.007
R65748 vdd.n35522 vdd.n35520 0.007
R65749 vdd.n35510 vdd.n35509 0.007
R65750 vdd.n35485 vdd.n35482 0.007
R65751 vdd.n35475 vdd.n35474 0.007
R65752 vdd.n35251 vdd.n35250 0.007
R65753 vdd.n35600 vdd.n35599 0.007
R65754 vdd.n35074 vdd.n35073 0.007
R65755 vdd.n35052 vdd.n35050 0.007
R65756 vdd.n35417 vdd.n35414 0.007
R65757 vdd.n35399 vdd.n35394 0.007
R65758 vdd.n35374 vdd.n35373 0.007
R65759 vdd.n35380 vdd.n35379 0.007
R65760 vdd.n35298 vdd.n35297 0.007
R65761 vdd.n34664 vdd.n34663 0.007
R65762 vdd.n34957 vdd.n34954 0.007
R65763 vdd.n34682 vdd.n34681 0.007
R65764 vdd.n34977 vdd.n34976 0.007
R65765 vdd.n34937 vdd.n34935 0.007
R65766 vdd.n34928 vdd.n34925 0.007
R65767 vdd.n35012 vdd.n35011 0.007
R65768 vdd.n34714 vdd.n34713 0.007
R65769 vdd.n34790 vdd.n34789 0.007
R65770 vdd.n34784 vdd.n34783 0.007
R65771 vdd.n34802 vdd.n34797 0.007
R65772 vdd.n34821 vdd.n34818 0.007
R65773 vdd.n34465 vdd.n34463 0.007
R65774 vdd.n34487 vdd.n34486 0.007
R65775 vdd.n34462 vdd.n34461 0.007
R65776 vdd.n34468 vdd.n34467 0.007
R65777 vdd.n34563 vdd.n34562 0.007
R65778 vdd.n34578 vdd.n34576 0.007
R65779 vdd.n34591 vdd.n34589 0.007
R65780 vdd.n34587 vdd.n34586 0.007
R65781 vdd.n34612 vdd.n34611 0.007
R65782 vdd.n736 vdd.n734 0.007
R65783 vdd.n742 vdd.n740 0.007
R65784 vdd.n767 vdd.n766 0.007
R65785 vdd.n710 vdd.n709 0.007
R65786 vdd.n992 vdd.n991 0.007
R65787 vdd.n986 vdd.n985 0.007
R65788 vdd.n1004 vdd.n999 0.007
R65789 vdd.n1013 vdd.n1011 0.007
R65790 vdd.n647 vdd.n646 0.007
R65791 vdd.n638 vdd.n636 0.007
R65792 vdd.n656 vdd.n655 0.007
R65793 vdd.n896 vdd.n895 0.007
R65794 vdd.n918 vdd.n915 0.007
R65795 vdd.n1104 vdd.n1103 0.007
R65796 vdd.n1095 vdd.n1094 0.007
R65797 vdd.n1098 vdd.n1095 0.007
R65798 vdd.n1059 vdd.n1058 0.007
R65799 vdd.n1076 vdd.n1075 0.007
R65800 vdd.n1133 vdd.n1132 0.007
R65801 vdd.n859 vdd.n858 0.007
R65802 vdd.n536 vdd.n534 0.007
R65803 vdd.n383 vdd.n382 0.007
R65804 vdd.n383 vdd.n381 0.007
R65805 vdd.n484 vdd.n483 0.007
R65806 vdd.n6 vdd.n5 0.007
R65807 vdd.n8 vdd.n7 0.007
R65808 vdd.n397 vdd.n396 0.007
R65809 vdd.n414 vdd.n411 0.007
R65810 vdd.n427 vdd.n425 0.007
R65811 vdd.n476 vdd.n475 0.007
R65812 vdd.n462 vdd.n461 0.007
R65813 vdd.n303 vdd.n227 0.007
R65814 vdd.n288 vdd.n285 0.007
R65815 vdd.n238 vdd.n237 0.007
R65816 vdd.n121 vdd.n118 0.007
R65817 vdd.n157 vdd.n155 0.007
R65818 vdd.n198 vdd.n197 0.007
R65819 vdd.n116 vdd.n115 0.007
R65820 vdd.n124 vdd.n123 0.007
R65821 vdd.n359 vdd.n358 0.007
R65822 vdd.n318 vdd.n317 0.007
R65823 vdd.n332 vdd.n331 0.007
R65824 vdd.n341 vdd.n340 0.007
R65825 vdd.n6302 vdd.n6300 0.007
R65826 vdd.n6289 vdd.n6287 0.007
R65827 vdd.n6274 vdd.n6273 0.007
R65828 vdd.n5971 vdd.n5968 0.007
R65829 vdd.n5980 vdd.n5978 0.007
R65830 vdd.n5990 vdd.n5989 0.007
R65831 vdd.n5815 vdd.n5814 0.007
R65832 vdd.n5830 vdd.n5820 0.007
R65833 vdd.n5792 vdd.n5791 0.007
R65834 vdd.n6035 vdd.n6034 0.007
R65835 vdd.n6179 vdd.n6178 0.007
R65836 vdd.n6200 vdd.n6197 0.007
R65837 vdd.n6208 vdd.n6207 0.007
R65838 vdd.n6090 vdd.n6085 0.007
R65839 vdd.n6064 vdd.n6063 0.007
R65840 vdd.n6070 vdd.n6069 0.007
R65841 vdd.n5889 vdd.n5888 0.007
R65842 vdd.n5411 vdd.n5410 0.007
R65843 vdd.n5704 vdd.n5701 0.007
R65844 vdd.n5429 vdd.n5428 0.007
R65845 vdd.n5724 vdd.n5723 0.007
R65846 vdd.n5684 vdd.n5682 0.007
R65847 vdd.n5675 vdd.n5672 0.007
R65848 vdd.n5759 vdd.n5758 0.007
R65849 vdd.n5461 vdd.n5460 0.007
R65850 vdd.n5537 vdd.n5536 0.007
R65851 vdd.n5531 vdd.n5530 0.007
R65852 vdd.n5549 vdd.n5544 0.007
R65853 vdd.n5568 vdd.n5565 0.007
R65854 vdd.n5212 vdd.n5210 0.007
R65855 vdd.n5234 vdd.n5233 0.007
R65856 vdd.n5209 vdd.n5208 0.007
R65857 vdd.n5215 vdd.n5214 0.007
R65858 vdd.n5310 vdd.n5309 0.007
R65859 vdd.n5325 vdd.n5323 0.007
R65860 vdd.n5338 vdd.n5336 0.007
R65861 vdd.n5334 vdd.n5333 0.007
R65862 vdd.n5359 vdd.n5358 0.007
R65863 vdd.n4652 vdd.n4650 0.007
R65864 vdd.n5143 vdd.n5142 0.007
R65865 vdd.n5134 vdd.n5132 0.007
R65866 vdd.n5112 vdd.n5109 0.007
R65867 vdd.n4856 vdd.n4852 0.007
R65868 vdd.n5118 vdd.n5117 0.007
R65869 vdd.n5125 vdd.n5124 0.007
R65870 vdd.n4783 vdd.n4782 0.007
R65871 vdd.n4777 vdd.n4776 0.007
R65872 vdd.n4765 vdd.n4760 0.007
R65873 vdd.n4731 vdd.n4729 0.007
R65874 vdd.n5001 vdd.n4998 0.007
R65875 vdd.n4984 vdd.n4983 0.007
R65876 vdd.n5014 vdd.n5013 0.007
R65877 vdd.n5016 vdd.n5015 0.007
R65878 vdd.n4699 vdd.n4698 0.007
R65879 vdd.n4930 vdd.n4929 0.007
R65880 vdd.n4241 vdd.n4240 0.007
R65881 vdd.n4531 vdd.n4528 0.007
R65882 vdd.n4539 vdd.n4538 0.007
R65883 vdd.n4554 vdd.n4553 0.007
R65884 vdd.n4511 vdd.n4509 0.007
R65885 vdd.n4502 vdd.n4499 0.007
R65886 vdd.n4589 vdd.n4588 0.007
R65887 vdd.n4288 vdd.n4287 0.007
R65888 vdd.n4364 vdd.n4363 0.007
R65889 vdd.n4358 vdd.n4357 0.007
R65890 vdd.n4376 vdd.n4371 0.007
R65891 vdd.n4394 vdd.n4391 0.007
R65892 vdd.n4042 vdd.n4040 0.007
R65893 vdd.n4064 vdd.n4063 0.007
R65894 vdd.n4039 vdd.n4038 0.007
R65895 vdd.n4141 vdd.n4140 0.007
R65896 vdd.n4156 vdd.n4154 0.007
R65897 vdd.n4169 vdd.n4167 0.007
R65898 vdd.n4190 vdd.n4189 0.007
R65899 vdd.n2675 vdd.n2674 0.007
R65900 vdd.n36987 vdd.n36986 0.007
R65901 vdd.n37007 vdd.n37000 0.007
R65902 vdd.n37022 vdd.n37015 0.007
R65903 vdd.n38198 vdd.n38197 0.007
R65904 vdd.n38184 vdd.n38183 0.007
R65905 vdd.n38172 vdd.n38169 0.007
R65906 vdd.n31167 vdd.n31162 0.007
R65907 vdd.n29825 vdd.n29824 0.007
R65908 vdd.n30007 vdd.n30006 0.007
R65909 vdd.n29861 vdd.n29854 0.007
R65910 vdd.n27942 vdd.n27941 0.007
R65911 vdd.n28865 vdd.n28864 0.007
R65912 vdd.n27999 vdd.n27997 0.007
R65913 vdd.n29846 vdd.n29810 0.007
R65914 vdd.n29727 vdd.n29725 0.007
R65915 vdd.n30647 vdd.n30645 0.007
R65916 vdd.n27620 vdd.n27619 0.007
R65917 vdd.n27629 vdd.n27626 0.007
R65918 vdd.n27255 vdd.n27254 0.007
R65919 vdd.n27480 vdd.n27477 0.007
R65920 vdd.n27515 vdd.n27514 0.007
R65921 vdd.n27524 vdd.n27521 0.007
R65922 vdd.n27539 vdd.n27538 0.007
R65923 vdd.n27380 vdd.n27377 0.007
R65924 vdd.n27399 vdd.n27398 0.007
R65925 vdd.n27408 vdd.n27406 0.007
R65926 vdd.n27418 vdd.n27415 0.007
R65927 vdd.n27460 vdd.n27459 0.007
R65928 vdd.n27326 vdd.n27325 0.007
R65929 vdd.n26041 vdd.n26040 0.007
R65930 vdd.n26050 vdd.n26047 0.007
R65931 vdd.n25677 vdd.n25676 0.007
R65932 vdd.n25718 vdd.n25715 0.007
R65933 vdd.n25926 vdd.n25925 0.007
R65934 vdd.n25952 vdd.n25951 0.007
R65935 vdd.n25961 vdd.n25958 0.007
R65936 vdd.n25976 vdd.n25975 0.007
R65937 vdd.n25823 vdd.n25820 0.007
R65938 vdd.n25845 vdd.n25844 0.007
R65939 vdd.n25854 vdd.n25852 0.007
R65940 vdd.n25864 vdd.n25861 0.007
R65941 vdd.n25906 vdd.n25905 0.007
R65942 vdd.n25778 vdd.n25777 0.007
R65943 vdd.n25636 vdd.n25635 0.007
R65944 vdd.n25593 vdd.n25592 0.007
R65945 vdd.n25436 vdd.n25434 0.007
R65946 vdd.n25531 vdd.n25436 0.007
R65947 vdd.n25544 vdd.n25543 0.007
R65948 vdd.n25471 vdd.n25470 0.007
R65949 vdd.n30925 vdd.n30924 0.007
R65950 vdd.n30839 vdd.n30838 0.007
R65951 vdd.n30844 vdd.n30843 0.007
R65952 vdd.n30020 vdd.n30019 0.007
R65953 vdd.n30024 vdd.n30022 0.007
R65954 vdd.n30019 vdd.n30018 0.007
R65955 vdd.n29620 vdd.n29619 0.007
R65956 vdd.n7162 vdd.n7161 0.007
R65957 vdd.n27714 vdd.n27713 0.007
R65958 vdd.n27668 vdd.n27665 0.007
R65959 vdd.n27667 vdd.n27666 0.007
R65960 vdd.n26546 vdd.n26545 0.007
R65961 vdd.n31312 vdd.n31311 0.007
R65962 vdd.n30994 vdd.n30992 0.007
R65963 vdd.n30810 vdd.n30809 0.007
R65964 vdd.n31301 vdd.n31300 0.007
R65965 vdd.n31293 vdd.n31292 0.007
R65966 vdd.n31296 vdd.n31294 0.007
R65967 vdd.n7194 vdd.n7193 0.007
R65968 vdd.n26391 vdd.n26388 0.007
R65969 vdd.n26472 vdd.n26450 0.007
R65970 vdd.n7185 vdd.n7179 0.007
R65971 vdd.n29530 vdd.n29522 0.007
R65972 vdd.n31441 vdd.n31434 0.007
R65973 vdd.n30813 vdd.n30788 0.007
R65974 vdd.n26258 vdd.n26257 0.007
R65975 vdd.n29398 vdd.n29397 0.007
R65976 vdd.n32582 vdd.n32581 0.007
R65977 vdd.n32583 vdd.n32582 0.007
R65978 vdd.n30711 vdd.n30709 0.007
R65979 vdd.n3692 vdd.n2697 0.007
R65980 vdd.n3967 vdd.n3768 0.007
R65981 vdd.n2530 vdd.n2431 0.007
R65982 vdd.n2480 vdd.n2457 0.007
R65983 vdd.n3658 vdd.n3657 0.007
R65984 vdd.n3676 vdd.n3675 0.007
R65985 vdd.n3683 vdd.n3682 0.007
R65986 vdd.n3695 vdd.n3694 0.007
R65987 vdd.n4000 vdd.n3999 0.007
R65988 vdd.n3985 vdd.n3984 0.007
R65989 vdd.n3970 vdd.n3969 0.007
R65990 vdd.n3959 vdd.n3958 0.007
R65991 vdd.n3943 vdd.n3942 0.007
R65992 vdd.n2253 vdd.n2252 0.007
R65993 vdd.n2260 vdd.n2259 0.007
R65994 vdd.n2268 vdd.n2267 0.007
R65995 vdd.n2316 vdd.n2315 0.007
R65996 vdd.n2335 vdd.n2334 0.007
R65997 vdd.n2354 vdd.n2353 0.007
R65998 vdd.n2369 vdd.n2368 0.007
R65999 vdd.n2560 vdd.n2559 0.007
R66000 vdd.n2645 vdd.n2644 0.007
R66001 vdd.n2660 vdd.n2659 0.007
R66002 vdd.n2096 vdd.n2084 0.007
R66003 vdd.n1957 vdd.n1952 0.007
R66004 vdd.n1927 vdd.n1925 0.007
R66005 vdd.n1915 vdd.n1913 0.007
R66006 vdd.n1845 vdd.n1843 0.007
R66007 vdd.n1892 vdd.n1891 0.007
R66008 vdd.n1783 vdd.n1772 0.007
R66009 vdd.n31808 vdd.n31807 0.007
R66010 vdd.n31827 vdd.n31826 0.007
R66011 vdd.n31852 vdd.n31851 0.007
R66012 vdd.n31937 vdd.n31936 0.007
R66013 vdd.n31951 vdd.n31950 0.007
R66014 vdd.n32024 vdd.n32022 0.007
R66015 vdd.n32138 vdd.n32135 0.007
R66016 vdd.n32166 vdd.n32164 0.007
R66017 vdd.n32188 vdd.n32187 0.007
R66018 vdd.n32210 vdd.n32206 0.007
R66019 vdd.n32278 vdd.n32277 0.007
R66020 vdd.n32297 vdd.n32296 0.007
R66021 vdd.n32307 vdd.n32306 0.007
R66022 vdd.n32476 vdd.n32474 0.007
R66023 vdd.n32465 vdd.n32463 0.007
R66024 vdd.n31052 vdd.n31051 0.007
R66025 vdd.n31075 vdd.n31073 0.007
R66026 vdd.n31104 vdd.n31099 0.007
R66027 vdd.n31967 vdd.n31966 0.007
R66028 vdd.n32106 vdd.n32094 0.007
R66029 vdd.n32340 vdd.n32339 0.007
R66030 vdd.n32511 vdd.n32413 0.007
R66031 vdd.n7176 vdd.n7175 0.007
R66032 vdd.n30776 vdd.n30775 0.007
R66033 vdd.n12573 vdd.n12572 0.007
R66034 vdd.n12507 vdd.n12506 0.007
R66035 vdd.n10640 vdd.n10639 0.007
R66036 vdd.n10734 vdd.n10733 0.007
R66037 vdd.n12360 vdd.n12359 0.007
R66038 vdd.n12300 vdd.n12299 0.007
R66039 vdd.n10967 vdd.n10965 0.007
R66040 vdd.n11082 vdd.n11081 0.007
R66041 vdd.n12155 vdd.n11131 0.007
R66042 vdd.n11227 vdd.n11224 0.007
R66043 vdd.n12054 vdd.n12053 0.007
R66044 vdd.n11994 vdd.n11993 0.007
R66045 vdd.n11520 vdd.n11519 0.007
R66046 vdd.n11543 vdd.n11451 0.007
R66047 vdd.n11950 vdd.n11543 0.007
R66048 vdd.n13923 vdd.n13922 0.007
R66049 vdd.n14029 vdd.n8546 0.007
R66050 vdd.n14213 vdd.n14212 0.007
R66051 vdd.n14366 vdd.n14365 0.007
R66052 vdd.n14476 vdd.n14475 0.007
R66053 vdd.n13751 vdd.n13750 0.007
R66054 vdd.n9258 vdd.n9253 0.007
R66055 vdd.n13156 vdd.n9236 0.007
R66056 vdd.n13171 vdd.n9229 0.007
R66057 vdd.n9114 vdd.n9110 0.007
R66058 vdd.n13469 vdd.n13462 0.007
R66059 vdd.n8893 vdd.n8889 0.007
R66060 vdd.n11510 vdd.n11502 0.007
R66061 vdd.n10422 vdd.n10310 0.007
R66062 vdd.n13066 vdd.n13065 0.007
R66063 vdd.n9392 vdd.n9391 0.007
R66064 vdd.n9492 vdd.n9491 0.007
R66065 vdd.n12913 vdd.n12912 0.007
R66066 vdd.n12858 vdd.n12857 0.007
R66067 vdd.n9752 vdd.n9751 0.007
R66068 vdd.n9852 vdd.n9851 0.007
R66069 vdd.n12705 vdd.n12704 0.007
R66070 vdd.n12650 vdd.n12649 0.007
R66071 vdd.n10174 vdd.n10052 0.007
R66072 vdd.n13785 ldomc_0.otaldom_0.pcsm_0.vdd 0.007
R66073 ldomc_0.otaldom_0.pcsm_0.vdd vdd.n8735 0.007
R66074 vdd.n24174 vdd.n24164 0.007
R66075 vdd.n24010 vdd.n24008 0.007
R66076 vdd.n23942 vdd.n23932 0.007
R66077 vdd.n23778 vdd.n23776 0.007
R66078 vdd.n23710 vdd.n23700 0.007
R66079 vdd.n23090 vdd.n23088 0.007
R66080 vdd.n23254 vdd.n23244 0.007
R66081 vdd.n23322 vdd.n23320 0.007
R66082 vdd.n23486 vdd.n23476 0.007
R66083 vdd.n23554 vdd.n23552 0.007
R66084 vdd.n22511 vdd.n22509 0.007
R66085 vdd.n22675 vdd.n22665 0.007
R66086 vdd.n22743 vdd.n22741 0.007
R66087 vdd.n22907 vdd.n22897 0.007
R66088 vdd.n22975 vdd.n22973 0.007
R66089 vdd.n15122 vdd.n15043 0.007
R66090 vdd.n16936 vdd.n16935 0.007
R66091 vdd.n17044 vdd.n17030 0.007
R66092 vdd.n17208 vdd.n17207 0.007
R66093 vdd.n17316 vdd.n17302 0.007
R66094 vdd.n17480 vdd.n17479 0.007
R66095 vdd.n17588 vdd.n17574 0.007
R66096 vdd.n17738 vdd.n17737 0.007
R66097 vdd.n17846 vdd.n17832 0.007
R66098 vdd.n18009 vdd.n18008 0.007
R66099 vdd.n18117 vdd.n18103 0.007
R66100 vdd.n18277 vdd.n18276 0.007
R66101 vdd.n18351 vdd.n18350 0.007
R66102 vdd.n18384 vdd.n18383 0.007
R66103 vdd.n18388 vdd.n18384 0.007
R66104 vdd.n19099 vdd.n19087 0.007
R66105 vdd.n18956 vdd.n18954 0.007
R66106 vdd.n18840 vdd.n18828 0.007
R66107 vdd.n18697 vdd.n18695 0.007
R66108 vdd.n18581 vdd.n18569 0.007
R66109 vdd.n21065 vdd.n21063 0.007
R66110 vdd.n21628 vdd.n21624 0.007
R66111 vdd.n21621 vdd.n21619 0.007
R66112 vdd.n21581 vdd.n21579 0.007
R66113 vdd.n21465 vdd.n21453 0.007
R66114 vdd.n21322 vdd.n21320 0.007
R66115 vdd.n21206 vdd.n21194 0.007
R66116 vdd.n16800 vdd.n16799 0.007
R66117 vdd.n15371 vdd.n15359 0.007
R66118 vdd.n15484 vdd.n15483 0.007
R66119 vdd.n15613 vdd.n15598 0.007
R66120 vdd.n15740 vdd.n15739 0.007
R66121 vdd.n15869 vdd.n15854 0.007
R66122 vdd.n15996 vdd.n15995 0.007
R66123 vdd.n16125 vdd.n16110 0.007
R66124 vdd.n16252 vdd.n16251 0.007
R66125 vdd.n16381 vdd.n16366 0.007
R66126 vdd.n16508 vdd.n16507 0.007
R66127 vdd.n16757 vdd.n16756 0.007
R66128 bandgapmd_0.otam_1.pcsm_0.vdd vdd.n19827 0.007
R66129 vdd.n19829 bandgapmd_0.otam_1.pcsm_0.vdd 0.007
R66130 vdd.n24529 vdd.n24528 0.007
R66131 vdd.n24907 vdd.n24906 0.007
R66132 vdd.n24944 vdd.n24943 0.007
R66133 vdd.n24564 vdd.n24563 0.007
R66134 ldomc_0.vdd vdd.n38217 0.007
R66135 vdd.n31209 vdd.n31208 0.007
R66136 vdd.n26134 vdd.n26133 0.007
R66137 vdd.n31382 vdd.n31380 0.007
R66138 vdd.n30684 vdd.n30683 0.007
R66139 vdd.n27892 vdd.n27891 0.007
R66140 vdd.n28050 vdd.n28049 0.007
R66141 vdd.n25264 vdd.n7964 0.007
R66142 vdd.n33482 vdd.n33481 0.007
R66143 vdd.n33716 vdd.n33715 0.007
R66144 vdd.n967 vdd.n966 0.007
R66145 vdd.n679 vdd.n678 0.007
R66146 vdd.n913 vdd.n905 0.007
R66147 vdd.n1150 vdd.n1149 0.007
R66148 vdd.n854 vdd.n851 0.007
R66149 vdd.n225 vdd.n221 0.007
R66150 vdd.n30948 vdd.n30946 0.007
R66151 vdd.n25662 vdd.n25661 0.007
R66152 vdd.n30953 vdd.n30952 0.007
R66153 vdd.n26453 vdd.n26452 0.007
R66154 vdd.n12576 vdd.n12575 0.007
R66155 vdd.n15045 vdd.n15044 0.007
R66156 vdd.n6136 vdd.n6135 0.007
R66157 vdd.n3886 vdd.n3880 0.006
R66158 vdd.n32311 vdd.n32310 0.006
R66159 vdd.n33751 vdd.n33750 0.006
R66160 vdd.n31314 vdd.n31312 0.006
R66161 vdd.n31379 vdd.n31377 0.006
R66162 vdd.n31003 vdd.n31002 0.006
R66163 vdd.n5067 vdd.n5060 0.006
R66164 vdd.n35604 vdd.n35603 0.006
R66165 vdd.n35340 vdd.n35339 0.006
R66166 vdd.n35016 vdd.n35015 0.006
R66167 vdd.n34756 vdd.n34755 0.006
R66168 vdd.n5763 vdd.n5762 0.006
R66169 vdd.n5503 vdd.n5502 0.006
R66170 vdd.n5176 vdd.n5175 0.006
R66171 vdd.n4934 vdd.n4933 0.006
R66172 vdd.n4593 vdd.n4592 0.006
R66173 vdd.n4330 vdd.n4329 0.006
R66174 vdd.n30966 vdd.n30964 0.006
R66175 vdd.n30833 vdd.n30832 0.006
R66176 vdd.n2632 vdd.n2631 0.006
R66177 vdd.n2632 vdd.n2584 0.006
R66178 vdd.n32515 vdd.n32513 0.006
R66179 vdd.n33460 vdd.n33459 0.006
R66180 vdd.n34342 vdd.n34341 0.006
R66181 vdd.n474 vdd.n473 0.006
R66182 vdd.n196 vdd.n195 0.006
R66183 vdd.n319 vdd.n316 0.006
R66184 vdd.n6044 vdd.n6043 0.006
R66185 vdd.n5859 vdd.n5857 0.006
R66186 vdd.n27966 vdd.n27868 0.006
R66187 vdd.n35611 vdd.n35465 0.006
R66188 vdd.n29434 vdd.n29433 0.006
R66189 vdd.n29534 vdd.n29532 0.006
R66190 vdd.n32645 vdd.n32643 0.006
R66191 vdd.n31430 vdd.n31429 0.006
R66192 vdd.n31227 vdd.n31226 0.006
R66193 vdd.n26322 vdd.n26321 0.006
R66194 vdd.n26476 vdd.n26474 0.006
R66195 vdd.n33391 vdd.n33381 0.006
R66196 vdd.n33357 vdd.n33356 0.006
R66197 vdd.n33700 vdd.n33699 0.006
R66198 vdd.n33779 vdd.n33778 0.006
R66199 vdd.n34216 vdd.n34215 0.006
R66200 vdd.n34063 vdd.n34062 0.006
R66201 vdd.n35049 vdd.n35048 0.006
R66202 vdd.n35190 vdd.n35189 0.006
R66203 vdd.n35336 vdd.n35335 0.006
R66204 vdd.n34752 vdd.n34751 0.006
R66205 vdd.n675 vdd.n674 0.006
R66206 vdd.n567 vdd.n566 0.006
R66207 vdd.n180 vdd.n179 0.006
R66208 vdd.n6218 vdd.n6217 0.006
R66209 vdd.n6323 vdd.n6322 0.006
R66210 vdd.n5917 vdd.n5916 0.006
R66211 vdd.n5499 vdd.n5498 0.006
R66212 vdd.n4326 vdd.n4325 0.006
R66213 vdd.n4223 vdd.n4122 0.006
R66214 vdd.n37221 vdd.n37220 0.006
R66215 vdd.n33064 vdd.n33063 0.006
R66216 vdd.n33023 vdd.n33022 0.006
R66217 vdd.n37364 vdd.n37345 0.006
R66218 vdd.n37411 vdd.n37410 0.006
R66219 vdd.n32919 vdd.n32918 0.006
R66220 vdd.n32878 vdd.n32877 0.006
R66221 vdd.n37551 vdd.n37543 0.006
R66222 vdd.n26757 vdd.n26755 0.006
R66223 vdd.n31288 vdd.n31279 0.006
R66224 vdd.n30209 vdd.n30208 0.006
R66225 vdd.n30012 vdd.n30008 0.006
R66226 vdd.n27817 vdd.n27816 0.006
R66227 vdd.n28178 vdd.n28177 0.006
R66228 vdd.n28852 vdd.n28849 0.006
R66229 vdd.n28925 vdd.n28924 0.006
R66230 vdd.n28933 vdd.n28928 0.006
R66231 vdd.n28041 vdd.n28040 0.006
R66232 vdd.n28008 vdd.n28006 0.006
R66233 vdd.n27947 vdd.n27944 0.006
R66234 vdd.n27926 vdd.n27924 0.006
R66235 vdd.n29736 vdd.n29734 0.006
R66236 vdd.n30634 vdd.n30631 0.006
R66237 vdd.n30626 vdd.n30624 0.006
R66238 vdd.n30536 vdd.n30535 0.006
R66239 vdd.n30524 vdd.n30521 0.006
R66240 vdd.n27348 vdd.n27347 0.006
R66241 vdd.n31014 vdd.n31013 0.006
R66242 vdd.n25800 vdd.n25799 0.006
R66243 vdd.n25441 vdd.n25437 0.006
R66244 vdd.n31334 vdd.n31333 0.006
R66245 vdd.n32601 vdd.n32600 0.006
R66246 vdd.n29376 vdd.n29375 0.006
R66247 vdd.n26237 vdd.n26236 0.006
R66248 vdd.n25343 vdd.n25342 0.006
R66249 vdd.n31246 vdd.n31245 0.006
R66250 vdd.n26467 vdd.n26458 0.006
R66251 vdd.n29513 vdd.n29504 0.006
R66252 vdd.n27673 vdd.n27668 0.006
R66253 vdd.n29578 vdd.n29573 0.006
R66254 vdd.n30883 vdd.n30878 0.006
R66255 vdd.n2506 vdd.n2505 0.006
R66256 vdd.n1861 vdd.n1858 0.006
R66257 vdd.n27241 vdd.n27240 0.006
R66258 vdd.n31745 vdd.n31744 0.006
R66259 vdd.n31762 vdd.n31761 0.006
R66260 vdd.n31869 vdd.n31868 0.006
R66261 vdd.n31894 vdd.n31881 0.006
R66262 vdd.n32043 vdd.n32040 0.006
R66263 vdd.n32116 vdd.n32111 0.006
R66264 vdd.n32233 vdd.n32232 0.006
R66265 vdd.n32259 vdd.n32254 0.006
R66266 vdd.n32473 vdd.n32471 0.006
R66267 vdd.n31121 vdd.n31120 0.006
R66268 vdd.n31181 vdd.n31180 0.006
R66269 vdd.n10548 vdd.n10547 0.006
R66270 vdd.n12448 vdd.n12447 0.006
R66271 vdd.n12408 vdd.n10697 0.006
R66272 vdd.n10836 vdd.n10810 0.006
R66273 vdd.n10891 vdd.n10872 0.006
R66274 vdd.n12247 vdd.n12246 0.006
R66275 vdd.n12215 vdd.n11039 0.006
R66276 vdd.n11174 vdd.n11151 0.006
R66277 vdd.n12110 vdd.n12109 0.006
R66278 vdd.n11345 vdd.n11319 0.006
R66279 vdd.n11400 vdd.n11381 0.006
R66280 vdd.n11494 vdd.n11493 0.006
R66281 vdd.n11534 vdd.n11533 0.006
R66282 vdd.n13939 vdd.n8638 0.006
R66283 vdd.n14028 vdd.n14027 0.006
R66284 vdd.n14229 vdd.n8416 0.006
R66285 vdd.n14315 vdd.n14314 0.006
R66286 vdd.n14536 vdd.n8193 0.006
R66287 vdd.n13750 vdd.n8759 0.006
R66288 vdd.n11612 vdd.n9250 0.006
R66289 vdd.n13157 vdd.n9231 0.006
R66290 vdd.n9117 vdd.n9116 0.006
R66291 vdd.n13451 vdd.n13450 0.006
R66292 vdd.n8896 vdd.n8895 0.006
R66293 vdd.n11610 vdd.n9252 0.006
R66294 vdd.n11495 vdd.n11465 0.006
R66295 vdd.n11594 vdd.n11584 0.006
R66296 vdd.n10176 vdd.n10175 0.006
R66297 vdd.n10252 vdd.n10128 0.006
R66298 vdd.n10410 vdd.n10409 0.006
R66299 vdd.n9302 vdd.n9295 0.006
R66300 vdd.n9396 vdd.n9393 0.006
R66301 vdd.n12966 vdd.n9458 0.006
R66302 vdd.n9587 vdd.n9583 0.006
R66303 vdd.n9662 vdd.n9656 0.006
R66304 vdd.n9756 vdd.n9753 0.006
R66305 vdd.n12758 vdd.n9818 0.006
R66306 vdd.n9947 vdd.n9943 0.006
R66307 vdd.n10022 vdd.n10016 0.006
R66308 vdd.n12600 vdd.n10053 0.006
R66309 vdd.n22214 vdd.n22213 0.006
R66310 vdd.n22077 vdd.n22067 0.006
R66311 vdd.n22329 vdd.n22328 0.006
R66312 vdd.n22326 vdd.n22325 0.006
R66313 vdd.n24322 vdd.n24321 0.006
R66314 vdd.n24301 vdd.n24300 0.006
R66315 vdd.n24298 vdd.n24297 0.006
R66316 vdd.n24205 vdd.n24204 0.006
R66317 vdd.n22470 vdd.n22469 0.006
R66318 vdd.n22377 vdd.n22376 0.006
R66319 vdd.n16903 vdd.n16889 0.006
R66320 vdd.n17077 vdd.n17076 0.006
R66321 vdd.n17175 vdd.n17161 0.006
R66322 vdd.n17349 vdd.n17348 0.006
R66323 vdd.n17447 vdd.n17433 0.006
R66324 vdd.n17607 vdd.n17606 0.006
R66325 vdd.n17705 vdd.n17691 0.006
R66326 vdd.n17878 vdd.n17877 0.006
R66327 vdd.n17976 vdd.n17962 0.006
R66328 vdd.n18150 vdd.n18149 0.006
R66329 vdd.n18246 vdd.n18233 0.006
R66330 vdd.n18314 vdd.n18313 0.006
R66331 vdd.n18372 vdd.n18370 0.006
R66332 vdd.n19071 vdd.n19069 0.006
R66333 vdd.n18974 vdd.n18972 0.006
R66334 vdd.n18812 vdd.n18810 0.006
R66335 vdd.n18715 vdd.n18713 0.006
R66336 vdd.n18553 vdd.n18551 0.006
R66337 vdd.n21063 vdd.n21061 0.006
R66338 vdd.n21678 vdd.n21677 0.006
R66339 vdd.n21599 vdd.n21597 0.006
R66340 vdd.n21437 vdd.n21435 0.006
R66341 vdd.n21340 vdd.n21338 0.006
R66342 vdd.n21178 vdd.n21176 0.006
R66343 vdd.n21691 vdd.n21690 0.006
R66344 vdd.n16806 vdd.n16805 0.006
R66345 vdd.n21699 vdd.n18431 0.006
R66346 vdd.n16772 vdd.n16771 0.006
R66347 vdd.n16790 vdd.n16789 0.006
R66348 vdd.n15386 vdd.n15385 0.006
R66349 vdd.n15466 vdd.n15448 0.006
R66350 vdd.n15631 vdd.n15630 0.006
R66351 vdd.n15722 vdd.n15704 0.006
R66352 vdd.n15887 vdd.n15886 0.006
R66353 vdd.n15978 vdd.n15960 0.006
R66354 vdd.n16143 vdd.n16142 0.006
R66355 vdd.n16234 vdd.n16216 0.006
R66356 vdd.n16399 vdd.n16398 0.006
R66357 vdd.n16490 vdd.n16472 0.006
R66358 vdd.n16752 vdd.n16743 0.006
R66359 vdd.n24745 vdd.n24744 0.006
R66360 vdd.n24758 vdd.n24750 0.006
R66361 vdd.n24833 vdd.n24832 0.006
R66362 vdd.n25254 vdd.n24833 0.006
R66363 vdd.n25251 vdd.n25250 0.006
R66364 vdd.n25250 bandgapmd_0.bg_pmosm_0.vdd 0.006
R66365 vdd.n25176 vdd.n25166 0.006
R66366 vdd.n25161 vdd.n25160 0.006
R66367 vdd.n772 vdd.n771 0.006
R66368 vdd.n2006 vdd.n2005 0.006
R66369 vdd.n771 vdd.n770 0.006
R66370 vdd.n2562 vdd.n2560 0.006
R66371 vdd.n2562 vdd.n2561 0.006
R66372 vdd.n30797 vdd.n30796 0.006
R66373 vdd.n24903 vdd.n24902 0.006
R66374 vdd.n30665 vdd.n30653 0.006
R66375 vdd.n28905 vdd.n28904 0.006
R66376 vdd.n28877 vdd.n28107 0.006
R66377 vdd.n684 vdd.n683 0.006
R66378 vdd.n1162 vdd.n1161 0.006
R66379 vdd.n866 vdd.n863 0.006
R66380 vdd.n30959 vdd.n30958 0.006
R66381 vdd.n34345 vdd.n34344 0.006
R66382 vdd.n26081 vdd.n26080 0.005
R66383 vdd.n27659 vdd.n27658 0.005
R66384 vdd.n30591 vdd.n30590 0.005
R66385 vdd.n35223 vdd.n35222 0.005
R66386 vdd.n34636 vdd.n34635 0.005
R66387 vdd.n5383 vdd.n5382 0.005
R66388 vdd.n4704 vdd.n4703 0.005
R66389 vdd.n4213 vdd.n4212 0.005
R66390 vdd.n35222 vdd.n35221 0.005
R66391 vdd.n34635 vdd.n34634 0.005
R66392 vdd.n282 vdd.n281 0.005
R66393 vdd.n5382 vdd.n5381 0.005
R66394 vdd.n4703 vdd.n4702 0.005
R66395 vdd.n4212 vdd.n4211 0.005
R66396 vdd.n11772 vdd.n11666 0.005
R66397 vdd.n11806 vdd.n11804 0.005
R66398 vdd.n21864 vdd.n21859 0.005
R66399 vdd.n21897 vdd.n21895 0.005
R66400 vdd.n26277 vdd.n26276 0.005
R66401 vdd.n29423 vdd.n29422 0.005
R66402 vdd.n6353 vdd.n6352 0.005
R66403 vdd.n35465 vdd.n35358 0.005
R66404 vdd.n6136 vdd.n6046 0.005
R66405 vdd.n680 vdd.n679 0.005
R66406 vdd.n968 vdd.n967 0.005
R66407 vdd.n1151 vdd.n1150 0.005
R66408 vdd.n854 vdd.n853 0.005
R66409 vdd.n33483 vdd.n33482 0.005
R66410 vdd.n32315 vdd.n32311 0.005
R66411 vdd.n25483 vdd.n25481 0.005
R66412 vdd.n29504 vdd.n29503 0.005
R66413 vdd.n10482 vdd.n10123 0.005
R66414 vdd.n15053 vdd.n15051 0.005
R66415 vdd.n32375 vdd.n32369 0.005
R66416 vdd.n32106 vdd.n32105 0.005
R66417 vdd.n32528 vdd.n32527 0.005
R66418 vdd.n27996 vdd.n27858 0.005
R66419 vdd.n24524 vdd.n24519 0.005
R66420 vdd.n35609 vdd.n35608 0.005
R66421 vdd.n35352 vdd.n35351 0.005
R66422 vdd.n35021 vdd.n35020 0.005
R66423 vdd.n34768 vdd.n34767 0.005
R66424 vdd.n5768 vdd.n5767 0.005
R66425 vdd.n5515 vdd.n5514 0.005
R66426 vdd.n4598 vdd.n4597 0.005
R66427 vdd.n4342 vdd.n4341 0.005
R66428 vdd.n24549 vdd.n24548 0.005
R66429 vdd.n7187 vdd.n7186 0.005
R66430 vdd.n32680 vdd.n32679 0.005
R66431 vdd.n29099 vdd.n29098 0.005
R66432 vdd.n2888 vdd.n2881 0.005
R66433 vdd.n2900 vdd.n2898 0.005
R66434 vdd.n3069 vdd.n3062 0.005
R66435 vdd.n3081 vdd.n3079 0.005
R66436 vdd.n3250 vdd.n3243 0.005
R66437 vdd.n3262 vdd.n3260 0.005
R66438 vdd.n3431 vdd.n3424 0.005
R66439 vdd.n3443 vdd.n3441 0.005
R66440 vdd.n3612 vdd.n3605 0.005
R66441 vdd.n3624 vdd.n3622 0.005
R66442 vdd.n33454 vdd.n33453 0.005
R66443 vdd.n33681 vdd.n33680 0.005
R66444 vdd.n33846 vdd.n33844 0.005
R66445 vdd.n34158 vdd.n34157 0.005
R66446 vdd.n34163 vdd.n34162 0.005
R66447 vdd.n35312 vdd.n35311 0.005
R66448 vdd.n35356 vdd.n35355 0.005
R66449 vdd.n34772 vdd.n34771 0.005
R66450 vdd.n34736 vdd.n34735 0.005
R66451 vdd.n1146 vdd.n1145 0.005
R66452 vdd.n847 vdd.n845 0.005
R66453 vdd.n468 vdd.n467 0.005
R66454 vdd.n186 vdd.n185 0.005
R66455 vdd.n379 vdd.n378 0.005
R66456 vdd.n374 vdd.n373 0.005
R66457 vdd.n5864 vdd.n5863 0.005
R66458 vdd.n6041 vdd.n6040 0.005
R66459 vdd.n5847 vdd.n5846 0.005
R66460 vdd.n5922 vdd.n5921 0.005
R66461 vdd.n5519 vdd.n5518 0.005
R66462 vdd.n5483 vdd.n5482 0.005
R66463 vdd.n4906 vdd.n4905 0.005
R66464 vdd.n4346 vdd.n4345 0.005
R66465 vdd.n4310 vdd.n4309 0.005
R66466 vdd.n36033 vdd.n36023 0.005
R66467 vdd.n36049 vdd.n36047 0.005
R66468 vdd.n36264 vdd.n36254 0.005
R66469 vdd.n36280 vdd.n36278 0.005
R66470 vdd.n36495 vdd.n36485 0.005
R66471 vdd.n36511 vdd.n36509 0.005
R66472 vdd.n36726 vdd.n36716 0.005
R66473 vdd.n36742 vdd.n36740 0.005
R66474 vdd.n36957 vdd.n36947 0.005
R66475 vdd.n37048 vdd.n37047 0.005
R66476 vdd.n33272 vdd.n33258 0.005
R66477 vdd.n37119 vdd.n37102 0.005
R66478 vdd.n33177 vdd.n33176 0.005
R66479 vdd.n37153 vdd.n37152 0.005
R66480 vdd.n33139 vdd.n33121 0.005
R66481 vdd.n37213 vdd.n37210 0.005
R66482 vdd.n33099 vdd.n33098 0.005
R66483 vdd.n37285 vdd.n37265 0.005
R66484 vdd.n37315 vdd.n37314 0.005
R66485 vdd.n32982 vdd.n32968 0.005
R66486 vdd.n32963 vdd.n32962 0.005
R66487 vdd.n37457 vdd.n37456 0.005
R66488 vdd.n37497 vdd.n37496 0.005
R66489 vdd.n35673 vdd.n35660 0.005
R66490 vdd.n37550 vdd.n37546 0.005
R66491 vdd.n38215 vdd.n38214 0.005
R66492 vdd.n38174 vdd.n38172 0.005
R66493 vdd.n38028 vdd.n38026 0.005
R66494 vdd.n38012 vdd.n38002 0.005
R66495 vdd.n37797 vdd.n37795 0.005
R66496 vdd.n37781 vdd.n37771 0.005
R66497 vdd.n28223 vdd.n28213 0.005
R66498 vdd.n28239 vdd.n28237 0.005
R66499 vdd.n28454 vdd.n28444 0.005
R66500 vdd.n28470 vdd.n28468 0.005
R66501 vdd.n28685 vdd.n28675 0.005
R66502 vdd.n28701 vdd.n28699 0.005
R66503 vdd.n1662 vdd.n1660 0.005
R66504 vdd.n1650 vdd.n1643 0.005
R66505 vdd.n1481 vdd.n1479 0.005
R66506 vdd.n1469 vdd.n1462 0.005
R66507 vdd.n1300 vdd.n1298 0.005
R66508 vdd.n26766 vdd.n26764 0.005
R66509 vdd.n26935 vdd.n26928 0.005
R66510 vdd.n26947 vdd.n26945 0.005
R66511 vdd.n27116 vdd.n27109 0.005
R66512 vdd.n27128 vdd.n27126 0.005
R66513 vdd.n31161 vdd.n31158 0.005
R66514 vdd.n30683 vdd.n30682 0.005
R66515 vdd.n29747 vdd.n29743 0.005
R66516 vdd.n27891 vdd.n27890 0.005
R66517 vdd.n27797 vdd.n27796 0.005
R66518 vdd.n28054 vdd.n28050 0.005
R66519 vdd.n28074 vdd.n28073 0.005
R66520 vdd.n28127 vdd.n28126 0.005
R66521 vdd.n28128 vdd.n28127 0.005
R66522 vdd.n30247 vdd.n30240 0.005
R66523 vdd.n28836 vdd.n28833 0.005
R66524 vdd.n28837 vdd.n28836 0.005
R66525 vdd.n28849 vdd.n28846 0.005
R66526 vdd.n28913 vdd.n28910 0.005
R66527 vdd.n28946 vdd.n28941 0.005
R66528 vdd.n28947 vdd.n28946 0.005
R66529 vdd.n28992 vdd.n28991 0.005
R66530 vdd.n29005 vdd.n29004 0.005
R66531 vdd.n28040 vdd.n28039 0.005
R66532 vdd.n28039 vdd.n28037 0.005
R66533 vdd.n28031 vdd.n28029 0.005
R66534 vdd.n28022 vdd.n28019 0.005
R66535 vdd.n28019 vdd.n28017 0.005
R66536 vdd.n28010 vdd.n28008 0.005
R66537 vdd.n27956 vdd.n27953 0.005
R66538 vdd.n27924 vdd.n27921 0.005
R66539 vdd.n29903 vdd.n29898 0.005
R66540 vdd.n29905 vdd.n29904 0.005
R66541 vdd.n29805 vdd.n29802 0.005
R66542 vdd.n29785 vdd.n29783 0.005
R66543 vdd.n29773 vdd.n29770 0.005
R66544 vdd.n29770 vdd.n29768 0.005
R66545 vdd.n29738 vdd.n29736 0.005
R66546 vdd.n30643 vdd.n30640 0.005
R66547 vdd.n30631 vdd.n30630 0.005
R66548 vdd.n30617 vdd.n30615 0.005
R66549 vdd.n25531 vdd.n25530 0.005
R66550 vdd.n30875 vdd.n30874 0.005
R66551 vdd.n30788 vdd.n30787 0.005
R66552 vdd.n30142 vdd.n30141 0.005
R66553 vdd.n32622 vdd.n32621 0.005
R66554 vdd.n29539 vdd.n29538 0.005
R66555 vdd.n29522 vdd.n29521 0.005
R66556 vdd.n29356 vdd.n29355 0.005
R66557 vdd.n26487 vdd.n26486 0.005
R66558 vdd.n26566 vdd.n26565 0.005
R66559 vdd.n31005 vdd.n31004 0.005
R66560 vdd.n31220 vdd.n31219 0.005
R66561 vdd.n31215 vdd.n31199 0.005
R66562 vdd.n26132 vdd.n26131 0.005
R66563 vdd.n25370 vdd.n25369 0.005
R66564 vdd.n25376 vdd.n25374 0.005
R66565 vdd.n32809 vdd.n6420 0.005
R66566 vdd.n32804 vdd.n6478 0.005
R66567 vdd.n32799 vdd.n6535 0.005
R66568 vdd.n32778 vdd.n6759 0.005
R66569 vdd.n32772 vdd.n6818 0.005
R66570 vdd.n32766 vdd.n6874 0.005
R66571 vdd.n32760 vdd.n6930 0.005
R66572 vdd.n32754 vdd.n6986 0.005
R66573 vdd.n32748 vdd.n7042 0.005
R66574 vdd.n32737 vdd.n7199 0.005
R66575 vdd.n31235 vdd.n31234 0.005
R66576 vdd.n30804 vdd.n30803 0.005
R66577 vdd.n32807 vdd.n6445 0.005
R66578 vdd.n32802 vdd.n6502 0.005
R66579 vdd.n32796 vdd.n6559 0.005
R66580 vdd.n32790 vdd.n6611 0.005
R66581 vdd.n32775 vdd.n6785 0.005
R66582 vdd.n26127 vdd.n26126 0.005
R66583 vdd.n26137 vdd.n26136 0.005
R66584 vdd.n25376 vdd.n25375 0.005
R66585 vdd.n26391 vdd.n26387 0.005
R66586 vdd.n26467 vdd.n26460 0.005
R66587 vdd.n7185 vdd.n7180 0.005
R66588 vdd.n29513 vdd.n29506 0.005
R66589 vdd.n26258 vdd.n26254 0.005
R66590 vdd.n27673 vdd.n27671 0.005
R66591 vdd.n29398 vdd.n29394 0.005
R66592 vdd.n29578 vdd.n29576 0.005
R66593 vdd.n30024 vdd.n30023 0.005
R66594 vdd.n32583 vdd.n32577 0.005
R66595 vdd.n30711 vdd.n30707 0.005
R66596 vdd.n30883 vdd.n30881 0.005
R66597 vdd.n3673 vdd.n2728 0.005
R66598 vdd.n3997 vdd.n3746 0.005
R66599 vdd.n2624 vdd.n2590 0.005
R66600 vdd.n3687 vdd.n3684 0.005
R66601 vdd.n3693 vdd.n3692 0.005
R66602 vdd.n3712 vdd.n3711 0.005
R66603 vdd.n4013 vdd.n4012 0.005
R66604 vdd.n3998 vdd.n3997 0.005
R66605 vdd.n3966 vdd.n3963 0.005
R66606 vdd.n3947 vdd.n3944 0.005
R66607 vdd.n3878 vdd.n3877 0.005
R66608 vdd.n2264 vdd.n2261 0.005
R66609 vdd.n2266 vdd.n2265 0.005
R66610 vdd.n2285 vdd.n2284 0.005
R66611 vdd.n2303 vdd.n2298 0.005
R66612 vdd.n2322 vdd.n2317 0.005
R66613 vdd.n2364 vdd.n2361 0.005
R66614 vdd.n2393 vdd.n2392 0.005
R66615 vdd.n2545 vdd.n2544 0.005
R66616 vdd.n2519 vdd.n2518 0.005
R66617 vdd.n2497 vdd.n2490 0.005
R66618 vdd.n2664 vdd.n2661 0.005
R66619 vdd.n2000 vdd.n1980 0.005
R66620 vdd.n1991 vdd.n1990 0.005
R66621 vdd.n2083 vdd.n2082 0.005
R66622 vdd.n1922 vdd.n1919 0.005
R66623 vdd.n1896 vdd.n1893 0.005
R66624 vdd.n1885 vdd.n1884 0.005
R66625 vdd.n1884 vdd.n1882 0.005
R66626 vdd.n1848 vdd.n1846 0.005
R66627 vdd.n1820 vdd.n1810 0.005
R66628 vdd.n1820 vdd.n1811 0.005
R66629 vdd.n31934 vdd.n31933 0.005
R66630 vdd.n26196 vdd.n26193 0.005
R66631 vdd.n26601 vdd.n26600 0.005
R66632 vdd.n26706 vdd.n26691 0.005
R66633 vdd.n26330 vdd.n26325 0.005
R66634 vdd.n26402 vdd.n26397 0.005
R66635 vdd.n31761 vdd.n31760 0.005
R66636 vdd.n31767 vdd.n31762 0.005
R66637 vdd.n31799 vdd.n31794 0.005
R66638 vdd.n31850 vdd.n31849 0.005
R66639 vdd.n31897 vdd.n31894 0.005
R66640 vdd.n31900 vdd.n31897 0.005
R66641 vdd.n31912 vdd.n31907 0.005
R66642 vdd.n31916 vdd.n31915 0.005
R66643 vdd.n31962 vdd.n31959 0.005
R66644 vdd.n31976 vdd.n31973 0.005
R66645 vdd.n31994 vdd.n31993 0.005
R66646 vdd.n32013 vdd.n32011 0.005
R66647 vdd.n32045 vdd.n32044 0.005
R66648 vdd.n32047 vdd.n32045 0.005
R66649 vdd.n32050 vdd.n32047 0.005
R66650 vdd.n32055 vdd.n32053 0.005
R66651 vdd.n32084 vdd.n32079 0.005
R66652 vdd.n32149 vdd.n32144 0.005
R66653 vdd.n32205 vdd.n32204 0.005
R66654 vdd.n32262 vdd.n32259 0.005
R66655 vdd.n32265 vdd.n32262 0.005
R66656 vdd.n32284 vdd.n32279 0.005
R66657 vdd.n32287 vdd.n32284 0.005
R66658 vdd.n32288 vdd.n32287 0.005
R66659 vdd.n32318 vdd.n32315 0.005
R66660 vdd.n32334 vdd.n32331 0.005
R66661 vdd.n32354 vdd.n32353 0.005
R66662 vdd.n32368 vdd.n32366 0.005
R66663 vdd.n32383 vdd.n32381 0.005
R66664 vdd.n32531 vdd.n32529 0.005
R66665 vdd.n32524 vdd.n32523 0.005
R66666 vdd.n32498 vdd.n32495 0.005
R66667 vdd.n32459 vdd.n32457 0.005
R66668 vdd.n31098 vdd.n31097 0.005
R66669 vdd.n31996 vdd.n31995 0.005
R66670 vdd.n32209 vdd.n32208 0.005
R66671 vdd.n32310 vdd.n32309 0.005
R66672 vdd.n31296 vdd.n31295 0.005
R66673 vdd.n32809 vdd.n6412 0.005
R66674 vdd.n32807 vdd.n6442 0.005
R66675 vdd.n32804 vdd.n6472 0.005
R66676 vdd.n32802 vdd.n6499 0.005
R66677 vdd.n32799 vdd.n6526 0.005
R66678 vdd.n32796 vdd.n6556 0.005
R66679 vdd.n32793 vdd.n6582 0.005
R66680 vdd.n32778 vdd.n6751 0.005
R66681 vdd.n32775 vdd.n6782 0.005
R66682 vdd.n32772 vdd.n6810 0.005
R66683 vdd.n32769 vdd.n6839 0.005
R66684 vdd.n32766 vdd.n6865 0.005
R66685 vdd.n32763 vdd.n6895 0.005
R66686 vdd.n32760 vdd.n6921 0.005
R66687 vdd.n32757 vdd.n6951 0.005
R66688 vdd.n32754 vdd.n6977 0.005
R66689 vdd.n32751 vdd.n7008 0.005
R66690 vdd.n32748 vdd.n7033 0.005
R66691 vdd.n32737 vdd.n7189 0.005
R66692 vdd.n25332 vdd.n7260 0.005
R66693 vdd.n12496 vdd.n12495 0.005
R66694 vdd.n12464 vdd.n10608 0.005
R66695 vdd.n10745 vdd.n10744 0.005
R66696 vdd.n10781 vdd.n10779 0.005
R66697 vdd.n10902 vdd.n10899 0.005
R66698 vdd.n10978 vdd.n10977 0.005
R66699 vdd.n12197 vdd.n12196 0.005
R66700 vdd.n12157 vdd.n11125 0.005
R66701 vdd.n11255 vdd.n11254 0.005
R66702 vdd.n11289 vdd.n11287 0.005
R66703 vdd.n11411 vdd.n11408 0.005
R66704 vdd.n11953 vdd.n11451 0.005
R66705 vdd.n13885 vdd.n13884 0.005
R66706 vdd.n14084 vdd.n14083 0.005
R66707 vdd.n14174 vdd.n14173 0.005
R66708 vdd.n8328 vdd.n8309 0.005
R66709 vdd.n14473 vdd.n8229 0.005
R66710 vdd.n13797 vdd.n13796 0.005
R66711 vdd.n13741 vdd.n8789 0.005
R66712 vdd.n13140 vdd.n9251 0.005
R66713 vdd.n13172 vdd.n9196 0.005
R66714 vdd.n13312 vdd.n13311 0.005
R66715 vdd.n13463 vdd.n8974 0.005
R66716 vdd.n13604 vdd.n13603 0.005
R66717 vdd.n10220 vdd.n10216 0.005
R66718 vdd.n10286 vdd.n10283 0.005
R66719 vdd.n10424 vdd.n10304 0.005
R66720 vdd.n13055 vdd.n13054 0.005
R66721 vdd.n9379 vdd.n9378 0.005
R66722 vdd.n9505 vdd.n9504 0.005
R66723 vdd.n12924 vdd.n9548 0.005
R66724 vdd.n12847 vdd.n12846 0.005
R66725 vdd.n9739 vdd.n9738 0.005
R66726 vdd.n9865 vdd.n9864 0.005
R66727 vdd.n12716 vdd.n9908 0.005
R66728 vdd.n12639 vdd.n12638 0.005
R66729 vdd.n12620 vdd.n10053 0.005
R66730 vdd.n11773 vdd.n11772 0.005
R66731 vdd.n11735 vdd.n11734 0.005
R66732 vdd.n11829 vdd.n11814 0.005
R66733 vdd.n11874 vdd.n11804 0.005
R66734 vdd.n11912 vdd.n11663 0.005
R66735 vdd.n13212 vdd.n13211 0.005
R66736 vdd.n13252 vdd.n9174 0.005
R66737 vdd.n14401 vdd.n14400 0.005
R66738 vdd.n14402 vdd.n8279 0.005
R66739 vdd.n14680 vdd.n8116 0.005
R66740 vdd.n14709 vdd.n14708 0.005
R66741 vdd.n14794 vdd.n14793 0.005
R66742 vdd.n14796 vdd.n14795 0.005
R66743 vdd.n14852 vdd.n8027 0.005
R66744 vdd.n14882 vdd.n14881 0.005
R66745 vdd.n22349 vdd.n22346 0.005
R66746 vdd.n22065 vdd.n22062 0.005
R66747 vdd.n22322 vdd.n22311 0.005
R66748 vdd.n22307 vdd.n22295 0.005
R66749 vdd.n24337 vdd.n24327 0.005
R66750 vdd.n24310 vdd.n24309 0.005
R66751 vdd.n24294 vdd.n24283 0.005
R66752 vdd.n24279 vdd.n24267 0.005
R66753 vdd.n24220 vdd.n24210 0.005
R66754 vdd.n24108 vdd.n24106 0.005
R66755 vdd.n24068 vdd.n24066 0.005
R66756 vdd.n23876 vdd.n23874 0.005
R66757 vdd.n23836 vdd.n23834 0.005
R66758 vdd.n23644 vdd.n23642 0.005
R66759 vdd.n23148 vdd.n23146 0.005
R66760 vdd.n23188 vdd.n23186 0.005
R66761 vdd.n23380 vdd.n23378 0.005
R66762 vdd.n23420 vdd.n23418 0.005
R66763 vdd.n23612 vdd.n23610 0.005
R66764 vdd.n22569 vdd.n22567 0.005
R66765 vdd.n22609 vdd.n22607 0.005
R66766 vdd.n22801 vdd.n22799 0.005
R66767 vdd.n22841 vdd.n22839 0.005
R66768 vdd.n23033 vdd.n23031 0.005
R66769 vdd.n22466 vdd.n22455 0.005
R66770 vdd.n22451 vdd.n22439 0.005
R66771 vdd.n22392 vdd.n22382 0.005
R66772 vdd.n22365 vdd.n22364 0.005
R66773 vdd.n16952 vdd.n16951 0.005
R66774 vdd.n17028 vdd.n17014 0.005
R66775 vdd.n17224 vdd.n17223 0.005
R66776 vdd.n17300 vdd.n17286 0.005
R66777 vdd.n17496 vdd.n17495 0.005
R66778 vdd.n17572 vdd.n17558 0.005
R66779 vdd.n17754 vdd.n17753 0.005
R66780 vdd.n17830 vdd.n17816 0.005
R66781 vdd.n18025 vdd.n18024 0.005
R66782 vdd.n18101 vdd.n18087 0.005
R66783 vdd.n18292 vdd.n18291 0.005
R66784 vdd.n18383 vdd.n18382 0.005
R66785 vdd.n19115 vdd.n19103 0.005
R66786 vdd.n18940 vdd.n18938 0.005
R66787 vdd.n18856 vdd.n18844 0.005
R66788 vdd.n18681 vdd.n18679 0.005
R66789 vdd.n18597 vdd.n18585 0.005
R66790 vdd.n21047 vdd.n21045 0.005
R66791 vdd.n21092 vdd.n21079 0.005
R66792 vdd.n21683 vdd.n21682 0.005
R66793 vdd.n21565 vdd.n21563 0.005
R66794 vdd.n21481 vdd.n21469 0.005
R66795 vdd.n21306 vdd.n21304 0.005
R66796 vdd.n21222 vdd.n21210 0.005
R66797 vdd.n16787 vdd.n16786 0.005
R66798 vdd.n15279 vdd.n15278 0.005
R66799 vdd.n15357 vdd.n15344 0.005
R66800 vdd.n15501 vdd.n15500 0.005
R66801 vdd.n15596 vdd.n15581 0.005
R66802 vdd.n15757 vdd.n15756 0.005
R66803 vdd.n15852 vdd.n15837 0.005
R66804 vdd.n16013 vdd.n16012 0.005
R66805 vdd.n16108 vdd.n16093 0.005
R66806 vdd.n16269 vdd.n16268 0.005
R66807 vdd.n16364 vdd.n16349 0.005
R66808 vdd.n16525 vdd.n16524 0.005
R66809 vdd.n16753 vdd.n16752 0.005
R66810 vdd.n20644 vdd.n20629 0.005
R66811 vdd.n20628 vdd.n20627 0.005
R66812 vdd.n20407 vdd.n20392 0.005
R66813 vdd.n20385 vdd.n20384 0.005
R66814 vdd.n20273 vdd.n20271 0.005
R66815 vdd.n20270 vdd.n20269 0.005
R66816 vdd.n20171 vdd.n20156 0.005
R66817 vdd.n20149 vdd.n20148 0.005
R66818 vdd.n19422 vdd.n19421 0.005
R66819 vdd.n19435 vdd.n19423 0.005
R66820 vdd.n21864 vdd.n21863 0.005
R66821 vdd.n21812 vdd.n21810 0.005
R66822 vdd.n21920 vdd.n21905 0.005
R66823 vdd.n21965 vdd.n21895 0.005
R66824 vdd.n21755 vdd.n21749 0.005
R66825 vdd.n24524 vdd.n24523 0.005
R66826 vdd.n25030 vdd.n25028 0.005
R66827 vdd.n25022 vdd.n25019 0.005
R66828 vdd.n24916 vdd.n24915 0.005
R66829 vdd.n24605 vdd.n24603 0.005
R66830 vdd.n24597 vdd.n24595 0.005
R66831 vdd.n24732 vdd.n24730 0.005
R66832 vdd.n24770 vdd.n24762 0.005
R66833 vdd.n24822 vdd.n24820 0.005
R66834 vdd.n25240 vdd.n25238 0.005
R66835 vdd.n25188 vdd.n25180 0.005
R66836 vdd.n25150 vdd.n25148 0.005
R66837 vdd.n2100 vdd.n2068 0.005
R66838 vdd.n2100 vdd.n2099 0.005
R66839 vdd.n25920 vdd.n25707 0.005
R66840 vdd.n881 vdd.n880 0.005
R66841 vdd.n31310 vdd.n31309 0.005
R66842 vdd.n4594 vdd.n4593 0.005
R66843 vdd.n4331 vdd.n4330 0.005
R66844 vdd.n5177 vdd.n5176 0.005
R66845 vdd.n4935 vdd.n4934 0.005
R66846 vdd.n5764 vdd.n5763 0.005
R66847 vdd.n5504 vdd.n5503 0.005
R66848 vdd.n35017 vdd.n35016 0.005
R66849 vdd.n34757 vdd.n34756 0.005
R66850 vdd.n35605 vdd.n35604 0.005
R66851 vdd.n35341 vdd.n35340 0.005
R66852 vdd.n205 vdd.n204 0.005
R66853 vdd.n306 vdd.n219 0.005
R66854 vdd.n29396 vdd.n29395 0.005
R66855 vdd.n26256 vdd.n26255 0.005
R66856 vdd.n24931 vdd.n24930 0.005
R66857 vdd.n1887 vdd.n1218 0.005
R66858 vdd.n27488 vdd.n27486 0.005
R66859 vdd.n31390 vdd.n31389 0.005
R66860 vdd.n30796 vdd.n30795 0.005
R66861 vdd.n30877 vdd.n30876 0.005
R66862 vdd.n29572 vdd.n29571 0.005
R66863 vdd.n30795 vdd.n30794 0.005
R66864 vdd.n35023 vdd.n35022 0.004
R66865 vdd.n780 vdd.n779 0.004
R66866 vdd.n5770 vdd.n5769 0.004
R66867 vdd.n4709 vdd.n4708 0.004
R66868 vdd.n4600 vdd.n4599 0.004
R66869 vdd.n779 vdd.n778 0.004
R66870 vdd.n4708 vdd.n4707 0.004
R66871 vdd.n34440 vdd.n34345 0.004
R66872 vdd.n5184 vdd.n5183 0.004
R66873 vdd.n4946 vdd.n4945 0.004
R66874 vdd.n7143 vdd.n7141 0.004
R66875 vdd.n7918 vdd.n7917 0.004
R66876 vdd.n7862 vdd.n7861 0.004
R66877 vdd.n7806 vdd.n7805 0.004
R66878 vdd.n7747 vdd.n7746 0.004
R66879 vdd.n7691 vdd.n7690 0.004
R66880 vdd.n7576 vdd.n7575 0.004
R66881 vdd.n7521 vdd.n7519 0.004
R66882 vdd.n7464 vdd.n7463 0.004
R66883 vdd.n7407 vdd.n7406 0.004
R66884 vdd.n7350 vdd.n7349 0.004
R66885 vdd.n7296 vdd.n7295 0.004
R66886 vdd.n7134 vdd.n7133 0.004
R66887 vdd.n7131 vdd.n7130 0.004
R66888 vdd.n6731 vdd.n6729 0.004
R66889 vdd.n6680 vdd.n6678 0.004
R66890 vdd.n6620 vdd.n6618 0.004
R66891 vdd.n7950 vdd.n7949 0.004
R66892 vdd.n7129 vdd.n7128 0.004
R66893 vdd.n7126 vdd.n7124 0.004
R66894 vdd.n7636 vdd.n7635 0.004
R66895 vdd.n7970 vdd.n7969 0.004
R66896 vdd.n7886 vdd.n7885 0.004
R66897 vdd.n7830 vdd.n7829 0.004
R66898 vdd.n7770 vdd.n7769 0.004
R66899 vdd.n7715 vdd.n7714 0.004
R66900 vdd.n7658 vdd.n7657 0.004
R66901 vdd.n7601 vdd.n7600 0.004
R66902 vdd.n7543 vdd.n7542 0.004
R66903 vdd.n7482 vdd.n7481 0.004
R66904 vdd.n7431 vdd.n7430 0.004
R66905 vdd.n7375 vdd.n7374 0.004
R66906 vdd.n7318 vdd.n7317 0.004
R66907 vdd.n7263 vdd.n7262 0.004
R66908 vdd.n7192 vdd.n7191 0.004
R66909 vdd.n7121 vdd.n7120 0.004
R66910 vdd.n7091 vdd.n7090 0.004
R66911 vdd.n7036 vdd.n7035 0.004
R66912 vdd.n6980 vdd.n6979 0.004
R66913 vdd.n6924 vdd.n6923 0.004
R66914 vdd.n6867 vdd.n6866 0.004
R66915 vdd.n6812 vdd.n6811 0.004
R66916 vdd.n6699 vdd.n6698 0.004
R66917 vdd.n6722 vdd.n6720 0.004
R66918 vdd.n6644 vdd.n6643 0.004
R66919 vdd.n6669 vdd.n6668 0.004
R66920 vdd.n7147 vdd.n7145 0.004
R66921 vdd.n7088 vdd.n7087 0.004
R66922 vdd.n7118 vdd.n7117 0.004
R66923 vdd.n7259 vdd.n7258 0.004
R66924 vdd.n7315 vdd.n7314 0.004
R66925 vdd.n7340 vdd.n7339 0.004
R66926 vdd.n7372 vdd.n7371 0.004
R66927 vdd.n7398 vdd.n7397 0.004
R66928 vdd.n7428 vdd.n7427 0.004
R66929 vdd.n7455 vdd.n7454 0.004
R66930 vdd.n7479 vdd.n7478 0.004
R66931 vdd.n7510 vdd.n7509 0.004
R66932 vdd.n7540 vdd.n7539 0.004
R66933 vdd.n7566 vdd.n7565 0.004
R66934 vdd.n7598 vdd.n7597 0.004
R66935 vdd.n7624 vdd.n7623 0.004
R66936 vdd.n7655 vdd.n7654 0.004
R66937 vdd.n7681 vdd.n7680 0.004
R66938 vdd.n7712 vdd.n7711 0.004
R66939 vdd.n7738 vdd.n7737 0.004
R66940 vdd.n7767 vdd.n7766 0.004
R66941 vdd.n7796 vdd.n7795 0.004
R66942 vdd.n7827 vdd.n7826 0.004
R66943 vdd.n7852 vdd.n7851 0.004
R66944 vdd.n7883 vdd.n7882 0.004
R66945 vdd.n7909 vdd.n7908 0.004
R66946 vdd.n7937 vdd.n7936 0.004
R66947 vdd.n6750 vdd.n6749 0.004
R66948 vdd.n6697 vdd.n6696 0.004
R66949 vdd.n6641 vdd.n6640 0.004
R66950 vdd.n6411 vdd.n6410 0.004
R66951 vdd.n685 vdd.n684 0.004
R66952 vdd.n1163 vdd.n1162 0.004
R66953 vdd.n866 vdd.n865 0.004
R66954 vdd.n29255 vdd.n29254 0.004
R66955 vdd.n31420 vdd.n31419 0.004
R66956 vdd.n30509 vdd.n30508 0.004
R66957 vdd.n25264 vdd.n7978 0.004
R66958 vdd.n32369 vdd.n32368 0.004
R66959 vdd.n387 vdd.n386 0.004
R66960 vdd.n4601 vdd.n4449 0.004
R66961 vdd.n29315 vdd.n29313 0.004
R66962 vdd.n30108 vdd.n30106 0.004
R66963 vdd.n30771 vdd.n30769 0.004
R66964 vdd.n7155 vdd.n7154 0.004
R66965 vdd.n26710 vdd.n26709 0.004
R66966 vdd.n26522 vdd.n26521 0.004
R66967 vdd.n25264 vdd.n7968 0.004
R66968 vdd.n32720 vdd.n32719 0.004
R66969 vdd.n27734 vdd.n27733 0.004
R66970 vdd.n31216 vdd.n31215 0.004
R66971 vdd.n33859 vdd.n33858 0.004
R66972 vdd.n33421 vdd.n33420 0.004
R66973 vdd.n33859 vdd.n33857 0.004
R66974 vdd.n33423 vdd.n33422 0.004
R66975 vdd.n33850 vdd.n33847 0.004
R66976 vdd.n33807 vdd.n33806 0.004
R66977 vdd.n33816 vdd.n33815 0.004
R66978 vdd.n34279 vdd.n34278 0.004
R66979 vdd.n34268 vdd.n34267 0.004
R66980 vdd.n34287 vdd.n34286 0.004
R66981 vdd.n34276 vdd.n34275 0.004
R66982 vdd.n35545 vdd.n35544 0.004
R66983 vdd.n35534 vdd.n35533 0.004
R66984 vdd.n35553 vdd.n35552 0.004
R66985 vdd.n35542 vdd.n35541 0.004
R66986 vdd.n34915 vdd.n34914 0.004
R66987 vdd.n34923 vdd.n34922 0.004
R66988 vdd.n34994 vdd.n34993 0.004
R66989 vdd.n34991 vdd.n34990 0.004
R66990 vdd.n960 vdd.n959 0.004
R66991 vdd.n745 vdd.n744 0.004
R66992 vdd.n960 vdd.n957 0.004
R66993 vdd.n748 vdd.n747 0.004
R66994 vdd.n851 vdd.n848 0.004
R66995 vdd.n814 vdd.n813 0.004
R66996 vdd.n834 vdd.n833 0.004
R66997 vdd.n409 vdd.n408 0.004
R66998 vdd.n404 vdd.n403 0.004
R66999 vdd.n417 vdd.n416 0.004
R67000 vdd.n324 vdd.n323 0.004
R67001 vdd.n5958 vdd.n5957 0.004
R67002 vdd.n5966 vdd.n5965 0.004
R67003 vdd.n6017 vdd.n6016 0.004
R67004 vdd.n6014 vdd.n6013 0.004
R67005 vdd.n5662 vdd.n5661 0.004
R67006 vdd.n5670 vdd.n5669 0.004
R67007 vdd.n5741 vdd.n5740 0.004
R67008 vdd.n5738 vdd.n5737 0.004
R67009 vdd.n4667 vdd.n4666 0.004
R67010 vdd.n4672 vdd.n4671 0.004
R67011 vdd.n4669 vdd.n4668 0.004
R67012 vdd.n4674 vdd.n4673 0.004
R67013 vdd.n4950 vdd.n4949 0.004
R67014 vdd.n4489 vdd.n4488 0.004
R67015 vdd.n4497 vdd.n4496 0.004
R67016 vdd.n4571 vdd.n4570 0.004
R67017 vdd.n4568 vdd.n4567 0.004
R67018 vdd.n37042 vdd.n37030 0.004
R67019 vdd.n33285 vdd.n33284 0.004
R67020 vdd.n37076 vdd.n37064 0.004
R67021 vdd.n33203 vdd.n33188 0.004
R67022 vdd.n37132 vdd.n37131 0.004
R67023 vdd.n33162 vdd.n33150 0.004
R67024 vdd.n37208 vdd.n37193 0.004
R67025 vdd.n33116 vdd.n33115 0.004
R67026 vdd.n37296 vdd.n37295 0.004
R67027 vdd.n35654 vdd.n35650 0.004
R67028 vdd.n32944 vdd.n32943 0.004
R67029 vdd.n37473 vdd.n37460 0.004
R67030 vdd.n32836 vdd.n32822 0.004
R67031 vdd.n37574 vdd.n37573 0.004
R67032 vdd.n29749 vdd.n29747 0.004
R67033 vdd.n29952 vdd.n29951 0.004
R67034 vdd.n29828 vdd.n29825 0.004
R67035 vdd.n27802 vdd.n27798 0.004
R67036 vdd.n28971 vdd.n28969 0.004
R67037 vdd.n28804 vdd.n28803 0.004
R67038 vdd.n28838 vdd.n28818 0.004
R67039 vdd.n28818 vdd.n28817 0.004
R67040 vdd.n28864 vdd.n28861 0.004
R67041 vdd.n28900 vdd.n28897 0.004
R67042 vdd.n28958 vdd.n28953 0.004
R67043 vdd.n28048 vdd.n28046 0.004
R67044 vdd.n28001 vdd.n27999 0.004
R67045 vdd.n27964 vdd.n27961 0.004
R67046 vdd.n29916 vdd.n29911 0.004
R67047 vdd.n29918 vdd.n29917 0.004
R67048 vdd.n29943 vdd.n29942 0.004
R67049 vdd.n29793 vdd.n29790 0.004
R67050 vdd.n29729 vdd.n29727 0.004
R67051 vdd.n30652 vdd.n30649 0.004
R67052 vdd.n30608 vdd.n30606 0.004
R67053 vdd.n30581 vdd.n30580 0.004
R67054 vdd.n30576 vdd.n30575 0.004
R67055 vdd.n30538 vdd.n30536 0.004
R67056 vdd.n32812 vdd.n6406 0.004
R67057 vdd.n32804 vdd.n6489 0.004
R67058 vdd.n32799 vdd.n6547 0.004
R67059 vdd.n32788 vdd.n6660 0.004
R67060 vdd.n32778 vdd.n6771 0.004
R67061 vdd.n32772 vdd.n6830 0.004
R67062 vdd.n32766 vdd.n6885 0.004
R67063 vdd.n32760 vdd.n6942 0.004
R67064 vdd.n32754 vdd.n6999 0.004
R67065 vdd.n32748 vdd.n7055 0.004
R67066 vdd.n32737 vdd.n7221 0.004
R67067 vdd.n32802 vdd.n6513 0.004
R67068 vdd.n32796 vdd.n6570 0.004
R67069 vdd.n32790 vdd.n6627 0.004
R67070 vdd.n32775 vdd.n6797 0.004
R67071 vdd.n32769 vdd.n6852 0.004
R67072 vdd.n32763 vdd.n6908 0.004
R67073 vdd.n32757 vdd.n6965 0.004
R67074 vdd.n32751 vdd.n7021 0.004
R67075 vdd.n32745 vdd.n7075 0.004
R67076 vdd.n30901 vdd.n30900 0.004
R67077 vdd.n32547 vdd.n32546 0.004
R67078 vdd.n29597 vdd.n29596 0.004
R67079 vdd.n29448 vdd.n29447 0.004
R67080 vdd.n29421 vdd.n29420 0.004
R67081 vdd.n27690 vdd.n27689 0.004
R67082 vdd.n26460 vdd.n26459 0.004
R67083 vdd.n26364 vdd.n26363 0.004
R67084 vdd.n26275 vdd.n26274 0.004
R67085 vdd.n30994 vdd.n30993 0.004
R67086 vdd.n26472 vdd.n26453 0.004
R67087 vdd.n29530 vdd.n29520 0.004
R67088 vdd.n30813 vdd.n30786 0.004
R67089 vdd.n31319 vdd.n31316 0.004
R67090 vdd.n27660 vdd.n27252 0.004
R67091 vdd.n35615 vdd.n35614 0.004
R67092 vdd.n35029 vdd.n35028 0.004
R67093 vdd.n6363 vdd.n1175 0.004
R67094 vdd.n6361 vdd.n6360 0.004
R67095 vdd.n3681 vdd.n3680 0.004
R67096 vdd.n3692 vdd.n3687 0.004
R67097 vdd.n3706 vdd.n3703 0.004
R67098 vdd.n3711 vdd.n3706 0.004
R67099 vdd.n4002 vdd.n4000 0.004
R67100 vdd.n3987 vdd.n3985 0.004
R67101 vdd.n3983 vdd.n3982 0.004
R67102 vdd.n3977 vdd.n3974 0.004
R67103 vdd.n3972 vdd.n3970 0.004
R67104 vdd.n3961 vdd.n3959 0.004
R67105 vdd.n3944 vdd.n3943 0.004
R67106 vdd.n3942 vdd.n3940 0.004
R67107 vdd.n3929 vdd.n3926 0.004
R67108 vdd.n3926 vdd.n3924 0.004
R67109 vdd.n3914 vdd.n3909 0.004
R67110 vdd.n3909 vdd.n3906 0.004
R67111 vdd.n3892 vdd.n3891 0.004
R67112 vdd.n3865 vdd.n3864 0.004
R67113 vdd.n3846 vdd.n3845 0.004
R67114 vdd.n3843 vdd.n3841 0.004
R67115 vdd.n2222 vdd.n2220 0.004
R67116 vdd.n2228 vdd.n2225 0.004
R67117 vdd.n2248 vdd.n2247 0.004
R67118 vdd.n2258 vdd.n2257 0.004
R67119 vdd.n2265 vdd.n2264 0.004
R67120 vdd.n2279 vdd.n2276 0.004
R67121 vdd.n2284 vdd.n2279 0.004
R67122 vdd.n2315 vdd.n2314 0.004
R67123 vdd.n2334 vdd.n2333 0.004
R67124 vdd.n2341 vdd.n2336 0.004
R67125 vdd.n2349 vdd.n2346 0.004
R67126 vdd.n2353 vdd.n2352 0.004
R67127 vdd.n2368 vdd.n2367 0.004
R67128 vdd.n2559 vdd.n2558 0.004
R67129 vdd.n2554 vdd.n2553 0.004
R67130 vdd.n2553 vdd.n2550 0.004
R67131 vdd.n2539 vdd.n2536 0.004
R67132 vdd.n2516 vdd.n2514 0.004
R67133 vdd.n2472 vdd.n2471 0.004
R67134 vdd.n2469 vdd.n2467 0.004
R67135 vdd.n2605 vdd.n2603 0.004
R67136 vdd.n2611 vdd.n2608 0.004
R67137 vdd.n2631 vdd.n2630 0.004
R67138 vdd.n2658 vdd.n2656 0.004
R67139 vdd.n2665 vdd.n2664 0.004
R67140 vdd.n1973 vdd.n1970 0.004
R67141 vdd.n1980 vdd.n1973 0.004
R67142 vdd.n1995 vdd.n1993 0.004
R67143 vdd.n2096 vdd.n2095 0.004
R67144 vdd.n1957 vdd.n1955 0.004
R67145 vdd.n1951 vdd.n1950 0.004
R67146 vdd.n1949 vdd.n1946 0.004
R67147 vdd.n1882 vdd.n1873 0.004
R67148 vdd.n1873 vdd.n1872 0.004
R67149 vdd.n1856 vdd.n1854 0.004
R67150 vdd.n1851 vdd.n1848 0.004
R67151 vdd.n1791 vdd.n1790 0.004
R67152 vdd.n1788 vdd.n1786 0.004
R67153 vdd.n26199 vdd.n26198 0.004
R67154 vdd.n26598 vdd.n26595 0.004
R67155 vdd.n31760 vdd.n31759 0.004
R67156 vdd.n31811 vdd.n31808 0.004
R67157 vdd.n31819 vdd.n31814 0.004
R67158 vdd.n31825 vdd.n31824 0.004
R67159 vdd.n31830 vdd.n31827 0.004
R67160 vdd.n31855 vdd.n31852 0.004
R67161 vdd.n31875 vdd.n31872 0.004
R67162 vdd.n31915 vdd.n31912 0.004
R67163 vdd.n31939 vdd.n31938 0.004
R67164 vdd.n31979 vdd.n31978 0.004
R67165 vdd.n31991 vdd.n31988 0.004
R67166 vdd.n32141 vdd.n32138 0.004
R67167 vdd.n32169 vdd.n32166 0.004
R67168 vdd.n32177 vdd.n32172 0.004
R67169 vdd.n32186 vdd.n32185 0.004
R67170 vdd.n32191 vdd.n32188 0.004
R67171 vdd.n32213 vdd.n32210 0.004
R67172 vdd.n32300 vdd.n32298 0.004
R67173 vdd.n32337 vdd.n32336 0.004
R67174 vdd.n32351 vdd.n32348 0.004
R67175 vdd.n32478 vdd.n32476 0.004
R67176 vdd.n32474 vdd.n32473 0.004
R67177 vdd.n32463 vdd.n32461 0.004
R67178 vdd.n31055 vdd.n31052 0.004
R67179 vdd.n31063 vdd.n31058 0.004
R67180 vdd.n31072 vdd.n31071 0.004
R67181 vdd.n31078 vdd.n31075 0.004
R67182 vdd.n31107 vdd.n31104 0.004
R67183 vdd.n29282 vdd.n29281 0.004
R67184 vdd.n29297 vdd.n29296 0.004
R67185 vdd.n29464 vdd.n29438 0.004
R67186 vdd.n29530 vdd.n29517 0.004
R67187 vdd.n32666 vdd.n32665 0.004
R67188 vdd.n29642 vdd.n29641 0.004
R67189 vdd.n29646 vdd.n29645 0.004
R67190 vdd.n30059 vdd.n30044 0.004
R67191 vdd.n30090 vdd.n30089 0.004
R67192 vdd.n30813 vdd.n30779 0.004
R67193 vdd.n30743 vdd.n30742 0.004
R67194 vdd.n31237 vdd.n31236 0.004
R67195 vdd.n31249 vdd.n31248 0.004
R67196 vdd.n30776 vdd.n30773 0.004
R67197 vdd.n26217 vdd.n26216 0.004
R67198 vdd.n26672 vdd.n26671 0.004
R67199 vdd.n26407 vdd.n26406 0.004
R67200 vdd.n26472 vdd.n26471 0.004
R67201 vdd.n29095 vdd.n29094 0.004
R67202 vdd.n10541 vdd.n10540 0.004
R67203 vdd.n12437 vdd.n12436 0.004
R67204 vdd.n12420 vdd.n12419 0.004
R67205 vdd.n10839 vdd.n10838 0.004
R67206 vdd.n10880 vdd.n10879 0.004
R67207 vdd.n11023 vdd.n10997 0.004
R67208 vdd.n12217 vdd.n11034 0.004
R67209 vdd.n12139 vdd.n12138 0.004
R67210 vdd.n11216 vdd.n11197 0.004
R67211 vdd.n11348 vdd.n11347 0.004
R67212 vdd.n11389 vdd.n11388 0.004
R67213 vdd.n11487 vdd.n11470 0.004
R67214 vdd.n11521 vdd.n11520 0.004
R67215 vdd.n13947 vdd.n8636 0.004
R67216 vdd.n14017 vdd.n14016 0.004
R67217 vdd.n14237 vdd.n8414 0.004
R67218 vdd.n14306 vdd.n8361 0.004
R67219 vdd.n14554 vdd.n14553 0.004
R67220 vdd.n9258 vdd.n9257 0.004
R67221 vdd.n9082 vdd.n9081 0.004
R67222 vdd.n9027 vdd.n9013 0.004
R67223 vdd.n8862 vdd.n8861 0.004
R67224 vdd.n8807 vdd.n8793 0.004
R67225 vdd.n10400 vdd.n10331 0.004
R67226 vdd.n10364 vdd.n10363 0.004
R67227 vdd.n13007 vdd.n13006 0.004
R67228 vdd.n12968 vdd.n9451 0.004
R67229 vdd.n9588 vdd.n9576 0.004
R67230 vdd.n9654 vdd.n9627 0.004
R67231 vdd.n12799 vdd.n12798 0.004
R67232 vdd.n12760 vdd.n9810 0.004
R67233 vdd.n9948 vdd.n9935 0.004
R67234 vdd.n10014 vdd.n9987 0.004
R67235 vdd.n11755 vdd.n11718 0.004
R67236 vdd.n11706 vdd.n11703 0.004
R67237 vdd.n11862 vdd.n11812 0.004
R67238 vdd.n11849 vdd.n11842 0.004
R67239 vdd.n13182 vdd.n9219 0.004
R67240 vdd.n9207 vdd.n9205 0.004
R67241 vdd.n9176 vdd.n9162 0.004
R67242 vdd.n13273 vdd.n13272 0.004
R67243 vdd.n14350 vdd.n8339 0.004
R67244 vdd.n14353 vdd.n14352 0.004
R67245 vdd.n14424 vdd.n14423 0.004
R67246 vdd.n14458 vdd.n8246 0.004
R67247 vdd.n14651 vdd.n14650 0.004
R67248 vdd.n14691 vdd.n14690 0.004
R67249 vdd.n14720 vdd.n14719 0.004
R67250 vdd.n14765 vdd.n8091 0.004
R67251 vdd.n14768 vdd.n14767 0.004
R67252 vdd.n14807 vdd.n8060 0.004
R67253 vdd.n14823 vdd.n14822 0.004
R67254 vdd.n14865 vdd.n14864 0.004
R67255 vdd.n14900 vdd.n14899 0.004
R67256 vdd.n14937 vdd.n14936 0.004
R67257 vdd.n22341 vdd.n22255 0.004
R67258 vdd.n22340 vdd.n22339 0.004
R67259 vdd.n24304 vdd.n22131 0.004
R67260 vdd.n24303 vdd.n22141 0.004
R67261 vdd.n22292 vdd.n22280 0.004
R67262 vdd.n24352 vdd.n24351 0.004
R67263 vdd.n24264 vdd.n24252 0.004
R67264 vdd.n24235 vdd.n24234 0.004
R67265 vdd.n24188 vdd.n24178 0.004
R67266 vdd.n23996 vdd.n23994 0.004
R67267 vdd.n23956 vdd.n23946 0.004
R67268 vdd.n23764 vdd.n23762 0.004
R67269 vdd.n23724 vdd.n23714 0.004
R67270 vdd.n23076 vdd.n23074 0.004
R67271 vdd.n23268 vdd.n23258 0.004
R67272 vdd.n23308 vdd.n23306 0.004
R67273 vdd.n23500 vdd.n23490 0.004
R67274 vdd.n23540 vdd.n23538 0.004
R67275 vdd.n22497 vdd.n22495 0.004
R67276 vdd.n22689 vdd.n22679 0.004
R67277 vdd.n22729 vdd.n22727 0.004
R67278 vdd.n22921 vdd.n22911 0.004
R67279 vdd.n22961 vdd.n22959 0.004
R67280 vdd.n22436 vdd.n22424 0.004
R67281 vdd.n22407 vdd.n22406 0.004
R67282 vdd.n16887 vdd.n16873 0.004
R67283 vdd.n17093 vdd.n17092 0.004
R67284 vdd.n17159 vdd.n17145 0.004
R67285 vdd.n17365 vdd.n17364 0.004
R67286 vdd.n17431 vdd.n17417 0.004
R67287 vdd.n17623 vdd.n17622 0.004
R67288 vdd.n17689 vdd.n17675 0.004
R67289 vdd.n17894 vdd.n17893 0.004
R67290 vdd.n17960 vdd.n17946 0.004
R67291 vdd.n18166 vdd.n18165 0.004
R67292 vdd.n18231 vdd.n18218 0.004
R67293 vdd.n18309 vdd.n18308 0.004
R67294 vdd.n18350 vdd.n18349 0.004
R67295 vdd.n19055 vdd.n19053 0.004
R67296 vdd.n18990 vdd.n18988 0.004
R67297 vdd.n18796 vdd.n18794 0.004
R67298 vdd.n18731 vdd.n18729 0.004
R67299 vdd.n18537 vdd.n18535 0.004
R67300 vdd.n21624 vdd.n21623 0.004
R67301 vdd.n21421 vdd.n21419 0.004
R67302 vdd.n21356 vdd.n21354 0.004
R67303 vdd.n21162 vdd.n21160 0.004
R67304 vdd.n21097 vdd.n21095 0.004
R67305 vdd.n15400 vdd.n15399 0.004
R67306 vdd.n15446 vdd.n15434 0.004
R67307 vdd.n15648 vdd.n15647 0.004
R67308 vdd.n15702 vdd.n15687 0.004
R67309 vdd.n15904 vdd.n15903 0.004
R67310 vdd.n15958 vdd.n15943 0.004
R67311 vdd.n16160 vdd.n16159 0.004
R67312 vdd.n16214 vdd.n16199 0.004
R67313 vdd.n16416 vdd.n16415 0.004
R67314 vdd.n16470 vdd.n16455 0.004
R67315 vdd.n20676 vdd.n20664 0.004
R67316 vdd.n20660 vdd.n20648 0.004
R67317 vdd.n20613 vdd.n20611 0.004
R67318 vdd.n20597 vdd.n20595 0.004
R67319 vdd.n20466 vdd.n20465 0.004
R67320 vdd.n20423 vdd.n20411 0.004
R67321 vdd.n20367 vdd.n20365 0.004
R67322 vdd.n20305 vdd.n20303 0.004
R67323 vdd.n20289 vdd.n20287 0.004
R67324 vdd.n20255 vdd.n20253 0.004
R67325 vdd.n20239 vdd.n20237 0.004
R67326 vdd.n20187 vdd.n20175 0.004
R67327 vdd.n20131 vdd.n20129 0.004
R67328 vdd.n20069 vdd.n20067 0.004
R67329 vdd.n19388 vdd.n19386 0.004
R67330 vdd.n19404 vdd.n19402 0.004
R67331 vdd.n19451 vdd.n19439 0.004
R67332 vdd.n19467 vdd.n19455 0.004
R67333 vdd.n21770 vdd.n21769 0.004
R67334 vdd.n21778 vdd.n21776 0.004
R67335 vdd.n21953 vdd.n21903 0.004
R67336 vdd.n21940 vdd.n21933 0.004
R67337 vdd.n24974 vdd.n24973 0.004
R67338 vdd.n25052 vdd.n25051 0.004
R67339 vdd.n24937 vdd.n24936 0.004
R67340 vdd.n24948 vdd.n24947 0.004
R67341 vdd.n24560 vdd.n24559 0.004
R67342 vdd.n24632 vdd.n24631 0.004
R67343 vdd.n24685 vdd.n24683 0.004
R67344 vdd.n24697 vdd.n24695 0.004
R67345 vdd.n24719 vdd.n24717 0.004
R67346 vdd.n24782 vdd.n24774 0.004
R67347 vdd.n24798 vdd.n24796 0.004
R67348 vdd.n24810 vdd.n24808 0.004
R67349 vdd.n25228 vdd.n25226 0.004
R67350 vdd.n25216 vdd.n25214 0.004
R67351 vdd.n25200 vdd.n25192 0.004
R67352 vdd.n25148 vdd.n25140 0.004
R67353 vdd.n25137 vdd.n25135 0.004
R67354 vdd.n25115 vdd.n25113 0.004
R67355 vdd.n25103 vdd.n25101 0.004
R67356 vdd.n35231 vdd.n35230 0.004
R67357 vdd.n34644 vdd.n34643 0.004
R67358 vdd.n5391 vdd.n5390 0.004
R67359 vdd.n4221 vdd.n4220 0.004
R67360 vdd.n35230 vdd.n35229 0.004
R67361 vdd.n34643 vdd.n34642 0.004
R67362 vdd.n5390 vdd.n5389 0.004
R67363 vdd.n4220 vdd.n4219 0.004
R67364 vdd.n29573 vdd.n29572 0.004
R67365 vdd.n30878 vdd.n30877 0.004
R67366 vdd.n30897 vdd.n30896 0.004
R67367 vdd.n29594 vdd.n29593 0.004
R67368 vdd.n27687 vdd.n27686 0.004
R67369 vdd.n31959 vdd.n31955 0.004
R67370 vdd.n35617 vdd.n34443 0.004
R67371 vdd.n5776 vdd.n5775 0.004
R67372 vdd.n5190 vdd.n5189 0.004
R67373 vdd.n4606 vdd.n4605 0.004
R67374 vdd.n35619 vdd.n33863 0.004
R67375 vdd.n4222 vdd.n4221 0.004
R67376 vdd.n4599 vdd.n4598 0.004
R67377 vdd.n4343 vdd.n4342 0.004
R67378 vdd.n4710 vdd.n4709 0.004
R67379 vdd.n5392 vdd.n5391 0.004
R67380 vdd.n5769 vdd.n5768 0.004
R67381 vdd.n5516 vdd.n5515 0.004
R67382 vdd.n34645 vdd.n34644 0.004
R67383 vdd.n35022 vdd.n35021 0.004
R67384 vdd.n34769 vdd.n34768 0.004
R67385 vdd.n35232 vdd.n35231 0.004
R67386 vdd.n35610 vdd.n35609 0.004
R67387 vdd.n35353 vdd.n35352 0.004
R67388 vdd.n1167 vdd.n1166 0.004
R67389 vdd.n882 vdd.n873 0.004
R67390 vdd.n4602 vdd.n4601 0.004
R67391 vdd.n35025 vdd.n35024 0.004
R67392 vdd.n5772 vdd.n5771 0.004
R67393 vdd.n28803 vdd.n28802 0.004
R67394 vdd.n31212 vdd.n31211 0.004
R67395 vdd.n33856 vdd.n33855 0.004
R67396 vdd.n956 vdd.n955 0.004
R67397 vdd.n30956 vdd.n30955 0.004
R67398 vdd.n467 vdd.n466 0.004
R67399 vdd.n185 vdd.n184 0.004
R67400 vdd.n380 vdd.n379 0.004
R67401 vdd.n33453 vdd.n33452 0.004
R67402 vdd.n30739 vdd.n30738 0.004
R67403 vdd.n32603 vdd.n32602 0.004
R67404 vdd.n29378 vdd.n29377 0.004
R67405 vdd.n26239 vdd.n26238 0.004
R67406 vdd.n24970 vdd.n24969 0.004
R67407 vdd.n25643 vdd.n25422 0.004
R67408 vdd.n7140 vdd.n7138 0.004
R67409 vdd.n6406 vdd.n6405 0.004
R67410 vdd.n6468 vdd.n6466 0.004
R67411 vdd.n6636 vdd.n6635 0.004
R67412 vdd.n6746 vdd.n6744 0.004
R67413 vdd.n7151 vdd.n7150 0.004
R67414 vdd.n7312 vdd.n7311 0.004
R67415 vdd.n7368 vdd.n7367 0.004
R67416 vdd.n7424 vdd.n7422 0.004
R67417 vdd.n7475 vdd.n7474 0.004
R67418 vdd.n7536 vdd.n7535 0.004
R67419 vdd.n7594 vdd.n7592 0.004
R67420 vdd.n7651 vdd.n7649 0.004
R67421 vdd.n7708 vdd.n7706 0.004
R67422 vdd.n7763 vdd.n7761 0.004
R67423 vdd.n7822 vdd.n7821 0.004
R67424 vdd.n7879 vdd.n7878 0.004
R67425 vdd.n7933 vdd.n7932 0.004
R67426 vdd.n6390 vdd.n6389 0.004
R67427 vdd.n6429 vdd.n6428 0.004
R67428 vdd.n6655 vdd.n6653 0.004
R67429 vdd.n6710 vdd.n6709 0.004
R67430 vdd.n7107 vdd.n7105 0.004
R67431 vdd.n7209 vdd.n7208 0.004
R67432 vdd.n7276 vdd.n7274 0.004
R67433 vdd.n7330 vdd.n7329 0.004
R67434 vdd.n7387 vdd.n7385 0.004
R67435 vdd.n7444 vdd.n7442 0.004
R67436 vdd.n7497 vdd.n7495 0.004
R67437 vdd.n7555 vdd.n7554 0.004
R67438 vdd.n7613 vdd.n7611 0.004
R67439 vdd.n7670 vdd.n7668 0.004
R67440 vdd.n7727 vdd.n7725 0.004
R67441 vdd.n7784 vdd.n7782 0.004
R67442 vdd.n7841 vdd.n7840 0.004
R67443 vdd.n7898 vdd.n7896 0.004
R67444 vdd.n7974 vdd.n7973 0.004
R67445 vdd.n4347 vdd.n4346 0.004
R67446 vdd.n5520 vdd.n5519 0.004
R67447 vdd.n34773 vdd.n34772 0.004
R67448 vdd.n35357 vdd.n35356 0.004
R67449 vdd.n10246 vdd.n10235 0.004
R67450 vdd.n16669 vdd.n16648 0.004
R67451 vdd.n5185 vdd.n5184 0.004
R67452 vdd.n4947 vdd.n4946 0.004
R67453 vdd.n781 vdd.n780 0.004
R67454 vdd.n6040 vdd.n6039 0.004
R67455 vdd.n5923 vdd.n5922 0.004
R67456 vdd.n34062 vdd.n34061 0.004
R67457 vdd.n24838 vdd.n24837 0.004
R67458 vdd.n686 vdd.n685 0.003
R67459 vdd.n1164 vdd.n1163 0.003
R67460 vdd.n865 vdd.n864 0.003
R67461 vdd.n5178 vdd.n5177 0.003
R67462 vdd.n4936 vdd.n4935 0.003
R67463 vdd.n6137 vdd.n6136 0.003
R67464 vdd.n26510 vdd.n26509 0.003
R67465 vdd.n4606 vdd.n4021 0.003
R67466 vdd.n35620 vdd.n35619 0.003
R67467 vdd.n34157 vdd.n34156 0.003
R67468 vdd.n30775 vdd.n30774 0.003
R67469 vdd.n5848 vdd.n5847 0.003
R67470 vdd.n11918 vdd.n11917 0.003
R67471 vdd.n22004 vdd.n22003 0.003
R67472 vdd.n10246 vdd.n10228 0.003
R67473 vdd.n16669 vdd.n16605 0.003
R67474 vdd.n30943 vdd.n30942 0.003
R67475 vdd.n2637 vdd.n2632 0.003
R67476 vdd.n32814 vdd.n32812 0.003
R67477 vdd.n31188 vdd.n31187 0.003
R67478 vdd.n25264 vdd.n7965 0.003
R67479 vdd.n26135 vdd.n26134 0.003
R67480 vdd.n33780 vdd.n33779 0.003
R67481 vdd.n26155 vdd.n26151 0.003
R67482 vdd.n4214 vdd.n4213 0.003
R67483 vdd.n5384 vdd.n5383 0.003
R67484 vdd.n1168 vdd.n1167 0.003
R67485 vdd.n882 vdd.n881 0.003
R67486 vdd.n34637 vdd.n34636 0.003
R67487 vdd.n35224 vdd.n35223 0.003
R67488 vdd.n30783 vdd.n30782 0.003
R67489 vdd.n30970 vdd.n30969 0.003
R67490 vdd.n30762 vdd.n30761 0.003
R67491 vdd.n31785 vdd.n31782 0.003
R67492 vdd.n32077 vdd.n32076 0.003
R67493 vdd.n32388 vdd.n32383 0.003
R67494 vdd.n33447 vdd.n33445 0.003
R67495 vdd.n33372 vdd.n33371 0.003
R67496 vdd.n33485 vdd.n33484 0.003
R67497 vdd.n33334 vdd.n33332 0.003
R67498 vdd.n33356 vdd.n33353 0.003
R67499 vdd.n33768 vdd.n33718 0.003
R67500 vdd.n33720 vdd.n33719 0.003
R67501 vdd.n33730 vdd.n33729 0.003
R67502 vdd.n33572 vdd.n33571 0.003
R67503 vdd.n33684 vdd.n33681 0.003
R67504 vdd.n33680 vdd.n33677 0.003
R67505 vdd.n33787 vdd.n33783 0.003
R67506 vdd.n33794 vdd.n33791 0.003
R67507 vdd.n33847 vdd.n33846 0.003
R67508 vdd.n33799 vdd.n33798 0.003
R67509 vdd.n34155 vdd.n34083 0.003
R67510 vdd.n34112 vdd.n34109 0.003
R67511 vdd.n34333 vdd.n34331 0.003
R67512 vdd.n34219 vdd.n34216 0.003
R67513 vdd.n34215 vdd.n34213 0.003
R67514 vdd.n34428 vdd.n34427 0.003
R67515 vdd.n34359 vdd.n34358 0.003
R67516 vdd.n33919 vdd.n33917 0.003
R67517 vdd.n33880 vdd.n33878 0.003
R67518 vdd.n33956 vdd.n33953 0.003
R67519 vdd.n33885 vdd.n33884 0.003
R67520 vdd.n35498 vdd.n35497 0.003
R67521 vdd.n35275 vdd.n35242 0.003
R67522 vdd.n35599 vdd.n35597 0.003
R67523 vdd.n35110 vdd.n35109 0.003
R67524 vdd.n35105 vdd.n35103 0.003
R67525 vdd.n35042 vdd.n35039 0.003
R67526 vdd.n35065 vdd.n35063 0.003
R67527 vdd.n35386 vdd.n35385 0.003
R67528 vdd.n35375 vdd.n35374 0.003
R67529 vdd.n35339 vdd.n35336 0.003
R67530 vdd.n35335 vdd.n35333 0.003
R67531 vdd.n34691 vdd.n34655 0.003
R67532 vdd.n34946 vdd.n34945 0.003
R67533 vdd.n35011 vdd.n35009 0.003
R67534 vdd.n34755 vdd.n34752 0.003
R67535 vdd.n34751 vdd.n34749 0.003
R67536 vdd.n34858 vdd.n34857 0.003
R67537 vdd.n34785 vdd.n34784 0.003
R67538 vdd.n34478 vdd.n34476 0.003
R67539 vdd.n34518 vdd.n34516 0.003
R67540 vdd.n34458 vdd.n34455 0.003
R67541 vdd.n34523 vdd.n34522 0.003
R67542 vdd.n766 vdd.n764 0.003
R67543 vdd.n594 vdd.n593 0.003
R67544 vdd.n972 vdd.n971 0.003
R67545 vdd.n623 vdd.n621 0.003
R67546 vdd.n674 vdd.n671 0.003
R67547 vdd.n911 vdd.n910 0.003
R67548 vdd.n884 vdd.n883 0.003
R67549 vdd.n939 vdd.n938 0.003
R67550 vdd.n1171 vdd.n1170 0.003
R67551 vdd.n1149 vdd.n1146 0.003
R67552 vdd.n1145 vdd.n1142 0.003
R67553 vdd.n863 vdd.n859 0.003
R67554 vdd.n858 vdd.n856 0.003
R67555 vdd.n848 vdd.n847 0.003
R67556 vdd.n830 vdd.n829 0.003
R67557 vdd.n525 vdd.n523 0.003
R67558 vdd.n566 vdd.n563 0.003
R67559 vdd.n582 vdd.n581 0.003
R67560 vdd.n503 vdd.n493 0.003
R67561 vdd.n25 vdd.n24 0.003
R67562 vdd.n30 vdd.n27 0.003
R67563 vdd.n36 vdd.n33 0.003
R67564 vdd.n20 vdd.n18 0.003
R67565 vdd.n54 vdd.n52 0.003
R67566 vdd.n396 vdd.n394 0.003
R67567 vdd.n461 vdd.n459 0.003
R67568 vdd.n263 vdd.n262 0.003
R67569 vdd.n271 vdd.n266 0.003
R67570 vdd.n110 vdd.n109 0.003
R67571 vdd.n179 vdd.n176 0.003
R67572 vdd.n377 vdd.n374 0.003
R67573 vdd.n373 vdd.n371 0.003
R67574 vdd.n5999 vdd.n5998 0.003
R67575 vdd.n5841 vdd.n5785 0.003
R67576 vdd.n6034 vdd.n6032 0.003
R67577 vdd.n6159 vdd.n6158 0.003
R67578 vdd.n6154 vdd.n6152 0.003
R67579 vdd.n6240 vdd.n6237 0.003
R67580 vdd.n6193 vdd.n6191 0.003
R67581 vdd.n6079 vdd.n6078 0.003
R67582 vdd.n6065 vdd.n6064 0.003
R67583 vdd.n5920 vdd.n5917 0.003
R67584 vdd.n5916 vdd.n5914 0.003
R67585 vdd.n5438 vdd.n5402 0.003
R67586 vdd.n5693 vdd.n5692 0.003
R67587 vdd.n5758 vdd.n5756 0.003
R67588 vdd.n5502 vdd.n5499 0.003
R67589 vdd.n5498 vdd.n5496 0.003
R67590 vdd.n5605 vdd.n5604 0.003
R67591 vdd.n5532 vdd.n5531 0.003
R67592 vdd.n5225 vdd.n5223 0.003
R67593 vdd.n5265 vdd.n5263 0.003
R67594 vdd.n5205 vdd.n5202 0.003
R67595 vdd.n5270 vdd.n5269 0.003
R67596 vdd.n5094 vdd.n5092 0.003
R67597 vdd.n4843 vdd.n4838 0.003
R67598 vdd.n4834 vdd.n4833 0.003
R67599 vdd.n4819 vdd.n4818 0.003
R67600 vdd.n4778 vdd.n4777 0.003
R67601 vdd.n4720 vdd.n4719 0.003
R67602 vdd.n4996 vdd.n4994 0.003
R67603 vdd.n5046 vdd.n5043 0.003
R67604 vdd.n4963 vdd.n4961 0.003
R67605 vdd.n4968 vdd.n4967 0.003
R67606 vdd.n4711 vdd.n4616 0.003
R67607 vdd.n4698 vdd.n4696 0.003
R67608 vdd.n4929 vdd.n4927 0.003
R67609 vdd.n4265 vdd.n4232 0.003
R67610 vdd.n4520 vdd.n4519 0.003
R67611 vdd.n4588 vdd.n4586 0.003
R67612 vdd.n4329 vdd.n4326 0.003
R67613 vdd.n4325 vdd.n4323 0.003
R67614 vdd.n4432 vdd.n4431 0.003
R67615 vdd.n4359 vdd.n4358 0.003
R67616 vdd.n4055 vdd.n4053 0.003
R67617 vdd.n4095 vdd.n4093 0.003
R67618 vdd.n4035 vdd.n4032 0.003
R67619 vdd.n4100 vdd.n4099 0.003
R67620 vdd.n2099 vdd.n2098 0.003
R67621 vdd.n36975 vdd.n36973 0.003
R67622 vdd.n36989 vdd.n36987 0.003
R67623 vdd.n37015 vdd.n37014 0.003
R67624 vdd.n37030 vdd.n37029 0.003
R67625 vdd.n33285 vdd.n33275 0.003
R67626 vdd.n37061 vdd.n37059 0.003
R67627 vdd.n33272 vdd.n33271 0.003
R67628 vdd.n33271 vdd.n33269 0.003
R67629 vdd.n37127 vdd.n37126 0.003
R67630 vdd.n33184 vdd.n33181 0.003
R67631 vdd.n37153 vdd.n37140 0.003
R67632 vdd.n37140 vdd.n37137 0.003
R67633 vdd.n37188 vdd.n37187 0.003
R67634 vdd.n37208 vdd.n37207 0.003
R67635 vdd.n33106 vdd.n33105 0.003
R67636 vdd.n33099 vdd.n33093 0.003
R67637 vdd.n37230 vdd.n37229 0.003
R67638 vdd.n37239 vdd.n37230 0.003
R67639 vdd.n37238 vdd.n37235 0.003
R67640 vdd.n33076 vdd.n33075 0.003
R67641 vdd.n33088 vdd.n33087 0.003
R67642 vdd.n37262 vdd.n37261 0.003
R67643 vdd.n33064 vdd.n33060 0.003
R67644 vdd.n33041 vdd.n33029 0.003
R67645 vdd.n33041 vdd.n33040 0.003
R67646 vdd.n37293 vdd.n37292 0.003
R67647 vdd.n33023 vdd.n33019 0.003
R67648 vdd.n37315 vdd.n37303 0.003
R67649 vdd.n32995 vdd.n32994 0.003
R67650 vdd.n33004 vdd.n32995 0.003
R67651 vdd.n33003 vdd.n33001 0.003
R67652 vdd.n37328 vdd.n37327 0.003
R67653 vdd.n37340 vdd.n37339 0.003
R67654 vdd.n37364 vdd.n37363 0.003
R67655 vdd.n32981 vdd.n32980 0.003
R67656 vdd.n37390 vdd.n37375 0.003
R67657 vdd.n37390 vdd.n37389 0.003
R67658 vdd.n32952 vdd.n32951 0.003
R67659 vdd.n37411 vdd.n37398 0.003
R67660 vdd.n37433 vdd.n37425 0.003
R67661 vdd.n37432 vdd.n37429 0.003
R67662 vdd.n32931 vdd.n32930 0.003
R67663 vdd.n32937 vdd.n32936 0.003
R67664 vdd.n37447 vdd.n37436 0.003
R67665 vdd.n37457 vdd.n37447 0.003
R67666 vdd.n32919 vdd.n32915 0.003
R67667 vdd.n37472 vdd.n37471 0.003
R67668 vdd.n32894 vdd.n32889 0.003
R67669 vdd.n32894 vdd.n32893 0.003
R67670 vdd.n32878 vdd.n32874 0.003
R67671 vdd.n37516 vdd.n37515 0.003
R67672 vdd.n32859 vdd.n32850 0.003
R67673 vdd.n32858 vdd.n32856 0.003
R67674 vdd.n37529 vdd.n37528 0.003
R67675 vdd.n37538 vdd.n37537 0.003
R67676 vdd.n37537 vdd.n37535 0.003
R67677 vdd.n35673 vdd.n35672 0.003
R67678 vdd.n32835 vdd.n32834 0.003
R67679 vdd.n37574 vdd.n37562 0.003
R67680 vdd.n38200 vdd.n38198 0.003
R67681 vdd.n38186 vdd.n38184 0.003
R67682 vdd.n30682 vdd.n30678 0.003
R67683 vdd.n30636 vdd.n30194 0.003
R67684 vdd.n29862 vdd.n29861 0.003
R67685 vdd.n27943 vdd.n27917 0.003
R67686 vdd.n27847 vdd.n27843 0.003
R67687 vdd.n27798 vdd.n27797 0.003
R67688 vdd.n28073 vdd.n28072 0.003
R67689 vdd.n30202 vdd.n30201 0.003
R67690 vdd.n30238 vdd.n30230 0.003
R67691 vdd.n30254 vdd.n30250 0.003
R67692 vdd.n30248 vdd.n30247 0.003
R67693 vdd.n28853 vdd.n28852 0.003
R67694 vdd.n28873 vdd.n28870 0.003
R67695 vdd.n28876 vdd.n28873 0.003
R67696 vdd.n28885 vdd.n28882 0.003
R67697 vdd.n28934 vdd.n28933 0.003
R67698 vdd.n29003 vdd.n28998 0.003
R67699 vdd.n29011 vdd.n29008 0.003
R67700 vdd.n29016 vdd.n29011 0.003
R67701 vdd.n28028 vdd.n28027 0.003
R67702 vdd.n28017 vdd.n28014 0.003
R67703 vdd.n27995 vdd.n27992 0.003
R67704 vdd.n27992 vdd.n27990 0.003
R67705 vdd.n27973 vdd.n27970 0.003
R67706 vdd.n29929 vdd.n29924 0.003
R67707 vdd.n29943 vdd.n29929 0.003
R67708 vdd.n29941 vdd.n29939 0.003
R67709 vdd.n29939 vdd.n29937 0.003
R67710 vdd.n29778 vdd.n29774 0.003
R67711 vdd.n30661 vdd.n30658 0.003
R67712 vdd.n30664 vdd.n30661 0.003
R67713 vdd.n30673 vdd.n30670 0.003
R67714 vdd.n30630 vdd.n30629 0.003
R67715 vdd.n30624 vdd.n30621 0.003
R67716 vdd.n30612 vdd.n30611 0.003
R67717 vdd.n30606 vdd.n30603 0.003
R67718 vdd.n30603 vdd.n30602 0.003
R67719 vdd.n30599 vdd.n30597 0.003
R67720 vdd.n30582 vdd.n30581 0.003
R67721 vdd.n30571 vdd.n30570 0.003
R67722 vdd.n30569 vdd.n30560 0.003
R67723 vdd.n30548 vdd.n30538 0.003
R67724 vdd.n30533 vdd.n30531 0.003
R67725 vdd.n27484 vdd.n27483 0.003
R67726 vdd.n27477 vdd.n27476 0.003
R67727 vdd.n27533 vdd.n27531 0.003
R67728 vdd.n27575 vdd.n27573 0.003
R67729 vdd.n27567 vdd.n27564 0.003
R67730 vdd.n27580 vdd.n27579 0.003
R67731 vdd.n27390 vdd.n27389 0.003
R67732 vdd.n27459 vdd.n27457 0.003
R67733 vdd.n27351 vdd.n27348 0.003
R67734 vdd.n29566 vdd.n29563 0.003
R67735 vdd.n25705 vdd.n25704 0.003
R67736 vdd.n25715 vdd.n25714 0.003
R67737 vdd.n25970 vdd.n25968 0.003
R67738 vdd.n25688 vdd.n25686 0.003
R67739 vdd.n25703 vdd.n25700 0.003
R67740 vdd.n25693 vdd.n25692 0.003
R67741 vdd.n25836 vdd.n25835 0.003
R67742 vdd.n25905 vdd.n25903 0.003
R67743 vdd.n25803 vdd.n25800 0.003
R67744 vdd.n25414 vdd.n25409 0.003
R67745 vdd.n25592 vdd.n25590 0.003
R67746 vdd.n25598 vdd.n25597 0.003
R67747 vdd.n25477 vdd.n25476 0.003
R67748 vdd.n30923 vdd.n30922 0.003
R67749 vdd.n30749 vdd.n30746 0.003
R67750 vdd.n30707 vdd.n30704 0.003
R67751 vdd.n30706 vdd.n30705 0.003
R67752 vdd.n32579 vdd.n32578 0.003
R67753 vdd.n32582 vdd.n32580 0.003
R67754 vdd.n29982 vdd.n29981 0.003
R67755 vdd.n29967 vdd.n29966 0.003
R67756 vdd.n29618 vdd.n29617 0.003
R67757 vdd.n32658 vdd.n32656 0.003
R67758 vdd.n27712 vdd.n27711 0.003
R67759 vdd.n26544 vdd.n26543 0.003
R67760 vdd.n26548 vdd.n26547 0.003
R67761 vdd.n25367 vdd.n25366 0.003
R67762 vdd.n31299 vdd.n31298 0.003
R67763 vdd.n31244 vdd.n31243 0.003
R67764 vdd.n26181 vdd.n26120 0.003
R67765 vdd.n26320 vdd.n26275 0.003
R67766 vdd.n29093 vdd.n29086 0.003
R67767 vdd.n29432 vdd.n29421 0.003
R67768 vdd.n32664 vdd.n32658 0.003
R67769 vdd.n31428 vdd.n31417 0.003
R67770 vdd.n30831 vdd.n30820 0.003
R67771 vdd.n30767 vdd.n30749 0.003
R67772 vdd.n31371 vdd.n31370 0.003
R67773 vdd.n30975 vdd.n30968 0.003
R67774 vdd.n26241 vdd.n26237 0.003
R67775 vdd.n26549 vdd.n26548 0.003
R67776 vdd.n27695 vdd.n27693 0.003
R67777 vdd.n29380 vdd.n29376 0.003
R67778 vdd.n29481 vdd.n29479 0.003
R67779 vdd.n29601 vdd.n29599 0.003
R67780 vdd.n30025 vdd.n30020 0.003
R67781 vdd.n32605 vdd.n32601 0.003
R67782 vdd.n30164 vdd.n30163 0.003
R67783 vdd.n30905 vdd.n30903 0.003
R67784 vdd.n2241 vdd.n2208 0.003
R67785 vdd.n2119 vdd.n2118 0.003
R67786 vdd.n2322 vdd.n2117 0.003
R67787 vdd.n2540 vdd.n2428 0.003
R67788 vdd.n3674 vdd.n3673 0.003
R67789 vdd.n4004 vdd.n4002 0.003
R67790 vdd.n3992 vdd.n3989 0.003
R67791 vdd.n3968 vdd.n3967 0.003
R67792 vdd.n3958 vdd.n3956 0.003
R67793 vdd.n3875 vdd.n3873 0.003
R67794 vdd.n3863 vdd.n3861 0.003
R67795 vdd.n2244 vdd.n2242 0.003
R67796 vdd.n2251 vdd.n2250 0.003
R67797 vdd.n2314 vdd.n2311 0.003
R67798 vdd.n2330 vdd.n2327 0.003
R67799 vdd.n2356 vdd.n2355 0.003
R67800 vdd.n2370 vdd.n2369 0.003
R67801 vdd.n2560 vdd.n2393 0.003
R67802 vdd.n2488 vdd.n2486 0.003
R67803 vdd.n2627 vdd.n2625 0.003
R67804 vdd.n2642 vdd.n2637 0.003
R67805 vdd.n2095 vdd.n2092 0.003
R67806 vdd.n2080 vdd.n2077 0.003
R67807 vdd.n1917 vdd.n1915 0.003
R67808 vdd.n1913 vdd.n1912 0.003
R67809 vdd.n1809 vdd.n1807 0.003
R67810 vdd.n26621 vdd.n26620 0.003
R67811 vdd.n26707 vdd.n26706 0.003
R67812 vdd.n27239 vdd.n27238 0.003
R67813 vdd.n26170 vdd.n26169 0.003
R67814 vdd.n26178 vdd.n26170 0.003
R67815 vdd.n26337 vdd.n26336 0.003
R67816 vdd.n31787 vdd.n31786 0.003
R67817 vdd.n31791 vdd.n31788 0.003
R67818 vdd.n31838 vdd.n31833 0.003
R67819 vdd.n31858 vdd.n31855 0.003
R67820 vdd.n31863 vdd.n31858 0.003
R67821 vdd.n31954 vdd.n31953 0.003
R67822 vdd.n31965 vdd.n31964 0.003
R67823 vdd.n31967 vdd.n31965 0.003
R67824 vdd.n32010 vdd.n32007 0.003
R67825 vdd.n32037 vdd.n32034 0.003
R67826 vdd.n32088 vdd.n32087 0.003
R67827 vdd.n32109 vdd.n32108 0.003
R67828 vdd.n32111 vdd.n32110 0.003
R67829 vdd.n32135 vdd.n32134 0.003
R67830 vdd.n32163 vdd.n32162 0.003
R67831 vdd.n32199 vdd.n32194 0.003
R67832 vdd.n32216 vdd.n32213 0.003
R67833 vdd.n32221 vdd.n32216 0.003
R67834 vdd.n32310 vdd.n32308 0.003
R67835 vdd.n32321 vdd.n32320 0.003
R67836 vdd.n32323 vdd.n32321 0.003
R67837 vdd.n32365 vdd.n32362 0.003
R67838 vdd.n32378 vdd.n32375 0.003
R67839 vdd.n32528 vdd.n32525 0.003
R67840 vdd.n32520 vdd.n32517 0.003
R67841 vdd.n32500 vdd.n32498 0.003
R67842 vdd.n32495 vdd.n32492 0.003
R67843 vdd.n32468 vdd.n32466 0.003
R67844 vdd.n32466 vdd.n32465 0.003
R67845 vdd.n31086 vdd.n31081 0.003
R67846 vdd.n31110 vdd.n31107 0.003
R67847 vdd.n31115 vdd.n31110 0.003
R67848 vdd.n32520 vdd.n32519 0.003
R67849 vdd.n31071 vdd.n31070 0.003
R67850 vdd.n31102 vdd.n31101 0.003
R67851 vdd.n29313 vdd.n29312 0.003
R67852 vdd.n32737 vdd.n7187 0.003
R67853 vdd.n32653 vdd.n32652 0.003
R67854 vdd.n29975 vdd.n29974 0.003
R67855 vdd.n30106 vdd.n30105 0.003
R67856 vdd.n30769 vdd.n30768 0.003
R67857 vdd.n31290 vdd.n31249 0.003
R67858 vdd.n26162 vdd.n26160 0.003
R67859 vdd.n31302 vdd.n31301 0.003
R67860 vdd.n26157 vdd.n26146 0.003
R67861 vdd.n26164 vdd.n26163 0.003
R67862 vdd.n26709 vdd.n26708 0.003
R67863 vdd.n26519 vdd.n26517 0.003
R67864 vdd.n29092 vdd.n29091 0.003
R67865 vdd.n29238 vdd.n29237 0.003
R67866 vdd.n7176 vdd.n7174 0.003
R67867 vdd.n12582 vdd.n12581 0.003
R67868 vdd.n10257 vdd.n10256 0.003
R67869 vdd.n10223 vdd.n10075 0.003
R67870 vdd.n10570 vdd.n10567 0.003
R67871 vdd.n12466 vdd.n10602 0.003
R67872 vdd.n12388 vdd.n12387 0.003
R67873 vdd.n10791 vdd.n10790 0.003
R67874 vdd.n10934 vdd.n10933 0.003
R67875 vdd.n10971 vdd.n10950 0.003
R67876 vdd.n12186 vdd.n12185 0.003
R67877 vdd.n12169 vdd.n12168 0.003
R67878 vdd.n11266 vdd.n11265 0.003
R67879 vdd.n11300 vdd.n11299 0.003
R67880 vdd.n11478 vdd.n11477 0.003
R67881 vdd.n11519 vdd.n11461 0.003
R67882 vdd.n11515 vdd.n11461 0.003
R67883 vdd.n11462 vdd.n11455 0.003
R67884 vdd.n11533 vdd.n11532 0.003
R67885 vdd.n11539 vdd.n11450 0.003
R67886 vdd.n11940 vdd.n11939 0.003
R67887 vdd.n11592 vdd.n11587 0.003
R67888 vdd.n11596 vdd.n11595 0.003
R67889 vdd.n11596 vdd.n11585 0.003
R67890 vdd.n13876 vdd.n8700 0.003
R67891 vdd.n14100 vdd.n8529 0.003
R67892 vdd.n14165 vdd.n8477 0.003
R67893 vdd.n14391 vdd.n14387 0.003
R67894 vdd.n14448 vdd.n14447 0.003
R67895 vdd.n13813 vdd.n8742 0.003
R67896 vdd.n11618 vdd.n11611 0.003
R67897 vdd.n11614 vdd.n11613 0.003
R67898 vdd.n13137 vdd.n9254 0.003
R67899 vdd.n9257 vdd.n9236 0.003
R67900 vdd.n13223 vdd.n13222 0.003
R67901 vdd.n9138 vdd.n9136 0.003
R67902 vdd.n13515 vdd.n13514 0.003
R67903 vdd.n8916 vdd.n8914 0.003
R67904 vdd.n11513 vdd.n11512 0.003
R67905 vdd.n11541 vdd.n11540 0.003
R67906 vdd.n10204 vdd.n10203 0.003
R67907 vdd.n10460 vdd.n10459 0.003
R67908 vdd.n10436 vdd.n10435 0.003
R67909 vdd.n9338 vdd.n9311 0.003
R67910 vdd.n9372 vdd.n9351 0.003
R67911 vdd.n9514 vdd.n9512 0.003
R67912 vdd.n9547 vdd.n9546 0.003
R67913 vdd.n9698 vdd.n9672 0.003
R67914 vdd.n9732 vdd.n9711 0.003
R67915 vdd.n9874 vdd.n9872 0.003
R67916 vdd.n9907 vdd.n9906 0.003
R67917 vdd.n10149 vdd.n10032 0.003
R67918 vdd.n10172 vdd.n10145 0.003
R67919 vdd.n13124 vdd.n13123 0.003
R67920 vdd.n13125 vdd.n9218 0.003
R67921 vdd.n13194 vdd.n13193 0.003
R67922 vdd.n13293 vdd.n13292 0.003
R67923 vdd.n13371 vdd.n13370 0.003
R67924 vdd.n13398 vdd.n9050 0.003
R67925 vdd.n13503 vdd.n13502 0.003
R67926 vdd.n13505 vdd.n13504 0.003
R67927 vdd.n13543 vdd.n8954 0.003
R67928 vdd.n13542 vdd.n8941 0.003
R67929 vdd.n13663 vdd.n13662 0.003
R67930 vdd.n13691 vdd.n8829 0.003
R67931 vdd.n13783 vdd.n13782 0.003
R67932 vdd.n13786 vdd.n13785 0.003
R67933 vdd.n13828 vdd.n8735 0.003
R67934 vdd.n13827 vdd.n8725 0.003
R67935 vdd.n8669 vdd.n8662 0.003
R67936 vdd.n13982 vdd.n8608 0.003
R67937 vdd.n14075 vdd.n8517 0.003
R67938 vdd.n14114 vdd.n14113 0.003
R67939 vdd.n14112 vdd.n14111 0.003
R67940 vdd.n8520 vdd.n8504 0.003
R67941 vdd.n8446 vdd.n8441 0.003
R67942 vdd.n14272 vdd.n8386 0.003
R67943 vdd.n14321 vdd.n8354 0.003
R67944 vdd.n8250 vdd.n8247 0.003
R67945 vdd.n8257 vdd.n8256 0.003
R67946 vdd.n14493 vdd.n14492 0.003
R67947 vdd.n8156 vdd.n8137 0.003
R67948 vdd.n14667 vdd.n14666 0.003
R67949 vdd.n8132 vdd.n8130 0.003
R67950 vdd.n14735 vdd.n14734 0.003
R67951 vdd.n14724 vdd.n8097 0.003
R67952 vdd.n14754 vdd.n14753 0.003
R67953 vdd.n14812 vdd.n8047 0.003
R67954 vdd.n14839 vdd.n14838 0.003
R67955 vdd.n8042 vdd.n8040 0.003
R67956 vdd.n14889 vdd.n14888 0.003
R67957 vdd.n14920 vdd.n14919 0.003
R67958 vdd.n14921 vdd.n8004 0.003
R67959 vdd.n24367 vdd.n24366 0.003
R67960 vdd.n24366 vdd.n24354 0.003
R67961 vdd.n24250 vdd.n24249 0.003
R67962 vdd.n24249 vdd.n24237 0.003
R67963 vdd.n22422 vdd.n22421 0.003
R67964 vdd.n22421 vdd.n22409 0.003
R67965 vdd.n15054 vdd.n15049 0.003
R67966 vdd.n15120 vdd.n15066 0.003
R67967 vdd.n16680 vdd.n16679 0.003
R67968 vdd.n16968 vdd.n16967 0.003
R67969 vdd.n17012 vdd.n16998 0.003
R67970 vdd.n17240 vdd.n17239 0.003
R67971 vdd.n17284 vdd.n17270 0.003
R67972 vdd.n17512 vdd.n17511 0.003
R67973 vdd.n17556 vdd.n17542 0.003
R67974 vdd.n17770 vdd.n17769 0.003
R67975 vdd.n17814 vdd.n17800 0.003
R67976 vdd.n18041 vdd.n18040 0.003
R67977 vdd.n18085 vdd.n18071 0.003
R67978 vdd.n18307 vdd.n18306 0.003
R67979 vdd.n18352 vdd.n18351 0.003
R67980 vdd.n18356 vdd.n18352 0.003
R67981 vdd.n18358 vdd.n18357 0.003
R67982 vdd.n18370 vdd.n18369 0.003
R67983 vdd.n18378 vdd.n18377 0.003
R67984 vdd.n18403 vdd.n18393 0.003
R67985 vdd.n18408 vdd.n18407 0.003
R67986 vdd.n18415 vdd.n18414 0.003
R67987 vdd.n21700 vdd.n18415 0.003
R67988 vdd.n19130 vdd.n19119 0.003
R67989 vdd.n18924 vdd.n18922 0.003
R67990 vdd.n18872 vdd.n18860 0.003
R67991 vdd.n18665 vdd.n18663 0.003
R67992 vdd.n18613 vdd.n18601 0.003
R67993 vdd.n21031 vdd.n21029 0.003
R67994 vdd.n21652 vdd.n21651 0.003
R67995 vdd.n21676 vdd.n21653 0.003
R67996 vdd.n21687 vdd.n21684 0.003
R67997 vdd.n21623 vdd.n21621 0.003
R67998 vdd.n21549 vdd.n21547 0.003
R67999 vdd.n21497 vdd.n21485 0.003
R68000 vdd.n21290 vdd.n21288 0.003
R68001 vdd.n21238 vdd.n21226 0.003
R68002 vdd.n18418 vdd.n18417 0.003
R68003 vdd.n18422 vdd.n18421 0.003
R68004 vdd.n16781 vdd.n16780 0.003
R68005 vdd.n15293 vdd.n15292 0.003
R68006 vdd.n15342 vdd.n15330 0.003
R68007 vdd.n15518 vdd.n15517 0.003
R68008 vdd.n15579 vdd.n15564 0.003
R68009 vdd.n15774 vdd.n15773 0.003
R68010 vdd.n15835 vdd.n15820 0.003
R68011 vdd.n16030 vdd.n16029 0.003
R68012 vdd.n16091 vdd.n16076 0.003
R68013 vdd.n16286 vdd.n16285 0.003
R68014 vdd.n16347 vdd.n16332 0.003
R68015 vdd.n16542 vdd.n16541 0.003
R68016 vdd.n16764 vdd.n16763 0.003
R68017 vdd.n20692 vdd.n20680 0.003
R68018 vdd.n20581 vdd.n20579 0.003
R68019 vdd.n20567 vdd.n20565 0.003
R68020 vdd.n20551 vdd.n20549 0.003
R68021 vdd.n20458 vdd.n20456 0.003
R68022 vdd.n20454 vdd.n20443 0.003
R68023 vdd.n20439 vdd.n20427 0.003
R68024 vdd.n20351 vdd.n20349 0.003
R68025 vdd.n20335 vdd.n20333 0.003
R68026 vdd.n20321 vdd.n20319 0.003
R68027 vdd.n20223 vdd.n20221 0.003
R68028 vdd.n20219 vdd.n20207 0.003
R68029 vdd.n20203 vdd.n20191 0.003
R68030 vdd.n20115 vdd.n20113 0.003
R68031 vdd.n20099 vdd.n20097 0.003
R68032 vdd.n20085 vdd.n20083 0.003
R68033 vdd.n19520 vdd.n19519 0.003
R68034 vdd.n19529 vdd.n19527 0.003
R68035 vdd.n19609 vdd.n19608 0.003
R68036 vdd.n19625 vdd.n19624 0.003
R68037 vdd.n19638 vdd.n19626 0.003
R68038 vdd.n19651 vdd.n19639 0.003
R68039 vdd.n19721 vdd.n19720 0.003
R68040 vdd.n19730 vdd.n19728 0.003
R68041 vdd.n19811 vdd.n19810 0.003
R68042 vdd.n19827 vdd.n19826 0.003
R68043 vdd.n19830 vdd.n19829 0.003
R68044 vdd.n20996 vdd.n19831 0.003
R68045 vdd.n20927 vdd.n20925 0.003
R68046 vdd.n20918 vdd.n20917 0.003
R68047 vdd.n20859 vdd.n20847 0.003
R68048 vdd.n20846 vdd.n20831 0.003
R68049 vdd.n20830 vdd.n20829 0.003
R68050 vdd.n20817 vdd.n20816 0.003
R68051 vdd.n20738 vdd.n20736 0.003
R68052 vdd.n20729 vdd.n20728 0.003
R68053 vdd.n19342 vdd.n19340 0.003
R68054 vdd.n19358 vdd.n19356 0.003
R68055 vdd.n19372 vdd.n19370 0.003
R68056 vdd.n19483 vdd.n19471 0.003
R68057 vdd.n24908 vdd.n24907 0.003
R68058 vdd.n24707 vdd.n24705 0.003
R68059 vdd.n24709 vdd.n24707 0.003
R68060 vdd.n24786 vdd.n24784 0.003
R68061 vdd.n24794 vdd.n24786 0.003
R68062 vdd.n25212 vdd.n25204 0.003
R68063 vdd.n25204 vdd.n25202 0.003
R68064 vdd.n25127 vdd.n25125 0.003
R68065 vdd.n25125 vdd.n25123 0.003
R68066 vdd.n35606 vdd.n35605 0.003
R68067 vdd.n35342 vdd.n35341 0.003
R68068 vdd.n35018 vdd.n35017 0.003
R68069 vdd.n34758 vdd.n34757 0.003
R68070 vdd.n5765 vdd.n5764 0.003
R68071 vdd.n5505 vdd.n5504 0.003
R68072 vdd.n4595 vdd.n4594 0.003
R68073 vdd.n4332 vdd.n4331 0.003
R68074 vdd.n30597 vdd.n30594 0.003
R68075 vdd.n31336 vdd.n31335 0.003
R68076 vdd.n31241 vdd.n31240 0.003
R68077 vdd.n25362 vdd.n25361 0.003
R68078 vdd.n32599 vdd.n32597 0.003
R68079 vdd.n29374 vdd.n29372 0.003
R68080 vdd.n26235 vdd.n26233 0.003
R68081 vdd.n6045 vdd.n6044 0.003
R68082 vdd.n5859 vdd.n5858 0.003
R68083 vdd.n475 vdd.n474 0.003
R68084 vdd.n197 vdd.n196 0.003
R68085 vdd.n319 vdd.n318 0.003
R68086 vdd.n34070 vdd.n34069 0.003
R68087 vdd.n34343 vdd.n34342 0.003
R68088 vdd.n33461 vdd.n33460 0.003
R68089 vdd.n26107 vdd.n26106 0.003
R68090 vdd.n32056 vdd.n32055 0.003
R68091 vdd.n31007 vdd.n31006 0.003
R68092 vdd.n26257 vdd.n26256 0.003
R68093 vdd.n29397 vdd.n29396 0.003
R68094 vdd.n26452 vdd.n26451 0.003
R68095 vdd.n31011 vdd.n31007 0.003
R68096 vdd.n3879 vdd.n3878 0.003
R68097 vdd.n30954 vdd.n30953 0.003
R68098 vdd.n2546 vdd.n2545 0.003
R68099 vdd.n26108 vdd.n26107 0.003
R68100 vdd.n26140 vdd.n26139 0.003
R68101 vdd.n27688 vdd.n27687 0.003
R68102 vdd.n29595 vdd.n29594 0.003
R68103 vdd.n30898 vdd.n30897 0.003
R68104 vdd.n32535 vdd.n32534 0.003
R68105 vdd.n31005 vdd.n31003 0.003
R68106 vdd.n31199 vdd.n31198 0.003
R68107 vdd.n4705 vdd.n4704 0.003
R68108 vdd.n773 vdd.n772 0.003
R68109 vdd.n30819 vdd.n30818 0.003
R68110 vdd.n30093 vdd.n30092 0.003
R68111 vdd.n29300 vdd.n29299 0.003
R68112 vdd.n26653 vdd.n26652 0.003
R68113 vdd.n6354 vdd.n6353 0.003
R68114 vdd.n2249 vdd.n2202 0.003
R68115 vdd.n30265 vdd.n30264 0.002
R68116 vdd.n30277 vdd.n30265 0.002
R68117 vdd.n29947 vdd.n29946 0.002
R68118 vdd.n681 vdd.n680 0.002
R68119 vdd.n1152 vdd.n1151 0.002
R68120 vdd.n853 vdd.n852 0.002
R68121 vdd.n30592 vdd.n30591 0.002
R68122 vdd.n30557 vdd.n30554 0.002
R68123 vdd.n30554 vdd.n30553 0.002
R68124 vdd.n30583 vdd.n30582 0.002
R68125 vdd.n30140 vdd.n30139 0.002
R68126 vdd.n29354 vdd.n29353 0.002
R68127 vdd.n29191 vdd.n29190 0.002
R68128 vdd.n26564 vdd.n26563 0.002
R68129 vdd.n25264 vdd.n7962 0.002
R68130 vdd.n31210 vdd.n31209 0.002
R68131 vdd.n31419 vdd.n31418 0.002
R68132 vdd.n27735 vdd.n27734 0.002
R68133 vdd.n32721 vdd.n32720 0.002
R68134 vdd.n31002 vdd.n31000 0.002
R68135 vdd.n31000 vdd.n30999 0.002
R68136 vdd.n5067 vdd.n5066 0.002
R68137 vdd.n29069 vdd.n29068 0.002
R68138 vdd.n35618 vdd.n35617 0.002
R68139 vdd.n35616 vdd.n35615 0.002
R68140 vdd.n35030 vdd.n35029 0.002
R68141 vdd.n6363 vdd.n6362 0.002
R68142 vdd.n6361 vdd.n5777 0.002
R68143 vdd.n5776 vdd.n5191 0.002
R68144 vdd.n5190 vdd.n4607 0.002
R68145 vdd.n34444 vdd.n6363 0.002
R68146 vdd.n29654 vdd.n29653 0.002
R68147 vdd.n27732 vdd.n27731 0.002
R68148 vdd.n31233 vdd.n31231 0.002
R68149 vdd.n30740 vdd.n30739 0.002
R68150 vdd.n30781 vdd.n30780 0.002
R68151 vdd.n32529 vdd.n32528 0.002
R68152 vdd.n6373 vdd.n6372 0.002
R68153 vdd.n6347 vdd.n6346 0.002
R68154 vdd.n576 vdd.n575 0.002
R68155 vdd.n206 vdd.n205 0.002
R68156 vdd.n306 vdd.n305 0.002
R68157 vdd.n33366 vdd.n33365 0.002
R68158 vdd.n33697 vdd.n33696 0.002
R68159 vdd.n33789 vdd.n33788 0.002
R68160 vdd.n2536 vdd.n2535 0.002
R68161 vdd.n32389 vdd.n32388 0.002
R68162 vdd.n3903 vdd.n3892 0.002
R68163 vdd.n24525 vdd.n24524 0.002
R68164 vdd.n32814 vdd.n32813 0.002
R68165 vdd.n30998 vdd.n30997 0.002
R68166 vdd.n34081 vdd.n34077 0.002
R68167 vdd.n35240 vdd.n35236 0.002
R68168 vdd.n34653 vdd.n34649 0.002
R68169 vdd.n5783 vdd.n5779 0.002
R68170 vdd.n5400 vdd.n5396 0.002
R68171 vdd.n4806 vdd.n4805 0.002
R68172 vdd.n4230 vdd.n4226 0.002
R68173 vdd.n29258 vdd.n29255 0.002
R68174 vdd.n26654 vdd.n26653 0.002
R68175 vdd.n29301 vdd.n29300 0.002
R68176 vdd.n30094 vdd.n30093 0.002
R68177 vdd.n31197 vdd.n31196 0.002
R68178 vdd.n31223 vdd.n31222 0.002
R68179 vdd.n31014 vdd.n31012 0.002
R68180 vdd.n2529 vdd.n2519 0.002
R68181 vdd.n30754 vdd.n30753 0.002
R68182 vdd.n1886 vdd.n1885 0.002
R68183 vdd.n3887 vdd.n3886 0.002
R68184 vdd.n34339 vdd.n34338 0.002
R68185 vdd.n34221 vdd.n34220 0.002
R68186 vdd.n2798 vdd.n2796 0.002
R68187 vdd.n2804 vdd.n2802 0.002
R68188 vdd.n2979 vdd.n2977 0.002
R68189 vdd.n2985 vdd.n2983 0.002
R68190 vdd.n3160 vdd.n3158 0.002
R68191 vdd.n3166 vdd.n3164 0.002
R68192 vdd.n3341 vdd.n3339 0.002
R68193 vdd.n3347 vdd.n3345 0.002
R68194 vdd.n3522 vdd.n3520 0.002
R68195 vdd.n3528 vdd.n3526 0.002
R68196 vdd.n183 vdd.n180 0.002
R68197 vdd.n316 vdd.n312 0.002
R68198 vdd.n311 vdd.n309 0.002
R68199 vdd.n4933 vdd.n4930 0.002
R68200 vdd.n2004 vdd.n2000 0.002
R68201 vdd.n35918 vdd.n35916 0.002
R68202 vdd.n35924 vdd.n35922 0.002
R68203 vdd.n36149 vdd.n36147 0.002
R68204 vdd.n36155 vdd.n36153 0.002
R68205 vdd.n36380 vdd.n36378 0.002
R68206 vdd.n36386 vdd.n36384 0.002
R68207 vdd.n36611 vdd.n36609 0.002
R68208 vdd.n36617 vdd.n36615 0.002
R68209 vdd.n36842 vdd.n36840 0.002
R68210 vdd.n36848 vdd.n36846 0.002
R68211 vdd.n36973 vdd.n36971 0.002
R68212 vdd.n36981 vdd.n36978 0.002
R68213 vdd.n36995 vdd.n36992 0.002
R68214 vdd.n37011 vdd.n37009 0.002
R68215 vdd.n37026 vdd.n37024 0.002
R68216 vdd.n37042 vdd.n37041 0.002
R68217 vdd.n37041 vdd.n37034 0.002
R68218 vdd.n33284 vdd.n33277 0.002
R68219 vdd.n37062 vdd.n37061 0.002
R68220 vdd.n37072 vdd.n37070 0.002
R68221 vdd.n33252 vdd.n33229 0.002
R68222 vdd.n33237 vdd.n33235 0.002
R68223 vdd.n37099 vdd.n37098 0.002
R68224 vdd.n37088 vdd.n37085 0.002
R68225 vdd.n33223 vdd.n33221 0.002
R68226 vdd.n33211 vdd.n33208 0.002
R68227 vdd.n37116 vdd.n37114 0.002
R68228 vdd.n33203 vdd.n33202 0.002
R68229 vdd.n33202 vdd.n33200 0.002
R68230 vdd.n37132 vdd.n37127 0.002
R68231 vdd.n37131 vdd.n37129 0.002
R68232 vdd.n33185 vdd.n33184 0.002
R68233 vdd.n33159 vdd.n33157 0.002
R68234 vdd.n37169 vdd.n37157 0.002
R68235 vdd.n37169 vdd.n37168 0.002
R68236 vdd.n37166 vdd.n37164 0.002
R68237 vdd.n35644 vdd.n35633 0.002
R68238 vdd.n35631 vdd.n35629 0.002
R68239 vdd.n37185 vdd.n37183 0.002
R68240 vdd.n33128 vdd.n33126 0.002
R68241 vdd.n37197 vdd.n37195 0.002
R68242 vdd.n33116 vdd.n33106 0.002
R68243 vdd.n33115 vdd.n33108 0.002
R68244 vdd.n33088 vdd.n33076 0.002
R68245 vdd.n33084 vdd.n33082 0.002
R68246 vdd.n33050 vdd.n33047 0.002
R68247 vdd.n37282 vdd.n37280 0.002
R68248 vdd.n33038 vdd.n33036 0.002
R68249 vdd.n37296 vdd.n37293 0.002
R68250 vdd.n37340 vdd.n37328 0.002
R68251 vdd.n37337 vdd.n37335 0.002
R68252 vdd.n37361 vdd.n37359 0.002
R68253 vdd.n32982 vdd.n32981 0.002
R68254 vdd.n37370 vdd.n37367 0.002
R68255 vdd.n37379 vdd.n37377 0.002
R68256 vdd.n32963 vdd.n32952 0.002
R68257 vdd.n37395 vdd.n37393 0.002
R68258 vdd.n37423 vdd.n37421 0.002
R68259 vdd.n37433 vdd.n37432 0.002
R68260 vdd.n37473 vdd.n37472 0.002
R68261 vdd.n32886 vdd.n32883 0.002
R68262 vdd.n37491 vdd.n37488 0.002
R68263 vdd.n32869 vdd.n32862 0.002
R68264 vdd.n32840 vdd.n32838 0.002
R68265 vdd.n32859 vdd.n32858 0.002
R68266 vdd.n32822 vdd.n32817 0.002
R68267 vdd.n32836 vdd.n32835 0.002
R68268 vdd.n37557 vdd.n37554 0.002
R68269 vdd.n37582 vdd.n37579 0.002
R68270 vdd.n38204 vdd.n38202 0.002
R68271 vdd.n38190 vdd.n38188 0.002
R68272 vdd.n38183 vdd.n38176 0.002
R68273 vdd.n38169 vdd.n38159 0.002
R68274 vdd.n37903 vdd.n37901 0.002
R68275 vdd.n37897 vdd.n37895 0.002
R68276 vdd.n37672 vdd.n37670 0.002
R68277 vdd.n37666 vdd.n37664 0.002
R68278 vdd.n28339 vdd.n28337 0.002
R68279 vdd.n28345 vdd.n28343 0.002
R68280 vdd.n28570 vdd.n28568 0.002
R68281 vdd.n28576 vdd.n28574 0.002
R68282 vdd.n28801 vdd.n28799 0.002
R68283 vdd.n1566 vdd.n1564 0.002
R68284 vdd.n1560 vdd.n1558 0.002
R68285 vdd.n1385 vdd.n1383 0.002
R68286 vdd.n1379 vdd.n1377 0.002
R68287 vdd.n26845 vdd.n26843 0.002
R68288 vdd.n26851 vdd.n26849 0.002
R68289 vdd.n27026 vdd.n27024 0.002
R68290 vdd.n27032 vdd.n27030 0.002
R68291 vdd.n27207 vdd.n27205 0.002
R68292 vdd.n26755 vdd.n26731 0.002
R68293 vdd.n31279 vdd.n31251 0.002
R68294 vdd.n29755 vdd.n29753 0.002
R68295 vdd.n29846 vdd.n29842 0.002
R68296 vdd.n29841 vdd.n29839 0.002
R68297 vdd.n27935 vdd.n27934 0.002
R68298 vdd.n27934 vdd.n27928 0.002
R68299 vdd.n27849 vdd.n27847 0.002
R68300 vdd.n27822 vdd.n27818 0.002
R68301 vdd.n27816 vdd.n27815 0.002
R68302 vdd.n28126 vdd.n28125 0.002
R68303 vdd.n28803 vdd.n28178 0.002
R68304 vdd.n30621 vdd.n30238 0.002
R68305 vdd.n28861 vdd.n28858 0.002
R68306 vdd.n28888 vdd.n28885 0.002
R68307 vdd.n28927 vdd.n28926 0.002
R68308 vdd.n28935 vdd.n28934 0.002
R68309 vdd.n28998 vdd.n28995 0.002
R68310 vdd.n29004 vdd.n29003 0.002
R68311 vdd.n28046 vdd.n28044 0.002
R68312 vdd.n28004 vdd.n28001 0.002
R68313 vdd.n27970 vdd.n27968 0.002
R68314 vdd.n27949 vdd.n27948 0.002
R68315 vdd.n27943 vdd.n27927 0.002
R68316 vdd.n29917 vdd.n29916 0.002
R68317 vdd.n29924 vdd.n29921 0.002
R68318 vdd.n29937 vdd.n29934 0.002
R68319 vdd.n29798 vdd.n29793 0.002
R68320 vdd.n29846 vdd.n29786 0.002
R68321 vdd.n29768 vdd.n29767 0.002
R68322 vdd.n29734 vdd.n29733 0.002
R68323 vdd.n29732 vdd.n29729 0.002
R68324 vdd.n30676 vdd.n30673 0.002
R68325 vdd.n30645 vdd.n30644 0.002
R68326 vdd.n30636 vdd.n30635 0.002
R68327 vdd.n30615 vdd.n30612 0.002
R68328 vdd.n30601 vdd.n30599 0.002
R68329 vdd.n30590 vdd.n30588 0.002
R68330 vdd.n30580 vdd.n30578 0.002
R68331 vdd.n30519 vdd.n30517 0.002
R68332 vdd.n25523 vdd.n25519 0.002
R68333 vdd.n31387 vdd.n31386 0.002
R68334 vdd.n31384 vdd.n31383 0.002
R68335 vdd.n31384 vdd.n31374 0.002
R68336 vdd.n32718 vdd.n32717 0.002
R68337 vdd.n32670 vdd.n32668 0.002
R68338 vdd.n29276 vdd.n29275 0.002
R68339 vdd.n29070 vdd.n29067 0.002
R68340 vdd.n25671 vdd.n25670 0.002
R68341 vdd.n32737 vdd.n7196 0.002
R68342 vdd.n32737 vdd.n7194 0.002
R68343 vdd.n26083 vdd.n25372 0.002
R68344 vdd.n31441 vdd.n31436 0.002
R68345 vdd.n31337 vdd.n31334 0.002
R68346 vdd.n32737 vdd.n7223 0.002
R68347 vdd.n6363 vdd.n589 0.002
R68348 vdd.n3673 vdd.n3672 0.002
R68349 vdd.n3675 vdd.n3674 0.002
R68350 vdd.n3720 vdd.n3717 0.002
R68351 vdd.n4016 vdd.n3720 0.002
R68352 vdd.n4012 vdd.n4007 0.002
R68353 vdd.n4007 vdd.n4004 0.002
R68354 vdd.n3997 vdd.n3992 0.002
R68355 vdd.n3989 vdd.n3987 0.002
R68356 vdd.n3982 vdd.n3977 0.002
R68357 vdd.n3969 vdd.n3968 0.002
R68358 vdd.n3967 vdd.n3966 0.002
R68359 vdd.n3956 vdd.n3955 0.002
R68360 vdd.n3955 vdd.n3947 0.002
R68361 vdd.n3932 vdd.n3930 0.002
R68362 vdd.n3930 vdd.n3929 0.002
R68363 vdd.n3906 vdd.n3904 0.002
R68364 vdd.n3889 vdd.n3887 0.002
R68365 vdd.n3877 vdd.n3875 0.002
R68366 vdd.n3864 vdd.n3863 0.002
R68367 vdd.n3845 vdd.n3843 0.002
R68368 vdd.n2220 vdd.n2219 0.002
R68369 vdd.n2225 vdd.n2222 0.002
R68370 vdd.n2242 vdd.n2241 0.002
R68371 vdd.n2247 vdd.n2244 0.002
R68372 vdd.n2252 vdd.n2251 0.002
R68373 vdd.n2293 vdd.n2290 0.002
R68374 vdd.n2294 vdd.n2293 0.002
R68375 vdd.n2308 vdd.n2303 0.002
R68376 vdd.n2311 vdd.n2308 0.002
R68377 vdd.n2327 vdd.n2322 0.002
R68378 vdd.n2333 vdd.n2330 0.002
R68379 vdd.n2346 vdd.n2341 0.002
R68380 vdd.n2355 vdd.n2354 0.002
R68381 vdd.n2361 vdd.n2356 0.002
R68382 vdd.n2387 vdd.n2370 0.002
R68383 vdd.n2392 vdd.n2387 0.002
R68384 vdd.n2558 vdd.n2557 0.002
R68385 vdd.n2550 vdd.n2549 0.002
R68386 vdd.n2542 vdd.n2540 0.002
R68387 vdd.n2540 vdd.n2539 0.002
R68388 vdd.n2505 vdd.n2503 0.002
R68389 vdd.n2503 vdd.n2501 0.002
R68390 vdd.n2490 vdd.n2488 0.002
R68391 vdd.n2471 vdd.n2469 0.002
R68392 vdd.n2603 vdd.n2602 0.002
R68393 vdd.n2608 vdd.n2605 0.002
R68394 vdd.n2625 vdd.n2624 0.002
R68395 vdd.n2630 vdd.n2627 0.002
R68396 vdd.n2644 vdd.n2642 0.002
R68397 vdd.n1998 vdd.n1995 0.002
R68398 vdd.n2092 vdd.n2089 0.002
R68399 vdd.n2082 vdd.n2080 0.002
R68400 vdd.n1950 vdd.n1949 0.002
R68401 vdd.n1925 vdd.n1924 0.002
R68402 vdd.n1924 vdd.n1923 0.002
R68403 vdd.n1923 vdd.n1922 0.002
R68404 vdd.n1912 vdd.n1897 0.002
R68405 vdd.n1897 vdd.n1896 0.002
R68406 vdd.n1890 vdd.n1889 0.002
R68407 vdd.n1841 vdd.n1839 0.002
R68408 vdd.n1831 vdd.n1829 0.002
R68409 vdd.n1829 vdd.n1827 0.002
R68410 vdd.n1810 vdd.n1809 0.002
R68411 vdd.n1790 vdd.n1788 0.002
R68412 vdd.n1783 vdd.n1775 0.002
R68413 vdd.n31881 vdd.n31690 0.002
R68414 vdd.n27240 vdd.n27239 0.002
R68415 vdd.n26169 vdd.n26168 0.002
R68416 vdd.n26198 vdd.n26196 0.002
R68417 vdd.n26213 vdd.n26199 0.002
R68418 vdd.n26600 vdd.n26598 0.002
R68419 vdd.n26691 vdd.n26690 0.002
R68420 vdd.n26683 vdd.n26682 0.002
R68421 vdd.n26682 vdd.n26680 0.002
R68422 vdd.n26297 vdd.n26296 0.002
R68423 vdd.n31758 vdd.n31745 0.002
R68424 vdd.n31759 vdd.n31758 0.002
R68425 vdd.n31786 vdd.n31785 0.002
R68426 vdd.n31804 vdd.n31799 0.002
R68427 vdd.n31806 vdd.n31805 0.002
R68428 vdd.n31807 vdd.n31806 0.002
R68429 vdd.n31824 vdd.n31819 0.002
R68430 vdd.n31833 vdd.n31830 0.002
R68431 vdd.n31849 vdd.n31838 0.002
R68432 vdd.n31868 vdd.n31863 0.002
R68433 vdd.n31880 vdd.n31875 0.002
R68434 vdd.n31953 vdd.n31951 0.002
R68435 vdd.n31964 vdd.n31962 0.002
R68436 vdd.n31978 vdd.n31976 0.002
R68437 vdd.n31981 vdd.n31979 0.002
R68438 vdd.n31993 vdd.n31991 0.002
R68439 vdd.n32011 vdd.n32010 0.002
R68440 vdd.n32019 vdd.n32016 0.002
R68441 vdd.n32022 vdd.n32019 0.002
R68442 vdd.n32044 vdd.n32043 0.002
R68443 vdd.n32078 vdd.n32077 0.002
R68444 vdd.n32079 vdd.n32078 0.002
R68445 vdd.n32087 vdd.n32084 0.002
R68446 vdd.n32108 vdd.n32107 0.002
R68447 vdd.n32117 vdd.n32116 0.002
R68448 vdd.n32162 vdd.n32149 0.002
R68449 vdd.n32164 vdd.n32163 0.002
R68450 vdd.n32185 vdd.n32177 0.002
R68451 vdd.n32194 vdd.n32191 0.002
R68452 vdd.n32204 vdd.n32199 0.002
R68453 vdd.n32232 vdd.n32221 0.002
R68454 vdd.n32248 vdd.n32245 0.002
R68455 vdd.n32253 vdd.n32248 0.002
R68456 vdd.n32308 vdd.n32307 0.002
R68457 vdd.n32320 vdd.n32318 0.002
R68458 vdd.n32336 vdd.n32334 0.002
R68459 vdd.n32340 vdd.n32337 0.002
R68460 vdd.n32353 vdd.n32351 0.002
R68461 vdd.n32366 vdd.n32365 0.002
R68462 vdd.n32381 vdd.n32378 0.002
R68463 vdd.n32534 vdd.n32533 0.002
R68464 vdd.n32525 vdd.n32524 0.002
R68465 vdd.n32523 vdd.n32520 0.002
R68466 vdd.n32492 vdd.n32487 0.002
R68467 vdd.n32471 vdd.n32468 0.002
R68468 vdd.n32457 vdd.n32454 0.002
R68469 vdd.n31051 vdd.n31050 0.002
R68470 vdd.n31071 vdd.n31063 0.002
R68471 vdd.n31081 vdd.n31078 0.002
R68472 vdd.n31097 vdd.n31086 0.002
R68473 vdd.n31120 vdd.n31115 0.002
R68474 vdd.n31187 vdd.n31186 0.002
R68475 vdd.n31186 vdd.n31184 0.002
R68476 vdd.n29187 vdd.n29186 0.002
R68477 vdd.n29284 vdd.n29283 0.002
R68478 vdd.n29336 vdd.n29284 0.002
R68479 vdd.n29312 vdd.n29311 0.002
R68480 vdd.n29296 vdd.n29295 0.002
R68481 vdd.n29419 vdd.n29418 0.002
R68482 vdd.n29432 vdd.n29419 0.002
R68483 vdd.n29464 vdd.n29435 0.002
R68484 vdd.n29437 vdd.n29436 0.002
R68485 vdd.n29532 vdd.n29531 0.002
R68486 vdd.n29531 vdd.n29530 0.002
R68487 vdd.n29514 vdd.n29513 0.002
R68488 vdd.n32664 vdd.n32653 0.002
R68489 vdd.n32667 vdd.n32666 0.002
R68490 vdd.n32681 vdd.n32680 0.002
R68491 vdd.n32703 vdd.n32681 0.002
R68492 vdd.n29644 vdd.n29643 0.002
R68493 vdd.n29671 vdd.n29644 0.002
R68494 vdd.n29976 vdd.n29975 0.002
R68495 vdd.n30043 vdd.n30042 0.002
R68496 vdd.n30059 vdd.n30043 0.002
R68497 vdd.n30077 vdd.n30076 0.002
R68498 vdd.n30125 vdd.n30077 0.002
R68499 vdd.n30105 vdd.n30104 0.002
R68500 vdd.n30089 vdd.n30088 0.002
R68501 vdd.n31415 vdd.n31414 0.002
R68502 vdd.n31428 vdd.n31415 0.002
R68503 vdd.n32563 vdd.n31431 0.002
R68504 vdd.n32536 vdd.n31441 0.002
R68505 vdd.n30814 vdd.n30813 0.002
R68506 vdd.n30778 vdd.n30777 0.002
R68507 vdd.n30777 vdd.n30776 0.002
R68508 vdd.n30768 vdd.n30767 0.002
R68509 vdd.n30742 vdd.n30741 0.002
R68510 vdd.n31193 vdd.n31192 0.002
R68511 vdd.n31225 vdd.n31193 0.002
R68512 vdd.n31236 vdd.n31228 0.002
R68513 vdd.n31239 vdd.n31238 0.002
R68514 vdd.n31247 vdd.n31239 0.002
R68515 vdd.n31247 vdd.n31246 0.002
R68516 vdd.n27245 vdd.n27243 0.002
R68517 vdd.n26180 vdd.n26164 0.002
R68518 vdd.n26217 vdd.n26215 0.002
R68519 vdd.n26622 vdd.n26585 0.002
R68520 vdd.n26711 vdd.n26622 0.002
R68521 vdd.n26708 vdd.n26673 0.002
R68522 vdd.n26671 vdd.n26670 0.002
R68523 vdd.n26319 vdd.n26286 0.002
R68524 vdd.n26320 vdd.n26319 0.002
R68525 vdd.n26407 vdd.n26351 0.002
R68526 vdd.n26405 vdd.n26404 0.002
R68527 vdd.n26404 vdd.n26391 0.002
R68528 vdd.n26523 vdd.n26522 0.002
R68529 vdd.n26474 vdd.n26473 0.002
R68530 vdd.n26473 vdd.n26472 0.002
R68531 vdd.n26468 vdd.n26467 0.002
R68532 vdd.n29093 vdd.n29092 0.002
R68533 vdd.n29096 vdd.n29095 0.002
R68534 vdd.n29100 vdd.n29099 0.002
R68535 vdd.n29101 vdd.n29100 0.002
R68536 vdd.n29136 vdd.n29118 0.002
R68537 vdd.n29165 vdd.n29163 0.002
R68538 vdd.n12600 vdd.n10070 0.002
R68539 vdd.n12600 vdd.n10076 0.002
R68540 vdd.n12600 vdd.n10091 0.002
R68541 vdd.n12600 vdd.n10079 0.002
R68542 vdd.n10223 vdd.n10222 0.002
R68543 vdd.n10266 vdd.n10255 0.002
R68544 vdd.n10223 vdd.n10134 0.002
R68545 vdd.n12600 vdd.n10087 0.002
R68546 vdd.n10683 vdd.n10659 0.002
R68547 vdd.n10695 vdd.n10677 0.002
R68548 vdd.n10851 vdd.n10850 0.002
R68549 vdd.n12329 vdd.n10852 0.002
R68550 vdd.n11024 vdd.n11017 0.002
R68551 vdd.n12229 vdd.n12228 0.002
R68552 vdd.n12128 vdd.n12127 0.002
R68553 vdd.n11205 vdd.n11204 0.002
R68554 vdd.n11360 vdd.n11359 0.002
R68555 vdd.n12023 vdd.n11361 0.002
R68556 vdd.n11503 vdd.n11435 0.002
R68557 vdd.n13956 vdd.n13955 0.002
R68558 vdd.n13998 vdd.n8585 0.002
R68559 vdd.n14246 vdd.n14245 0.002
R68560 vdd.n14289 vdd.n8365 0.002
R68561 vdd.n14543 vdd.n8178 0.002
R68562 vdd.n9254 vdd.n9251 0.002
R68563 vdd.n9083 vdd.n9059 0.002
R68564 vdd.n13433 vdd.n13432 0.002
R68565 vdd.n8863 vdd.n8839 0.002
R68566 vdd.n13725 vdd.n13724 0.002
R68567 vdd.n10335 vdd.n10332 0.002
R68568 vdd.n10373 vdd.n10352 0.002
R68569 vdd.n9428 vdd.n9426 0.002
R68570 vdd.n12980 vdd.n12979 0.002
R68571 vdd.n12895 vdd.n9602 0.002
R68572 vdd.n9643 vdd.n9642 0.002
R68573 vdd.n9788 vdd.n9786 0.002
R68574 vdd.n12772 vdd.n12771 0.002
R68575 vdd.n12687 vdd.n9962 0.002
R68576 vdd.n10003 vdd.n10002 0.002
R68577 vdd.n10162 vdd.n10161 0.002
R68578 vdd.n11768 vdd.n11675 0.002
R68579 vdd.n11718 vdd.n11686 0.002
R68580 vdd.n11699 vdd.n11698 0.002
R68581 vdd.n11711 vdd.n11700 0.002
R68582 vdd.n11862 vdd.n11809 0.002
R68583 vdd.n11858 vdd.n11857 0.002
R68584 vdd.n11851 vdd.n11839 0.002
R68585 vdd.n11912 vdd.n11909 0.002
R68586 vdd.n13085 vdd.n9284 0.002
R68587 vdd.n13123 vdd.n9270 0.002
R68588 vdd.n13126 vdd.n13125 0.002
R68589 vdd.n13193 vdd.n13192 0.002
R68590 vdd.n13292 vdd.n9147 0.002
R68591 vdd.n13341 vdd.n9100 0.002
R68592 vdd.n13343 vdd.n9066 0.002
R68593 vdd.n13397 vdd.n13396 0.002
R68594 vdd.n13416 vdd.n13415 0.002
R68595 vdd.n13488 vdd.n13487 0.002
R68596 vdd.n13476 vdd.n8999 0.002
R68597 vdd.n13565 vdd.n13564 0.002
R68598 vdd.n13585 vdd.n13584 0.002
R68599 vdd.n13633 vdd.n8879 0.002
R68600 vdd.n13635 vdd.n8846 0.002
R68601 vdd.n13689 vdd.n13688 0.002
R68602 vdd.n13710 vdd.n13709 0.002
R68603 vdd.n13768 vdd.n13767 0.002
R68604 vdd.n13756 vdd.n8782 0.002
R68605 vdd.n13853 vdd.n13846 0.002
R68606 vdd.n13847 vdd.n8687 0.002
R68607 vdd.n8688 vdd.n8673 0.002
R68608 vdd.n13910 vdd.n8671 0.002
R68609 vdd.n13984 vdd.n13983 0.002
R68610 vdd.n13985 vdd.n8570 0.002
R68611 vdd.n14046 vdd.n8571 0.002
R68612 vdd.n14044 vdd.n8556 0.002
R68613 vdd.n14142 vdd.n14135 0.002
R68614 vdd.n14136 vdd.n8463 0.002
R68615 vdd.n8465 vdd.n8449 0.002
R68616 vdd.n14200 vdd.n8447 0.002
R68617 vdd.n14274 vdd.n14273 0.002
R68618 vdd.n14275 vdd.n8353 0.002
R68619 vdd.n14321 vdd.n14320 0.002
R68620 vdd.n14457 vdd.n8247 0.002
R68621 vdd.n8256 vdd.n8219 0.002
R68622 vdd.n14495 vdd.n14493 0.002
R68623 vdd.n8156 vdd.n8152 0.002
R68624 vdd.n14668 vdd.n14667 0.002
R68625 vdd.n14679 vdd.n8130 0.002
R68626 vdd.n14736 vdd.n14735 0.002
R68627 vdd.n14724 vdd.n14721 0.002
R68628 vdd.n14755 vdd.n14754 0.002
R68629 vdd.n14812 vdd.n14808 0.002
R68630 vdd.n14840 vdd.n14839 0.002
R68631 vdd.n14851 vdd.n8040 0.002
R68632 vdd.n14889 vdd.n14883 0.002
R68633 vdd.n14919 vdd.n8013 0.002
R68634 vdd.n14935 vdd.n8004 0.002
R68635 vdd.n22341 vdd.n22256 0.002
R68636 vdd.n22343 vdd.n22230 0.002
R68637 vdd.n22363 vdd.n22362 0.002
R68638 vdd.n24304 vdd.n22133 0.002
R68639 vdd.n24306 vdd.n22117 0.002
R68640 vdd.n24308 vdd.n22091 0.002
R68641 vdd.n22308 vdd.n22307 0.002
R68642 vdd.n22293 vdd.n22292 0.002
R68643 vdd.n24351 vdd.n24339 0.002
R68644 vdd.n24280 vdd.n24279 0.002
R68645 vdd.n24265 vdd.n24264 0.002
R68646 vdd.n24234 vdd.n24222 0.002
R68647 vdd.n24094 vdd.n24092 0.002
R68648 vdd.n24082 vdd.n24080 0.002
R68649 vdd.n23862 vdd.n23860 0.002
R68650 vdd.n23850 vdd.n23848 0.002
R68651 vdd.n23630 vdd.n23628 0.002
R68652 vdd.n23162 vdd.n23160 0.002
R68653 vdd.n23174 vdd.n23172 0.002
R68654 vdd.n23394 vdd.n23392 0.002
R68655 vdd.n23406 vdd.n23404 0.002
R68656 vdd.n23626 vdd.n23624 0.002
R68657 vdd.n22583 vdd.n22581 0.002
R68658 vdd.n22595 vdd.n22593 0.002
R68659 vdd.n22815 vdd.n22813 0.002
R68660 vdd.n22827 vdd.n22825 0.002
R68661 vdd.n23050 vdd.n23045 0.002
R68662 vdd.n22452 vdd.n22451 0.002
R68663 vdd.n22437 vdd.n22436 0.002
R68664 vdd.n22406 vdd.n22394 0.002
R68665 vdd.n16743 vdd.n16595 0.002
R68666 vdd.n16743 vdd.n16689 0.002
R68667 vdd.n16743 vdd.n16738 0.002
R68668 vdd.n16743 vdd.n16702 0.002
R68669 vdd.n16679 vdd.n16672 0.002
R68670 vdd.n15040 vdd.n15039 0.002
R68671 vdd.n16679 vdd.n16600 0.002
R68672 vdd.n16743 vdd.n16730 0.002
R68673 vdd.n17109 vdd.n17108 0.002
R68674 vdd.n17143 vdd.n17129 0.002
R68675 vdd.n17381 vdd.n17380 0.002
R68676 vdd.n17415 vdd.n17401 0.002
R68677 vdd.n17639 vdd.n17638 0.002
R68678 vdd.n17673 vdd.n17659 0.002
R68679 vdd.n17910 vdd.n17909 0.002
R68680 vdd.n17944 vdd.n17930 0.002
R68681 vdd.n18182 vdd.n18181 0.002
R68682 vdd.n18216 vdd.n18202 0.002
R68683 vdd.n18331 vdd.n18330 0.002
R68684 vdd.n19039 vdd.n19037 0.002
R68685 vdd.n19006 vdd.n19004 0.002
R68686 vdd.n18780 vdd.n18778 0.002
R68687 vdd.n18747 vdd.n18745 0.002
R68688 vdd.n18521 vdd.n18519 0.002
R68689 vdd.n21684 vdd.n21683 0.002
R68690 vdd.n21405 vdd.n21403 0.002
R68691 vdd.n21372 vdd.n21370 0.002
R68692 vdd.n21146 vdd.n21144 0.002
R68693 vdd.n21113 vdd.n21111 0.002
R68694 vdd.n15415 vdd.n15414 0.002
R68695 vdd.n15432 vdd.n15420 0.002
R68696 vdd.n15665 vdd.n15664 0.002
R68697 vdd.n15685 vdd.n15670 0.002
R68698 vdd.n15921 vdd.n15920 0.002
R68699 vdd.n15941 vdd.n15926 0.002
R68700 vdd.n16177 vdd.n16176 0.002
R68701 vdd.n16197 vdd.n16182 0.002
R68702 vdd.n16433 vdd.n16432 0.002
R68703 vdd.n16453 vdd.n16438 0.002
R68704 vdd.n16576 vdd.n16575 0.002
R68705 vdd.n20680 vdd.n20678 0.002
R68706 vdd.n20583 vdd.n20581 0.002
R68707 vdd.n20565 vdd.n20563 0.002
R68708 vdd.n20549 vdd.n20547 0.002
R68709 vdd.n20464 vdd.n20458 0.002
R68710 vdd.n20443 vdd.n20441 0.002
R68711 vdd.n20427 vdd.n20425 0.002
R68712 vdd.n20353 vdd.n20351 0.002
R68713 vdd.n20337 vdd.n20335 0.002
R68714 vdd.n20319 vdd.n20317 0.002
R68715 vdd.n20235 vdd.n20223 0.002
R68716 vdd.n20207 vdd.n20205 0.002
R68717 vdd.n20191 vdd.n20189 0.002
R68718 vdd.n20117 vdd.n20115 0.002
R68719 vdd.n20101 vdd.n20099 0.002
R68720 vdd.n20083 vdd.n20081 0.002
R68721 vdd.n19502 vdd.n19500 0.002
R68722 vdd.n19517 vdd.n19516 0.002
R68723 vdd.n19532 vdd.n19530 0.002
R68724 vdd.n19548 vdd.n19546 0.002
R68725 vdd.n19578 vdd.n19576 0.002
R68726 vdd.n19594 vdd.n19592 0.002
R68727 vdd.n19667 vdd.n19655 0.002
R68728 vdd.n19683 vdd.n19671 0.002
R68729 vdd.n19703 vdd.n19701 0.002
R68730 vdd.n19718 vdd.n19717 0.002
R68731 vdd.n19734 vdd.n19732 0.002
R68732 vdd.n19750 vdd.n19748 0.002
R68733 vdd.n19780 vdd.n19778 0.002
R68734 vdd.n19796 vdd.n19794 0.002
R68735 vdd.n20993 vdd.n20991 0.002
R68736 vdd.n20977 vdd.n20975 0.002
R68737 vdd.n20947 vdd.n20945 0.002
R68738 vdd.n20931 vdd.n20929 0.002
R68739 vdd.n20915 vdd.n20914 0.002
R68740 vdd.n20900 vdd.n20898 0.002
R68741 vdd.n20880 vdd.n20868 0.002
R68742 vdd.n20864 vdd.n20863 0.002
R68743 vdd.n20802 vdd.n20800 0.002
R68744 vdd.n20786 vdd.n20784 0.002
R68745 vdd.n20757 vdd.n20755 0.002
R68746 vdd.n20741 vdd.n20739 0.002
R68747 vdd.n20726 vdd.n20725 0.002
R68748 vdd.n20711 vdd.n20709 0.002
R68749 vdd.n19340 vdd.n19338 0.002
R68750 vdd.n19356 vdd.n19354 0.002
R68751 vdd.n19374 vdd.n19372 0.002
R68752 vdd.n19471 vdd.n19469 0.002
R68753 vdd.n21853 vdd.n21851 0.002
R68754 vdd.n21771 vdd.n21770 0.002
R68755 vdd.n21793 vdd.n21791 0.002
R68756 vdd.n21785 vdd.n21783 0.002
R68757 vdd.n21953 vdd.n21900 0.002
R68758 vdd.n21949 vdd.n21948 0.002
R68759 vdd.n21942 vdd.n21930 0.002
R68760 vdd.n21749 vdd.n21748 0.002
R68761 vdd.n21746 vdd.n14976 0.002
R68762 vdd.n24932 vdd.n24916 0.002
R68763 vdd.n24885 vdd.n24884 0.002
R68764 vdd.n24622 vdd.n24621 0.002
R68765 vdd.n24631 vdd.n24629 0.002
R68766 vdd.n24683 vdd.n24681 0.002
R68767 vdd.n24695 vdd.n24693 0.002
R68768 vdd.n24721 vdd.n24719 0.002
R68769 vdd.n24730 vdd.n24722 0.002
R68770 vdd.n24774 vdd.n24772 0.002
R68771 vdd.n24806 vdd.n24798 0.002
R68772 vdd.n24818 vdd.n24810 0.002
R68773 vdd.n25236 vdd.n25228 0.002
R68774 vdd.n25224 vdd.n25216 0.002
R68775 vdd.n25192 vdd.n25190 0.002
R68776 vdd.n25139 vdd.n25137 0.002
R68777 vdd.n25113 vdd.n25111 0.002
R68778 vdd.n25101 vdd.n25099 0.002
R68779 vdd.n30560 vdd.n30558 0.002
R68780 vdd.n10249 vdd.n10224 0.002
R68781 vdd.n16670 vdd.n16604 0.002
R68782 vdd.n2549 vdd.n2548 0.002
R68783 vdd.n29641 vdd.n29636 0.002
R68784 vdd.n27246 vdd.n27245 0.002
R68785 vdd.n26297 vdd.n26292 0.002
R68786 vdd.n31221 vdd.n31218 0.002
R68787 vdd.n24908 vdd.n24903 0.002
R68788 vdd.n32534 vdd.n32390 0.002
R68789 vdd.n30951 vdd.n30950 0.002
R68790 vdd.n30952 vdd.n30951 0.002
R68791 vdd.n26673 vdd.n26655 0.002
R68792 vdd.n29311 vdd.n29298 0.002
R68793 vdd.n30104 vdd.n30091 0.002
R68794 vdd.n31355 vdd.n31354 0.002
R68795 vdd.n31230 vdd.n31229 0.002
R68796 vdd.n7219 vdd.n7211 0.002
R68797 vdd.n7177 vdd.n7176 0.002
R68798 vdd.n29714 vdd.n29713 0.002
R68799 vdd.n31785 vdd.n31784 0.002
R68800 vdd.n30756 vdd.n30755 0.002
R68801 vdd.n30510 vdd.n30509 0.002
R68802 vdd.n32739 vdd.n7116 0.002
R68803 vdd.n31196 vdd.n31195 0.002
R68804 vdd.n572 vdd.n571 0.002
R68805 vdd.n33362 vdd.n33361 0.002
R68806 vdd.n33686 vdd.n33685 0.002
R68807 vdd.n33852 vdd.n33851 0.002
R68808 vdd.n32763 vdd.n6892 0.002
R68809 vdd.n32766 vdd.n6862 0.002
R68810 vdd.n32772 vdd.n6808 0.002
R68811 vdd.n32778 vdd.n6748 0.002
R68812 vdd.n32782 vdd.n6695 0.002
R68813 vdd.n32788 vdd.n6638 0.002
R68814 vdd.n32793 vdd.n6580 0.002
R68815 vdd.n32799 vdd.n6524 0.002
R68816 vdd.n32804 vdd.n6470 0.002
R68817 vdd.n32809 vdd.n6408 0.002
R68818 vdd.n2535 vdd.n2530 0.002
R68819 vdd.n3904 vdd.n3903 0.002
R68820 vdd.n31374 vdd.n31372 0.002
R68821 vdd.n31305 vdd.n31304 0.002
R68822 vdd.n31347 vdd.n31341 0.002
R68823 vdd.n31400 vdd.n31394 0.002
R68824 vdd.n30915 vdd.n30909 0.002
R68825 vdd.n30720 vdd.n30714 0.002
R68826 vdd.n30173 vdd.n30167 0.002
R68827 vdd.n32593 vdd.n32587 0.002
R68828 vdd.n30155 vdd.n30149 0.002
R68829 vdd.n30068 vdd.n30062 0.002
R68830 vdd.n30035 vdd.n30029 0.002
R68831 vdd.n32634 vdd.n32628 0.002
R68832 vdd.n32731 vdd.n32725 0.002
R68833 vdd.n29610 vdd.n29604 0.002
R68834 vdd.n29561 vdd.n29555 0.002
R68835 vdd.n29491 vdd.n29486 0.002
R68836 vdd.n29405 vdd.n29400 0.002
R68837 vdd.n29367 vdd.n29361 0.002
R68838 vdd.n29266 vdd.n29261 0.002
R68839 vdd.n29248 vdd.n29243 0.002
R68840 vdd.n29144 vdd.n29139 0.002
R68841 vdd.n27743 vdd.n27738 0.002
R68842 vdd.n27704 vdd.n27698 0.002
R68843 vdd.n26534 vdd.n26528 0.002
R68844 vdd.n26557 vdd.n26552 0.002
R68845 vdd.n26267 vdd.n26261 0.002
R68846 vdd.n26578 vdd.n26572 0.002
R68847 vdd.n26226 vdd.n26220 0.002
R68848 vdd.n26092 vdd.n26086 0.002
R68849 vdd.n31326 vdd.n31321 0.002
R68850 vdd.n27251 vdd.n27248 0.002
R68851 vdd.n26092 vdd.n26085 0.002
R68852 vdd.n25354 vdd.n25348 0.002
R68853 vdd.n25354 vdd.n25346 0.002
R68854 vdd.n26226 vdd.n26218 0.002
R68855 vdd.n26718 vdd.n26715 0.002
R68856 vdd.n26718 vdd.n26713 0.002
R68857 vdd.n26578 vdd.n26570 0.002
R68858 vdd.n26250 vdd.n26245 0.002
R68859 vdd.n26250 vdd.n26243 0.002
R68860 vdd.n26267 vdd.n26259 0.002
R68861 vdd.n26415 vdd.n26411 0.002
R68862 vdd.n26415 vdd.n26409 0.002
R68863 vdd.n26557 vdd.n26551 0.002
R68864 vdd.n26438 vdd.n26433 0.002
R68865 vdd.n26438 vdd.n26431 0.002
R68866 vdd.n26534 vdd.n26526 0.002
R68867 vdd.n27681 vdd.n27677 0.002
R68868 vdd.n27681 vdd.n27675 0.002
R68869 vdd.n27704 vdd.n27697 0.002
R68870 vdd.n27723 vdd.n27719 0.002
R68871 vdd.n27723 vdd.n27717 0.002
R68872 vdd.n27743 vdd.n27737 0.002
R68873 vdd.n29110 vdd.n29105 0.002
R68874 vdd.n29110 vdd.n29103 0.002
R68875 vdd.n29144 vdd.n29137 0.002
R68876 vdd.n29172 vdd.n29169 0.002
R68877 vdd.n29172 vdd.n29167 0.002
R68878 vdd.n29248 vdd.n29242 0.002
R68879 vdd.n29214 vdd.n29210 0.002
R68880 vdd.n29214 vdd.n29208 0.002
R68881 vdd.n29266 vdd.n29260 0.002
R68882 vdd.n29346 vdd.n29340 0.002
R68883 vdd.n29346 vdd.n29338 0.002
R68884 vdd.n29367 vdd.n29360 0.002
R68885 vdd.n29389 vdd.n29384 0.002
R68886 vdd.n29389 vdd.n29382 0.002
R68887 vdd.n29405 vdd.n29399 0.002
R68888 vdd.n29472 vdd.n29468 0.002
R68889 vdd.n29472 vdd.n29466 0.002
R68890 vdd.n29491 vdd.n29484 0.002
R68891 vdd.n7218 vdd.n7215 0.002
R68892 vdd.n29561 vdd.n29554 0.002
R68893 vdd.n29588 vdd.n29582 0.002
R68894 vdd.n29588 vdd.n29580 0.002
R68895 vdd.n29610 vdd.n29602 0.002
R68896 vdd.n29628 vdd.n29625 0.002
R68897 vdd.n29628 vdd.n29623 0.002
R68898 vdd.n32731 vdd.n32723 0.002
R68899 vdd.n32711 vdd.n32707 0.002
R68900 vdd.n32711 vdd.n32705 0.002
R68901 vdd.n32634 vdd.n32626 0.002
R68902 vdd.n29679 vdd.n29675 0.002
R68903 vdd.n29679 vdd.n29673 0.002
R68904 vdd.n30035 vdd.n30027 0.002
R68905 vdd.n30004 vdd.n29999 0.002
R68906 vdd.n30004 vdd.n29997 0.002
R68907 vdd.n30068 vdd.n30060 0.002
R68908 vdd.n30133 vdd.n30129 0.002
R68909 vdd.n30133 vdd.n30127 0.002
R68910 vdd.n30155 vdd.n30147 0.002
R68911 vdd.n32613 vdd.n32609 0.002
R68912 vdd.n32613 vdd.n32607 0.002
R68913 vdd.n32593 vdd.n32585 0.002
R68914 vdd.n32571 vdd.n32567 0.002
R68915 vdd.n32571 vdd.n32565 0.002
R68916 vdd.n30173 vdd.n30166 0.002
R68917 vdd.n30869 vdd.n30864 0.002
R68918 vdd.n30869 vdd.n30862 0.002
R68919 vdd.n30720 vdd.n30713 0.002
R68920 vdd.n30892 vdd.n30887 0.002
R68921 vdd.n30892 vdd.n30885 0.002
R68922 vdd.n30915 vdd.n30907 0.002
R68923 vdd.n30936 vdd.n30931 0.002
R68924 vdd.n30936 vdd.n30929 0.002
R68925 vdd.n31400 vdd.n31392 0.002
R68926 vdd.n31364 vdd.n31360 0.002
R68927 vdd.n31364 vdd.n31358 0.002
R68928 vdd.n31347 vdd.n31339 0.002
R68929 vdd.n30984 vdd.n30980 0.002
R68930 vdd.n30984 vdd.n30982 0.002
R68931 vdd.n27245 vdd.n26729 0.002
R68932 vdd.n24554 vdd.n24549 0.002
R68933 vdd.n32016 vdd.n32014 0.002
R68934 vdd.n32359 vdd.n32357 0.002
R68935 vdd.n25673 vdd.n25672 0.002
R68936 vdd.n27251 vdd.n27247 0.002
R68937 vdd.n27251 vdd.n27250 0.002
R68938 vdd.n26092 vdd.n26088 0.002
R68939 vdd.n31391 vdd.n31369 0.002
R68940 vdd.n30860 vdd.n30837 0.002
R68941 vdd.n32563 vdd.n32544 0.002
R68942 vdd.n32563 vdd.n32541 0.002
R68943 vdd.n30125 vdd.n30112 0.002
R68944 vdd.n30125 vdd.n30110 0.002
R68945 vdd.n29995 vdd.n29979 0.002
R68946 vdd.n30059 vdd.n30046 0.002
R68947 vdd.n29671 vdd.n29651 0.002
R68948 vdd.n29671 vdd.n29648 0.002
R68949 vdd.n32703 vdd.n32685 0.002
R68950 vdd.n32703 vdd.n32683 0.002
R68951 vdd.n32721 vdd.n32716 0.002
R68952 vdd.n29552 vdd.n29537 0.002
R68953 vdd.n29464 vdd.n29445 0.002
R68954 vdd.n29464 vdd.n29442 0.002
R68955 vdd.n29336 vdd.n29319 0.002
R68956 vdd.n29336 vdd.n29317 0.002
R68957 vdd.n29206 vdd.n29189 0.002
R68958 vdd.n29258 vdd.n29257 0.002
R68959 vdd.n29165 vdd.n29159 0.002
R68960 vdd.n29240 vdd.n29234 0.002
R68961 vdd.n29101 vdd.n29049 0.002
R68962 vdd.n29136 vdd.n29123 0.002
R68963 vdd.n27735 vdd.n27729 0.002
R68964 vdd.n26429 vdd.n26428 0.002
R68965 vdd.n26524 vdd.n26484 0.002
R68966 vdd.n26407 vdd.n26361 0.002
R68967 vdd.n26407 vdd.n26358 0.002
R68968 vdd.n26711 vdd.n26629 0.002
R68969 vdd.n26711 vdd.n26627 0.002
R68970 vdd.n26217 vdd.n26112 0.002
R68971 vdd.n26711 vdd.n26632 0.002
R68972 vdd.n26407 vdd.n26366 0.002
R68973 vdd.n29464 vdd.n29450 0.002
R68974 vdd.n29671 vdd.n29657 0.002
R68975 vdd.n30125 vdd.n30115 0.002
R68976 vdd.n32563 vdd.n32549 0.002
R68977 vdd.n31319 vdd.n31318 0.002
R68978 vdd.n30975 vdd.n30973 0.002
R68979 vdd.n30860 vdd.n30846 0.002
R68980 vdd.n29995 vdd.n29984 0.002
R68981 vdd.n30059 vdd.n30050 0.002
R68982 vdd.n29552 vdd.n29541 0.002
R68983 vdd.n29240 vdd.n29230 0.002
R68984 vdd.n29206 vdd.n29195 0.002
R68985 vdd.n29136 vdd.n29127 0.002
R68986 vdd.n29165 vdd.n29156 0.002
R68987 vdd.n26083 vdd.n25674 0.002
R68988 vdd.n30831 vdd.n30822 0.002
R68989 vdd.n31441 vdd.n31437 0.002
R68990 vdd.n31428 vdd.n31422 0.002
R68991 vdd.n30104 vdd.n30095 0.002
R68992 vdd.n30059 vdd.n30051 0.002
R68993 vdd.n29973 vdd.n29969 0.002
R68994 vdd.n29641 vdd.n29637 0.002
R68995 vdd.n32678 vdd.n32672 0.002
R68996 vdd.n29513 vdd.n29507 0.002
R68997 vdd.n29552 vdd.n29543 0.002
R68998 vdd.n7185 vdd.n7181 0.002
R68999 vdd.n7185 vdd.n7182 0.002
R69000 vdd.n29432 vdd.n29426 0.002
R69001 vdd.n29311 vdd.n29302 0.002
R69002 vdd.n29281 vdd.n29277 0.002
R69003 vdd.n29240 vdd.n29228 0.002
R69004 vdd.n29136 vdd.n29128 0.002
R69005 vdd.n29097 vdd.n29072 0.002
R69006 vdd.n26467 vdd.n26461 0.002
R69007 vdd.n26524 vdd.n26493 0.002
R69008 vdd.n26391 vdd.n26385 0.002
R69009 vdd.n26320 vdd.n26280 0.002
R69010 vdd.n26673 vdd.n26651 0.002
R69011 vdd.n26217 vdd.n26104 0.002
R69012 vdd.n29165 vdd.n29149 0.002
R69013 vdd.n27245 vdd.n26726 0.002
R69014 vdd.n26181 vdd.n26130 0.002
R69015 vdd.n26181 vdd.n26145 0.002
R69016 vdd.n26217 vdd.n26097 0.002
R69017 vdd.n26711 vdd.n26640 0.002
R69018 vdd.n26673 vdd.n26646 0.002
R69019 vdd.n26665 vdd.n26664 0.002
R69020 vdd.n26320 vdd.n26285 0.002
R69021 vdd.n26407 vdd.n26378 0.002
R69022 vdd.n26391 vdd.n26381 0.002
R69023 vdd.n26520 vdd.n26504 0.002
R69024 vdd.n26524 vdd.n26502 0.002
R69025 vdd.n26472 vdd.n26445 0.002
R69026 vdd.n26467 vdd.n26465 0.002
R69027 vdd.n29093 vdd.n29078 0.002
R69028 vdd.n29097 vdd.n29077 0.002
R69029 vdd.n29101 vdd.n29063 0.002
R69030 vdd.n29136 vdd.n29135 0.002
R69031 vdd.n29240 vdd.n29222 0.002
R69032 vdd.n29206 vdd.n29204 0.002
R69033 vdd.n29281 vdd.n29280 0.002
R69034 vdd.n29336 vdd.n29334 0.002
R69035 vdd.n29311 vdd.n29309 0.002
R69036 vdd.n29294 vdd.n29293 0.002
R69037 vdd.n29432 vdd.n29431 0.002
R69038 vdd.n29464 vdd.n29462 0.002
R69039 vdd.n7185 vdd.n7184 0.002
R69040 vdd.n7173 vdd.n7171 0.002
R69041 vdd.n29552 vdd.n29550 0.002
R69042 vdd.n29530 vdd.n29528 0.002
R69043 vdd.n29513 vdd.n29512 0.002
R69044 vdd.n32664 vdd.n32663 0.002
R69045 vdd.n32678 vdd.n32677 0.002
R69046 vdd.n32703 vdd.n32701 0.002
R69047 vdd.n29641 vdd.n29640 0.002
R69048 vdd.n29671 vdd.n29669 0.002
R69049 vdd.n29973 vdd.n29972 0.002
R69050 vdd.n29995 vdd.n29994 0.002
R69051 vdd.n30059 vdd.n30058 0.002
R69052 vdd.n30125 vdd.n30123 0.002
R69053 vdd.n30104 vdd.n30102 0.002
R69054 vdd.n30087 vdd.n30086 0.002
R69055 vdd.n31428 vdd.n31427 0.002
R69056 vdd.n32563 vdd.n32561 0.002
R69057 vdd.n31441 vdd.n31440 0.002
R69058 vdd.n30860 vdd.n30858 0.002
R69059 vdd.n30831 vdd.n30829 0.002
R69060 vdd.n30813 vdd.n30812 0.002
R69061 vdd.n30767 vdd.n30765 0.002
R69062 vdd.n27245 vdd.n26728 0.002
R69063 vdd.n26181 vdd.n26142 0.002
R69064 vdd.n26181 vdd.n26143 0.002
R69065 vdd.n26217 vdd.n26102 0.002
R69066 vdd.n26217 vdd.n26100 0.002
R69067 vdd.n26711 vdd.n26636 0.002
R69068 vdd.n26711 vdd.n26638 0.002
R69069 vdd.n26673 vdd.n26649 0.002
R69070 vdd.n26673 vdd.n26648 0.002
R69071 vdd.n26665 vdd.n26662 0.002
R69072 vdd.n26665 vdd.n26663 0.002
R69073 vdd.n26320 vdd.n26282 0.002
R69074 vdd.n26320 vdd.n26283 0.002
R69075 vdd.n26407 vdd.n26372 0.002
R69076 vdd.n26407 vdd.n26374 0.002
R69077 vdd.n26391 vdd.n26384 0.002
R69078 vdd.n26391 vdd.n26383 0.002
R69079 vdd.n26520 vdd.n26507 0.002
R69080 vdd.n26520 vdd.n26505 0.002
R69081 vdd.n26524 vdd.n26496 0.002
R69082 vdd.n26524 vdd.n26498 0.002
R69083 vdd.n26472 vdd.n26448 0.002
R69084 vdd.n26472 vdd.n26447 0.002
R69085 vdd.n26467 vdd.n26462 0.002
R69086 vdd.n26467 vdd.n26464 0.002
R69087 vdd.n29093 vdd.n29082 0.002
R69088 vdd.n29093 vdd.n29080 0.002
R69089 vdd.n29097 vdd.n29074 0.002
R69090 vdd.n29097 vdd.n29075 0.002
R69091 vdd.n29101 vdd.n29058 0.002
R69092 vdd.n29101 vdd.n29060 0.002
R69093 vdd.n29136 vdd.n29130 0.002
R69094 vdd.n29136 vdd.n29132 0.002
R69095 vdd.n29165 vdd.n29153 0.002
R69096 vdd.n29165 vdd.n29151 0.002
R69097 vdd.n29240 vdd.n29226 0.002
R69098 vdd.n29240 vdd.n29224 0.002
R69099 vdd.n29206 vdd.n29200 0.002
R69100 vdd.n29206 vdd.n29202 0.002
R69101 vdd.n29281 vdd.n29278 0.002
R69102 vdd.n29281 vdd.n29279 0.002
R69103 vdd.n29336 vdd.n29329 0.002
R69104 vdd.n29336 vdd.n29331 0.002
R69105 vdd.n29311 vdd.n29304 0.002
R69106 vdd.n29311 vdd.n29306 0.002
R69107 vdd.n29294 vdd.n29291 0.002
R69108 vdd.n29294 vdd.n29292 0.002
R69109 vdd.n29432 vdd.n29428 0.002
R69110 vdd.n29432 vdd.n29429 0.002
R69111 vdd.n29464 vdd.n29456 0.002
R69112 vdd.n29464 vdd.n29458 0.002
R69113 vdd.n7185 vdd.n7183 0.002
R69114 vdd.n7173 vdd.n7167 0.002
R69115 vdd.n29552 vdd.n29545 0.002
R69116 vdd.n29552 vdd.n29547 0.002
R69117 vdd.n29530 vdd.n29524 0.002
R69118 vdd.n29530 vdd.n29526 0.002
R69119 vdd.n29513 vdd.n29508 0.002
R69120 vdd.n29513 vdd.n29510 0.002
R69121 vdd.n32664 vdd.n32661 0.002
R69122 vdd.n32664 vdd.n32662 0.002
R69123 vdd.n32678 vdd.n32674 0.002
R69124 vdd.n32678 vdd.n32675 0.002
R69125 vdd.n32703 vdd.n32696 0.002
R69126 vdd.n32703 vdd.n32698 0.002
R69127 vdd.n29641 vdd.n29638 0.002
R69128 vdd.n29641 vdd.n29639 0.002
R69129 vdd.n29671 vdd.n29663 0.002
R69130 vdd.n29671 vdd.n29665 0.002
R69131 vdd.n29973 vdd.n29970 0.002
R69132 vdd.n29973 vdd.n29971 0.002
R69133 vdd.n29995 vdd.n29988 0.002
R69134 vdd.n29995 vdd.n29990 0.002
R69135 vdd.n30059 vdd.n30053 0.002
R69136 vdd.n30059 vdd.n30055 0.002
R69137 vdd.n30125 vdd.n30119 0.002
R69138 vdd.n30125 vdd.n30121 0.002
R69139 vdd.n30104 vdd.n30097 0.002
R69140 vdd.n30104 vdd.n30099 0.002
R69141 vdd.n30087 vdd.n30084 0.002
R69142 vdd.n30087 vdd.n30085 0.002
R69143 vdd.n31428 vdd.n31424 0.002
R69144 vdd.n31428 vdd.n31425 0.002
R69145 vdd.n32563 vdd.n32555 0.002
R69146 vdd.n32563 vdd.n32557 0.002
R69147 vdd.n31441 vdd.n31438 0.002
R69148 vdd.n31441 vdd.n31439 0.002
R69149 vdd.n30860 vdd.n30852 0.002
R69150 vdd.n30860 vdd.n30854 0.002
R69151 vdd.n30831 vdd.n30824 0.002
R69152 vdd.n30831 vdd.n30826 0.002
R69153 vdd.n30813 vdd.n30792 0.002
R69154 vdd.n30813 vdd.n30802 0.002
R69155 vdd.n30767 vdd.n30758 0.002
R69156 vdd.n26711 vdd.n26634 0.002
R69157 vdd.n26407 vdd.n26369 0.002
R69158 vdd.n29101 vdd.n29053 0.002
R69159 vdd.n29101 vdd.n29055 0.002
R69160 vdd.n29165 vdd.n29154 0.002
R69161 vdd.n29206 vdd.n29198 0.002
R69162 vdd.n29336 vdd.n29323 0.002
R69163 vdd.n29336 vdd.n29326 0.002
R69164 vdd.n29464 vdd.n29453 0.002
R69165 vdd.n7173 vdd.n7164 0.002
R69166 vdd.n32703 vdd.n32689 0.002
R69167 vdd.n32703 vdd.n32693 0.002
R69168 vdd.n29671 vdd.n29660 0.002
R69169 vdd.n29995 vdd.n29985 0.002
R69170 vdd.n30125 vdd.n30117 0.002
R69171 vdd.n32563 vdd.n32552 0.002
R69172 vdd.n30860 vdd.n30849 0.002
R69173 vdd.n26083 vdd.n25365 0.002
R69174 vdd.n26217 vdd.n26110 0.002
R69175 vdd.n26524 vdd.n26488 0.002
R69176 vdd.n29101 vdd.n29050 0.002
R69177 vdd.n29136 vdd.n29125 0.002
R69178 vdd.n29165 vdd.n29157 0.002
R69179 vdd.n29240 vdd.n29232 0.002
R69180 vdd.n29206 vdd.n29193 0.002
R69181 vdd.n7173 vdd.n7159 0.002
R69182 vdd.n29552 vdd.n29540 0.002
R69183 vdd.n29995 vdd.n29980 0.002
R69184 vdd.n30059 vdd.n30048 0.002
R69185 vdd.n30860 vdd.n30841 0.002
R69186 vdd.n30975 vdd.n30940 0.002
R69187 vdd.n27251 vdd.n27249 0.002
R69188 vdd.n26092 vdd.n26090 0.002
R69189 vdd.n25354 vdd.n25352 0.002
R69190 vdd.n25354 vdd.n25350 0.002
R69191 vdd.n26226 vdd.n26224 0.002
R69192 vdd.n26226 vdd.n26222 0.002
R69193 vdd.n26718 vdd.n26717 0.002
R69194 vdd.n26718 vdd.n26716 0.002
R69195 vdd.n26578 vdd.n26576 0.002
R69196 vdd.n26578 vdd.n26574 0.002
R69197 vdd.n26250 vdd.n26248 0.002
R69198 vdd.n26250 vdd.n26247 0.002
R69199 vdd.n26267 vdd.n26265 0.002
R69200 vdd.n26267 vdd.n26263 0.002
R69201 vdd.n26415 vdd.n26413 0.002
R69202 vdd.n26415 vdd.n26412 0.002
R69203 vdd.n26557 vdd.n26556 0.002
R69204 vdd.n26557 vdd.n26554 0.002
R69205 vdd.n26438 vdd.n26436 0.002
R69206 vdd.n26438 vdd.n26434 0.002
R69207 vdd.n26534 vdd.n26532 0.002
R69208 vdd.n26534 vdd.n26530 0.002
R69209 vdd.n27681 vdd.n27679 0.002
R69210 vdd.n27681 vdd.n27678 0.002
R69211 vdd.n27704 vdd.n27702 0.002
R69212 vdd.n27704 vdd.n27700 0.002
R69213 vdd.n27723 vdd.n27722 0.002
R69214 vdd.n27723 vdd.n27720 0.002
R69215 vdd.n27743 vdd.n27742 0.002
R69216 vdd.n27743 vdd.n27740 0.002
R69217 vdd.n29110 vdd.n29109 0.002
R69218 vdd.n29110 vdd.n29107 0.002
R69219 vdd.n29144 vdd.n29143 0.002
R69220 vdd.n29144 vdd.n29141 0.002
R69221 vdd.n29172 vdd.n29171 0.002
R69222 vdd.n29172 vdd.n29170 0.002
R69223 vdd.n29248 vdd.n29247 0.002
R69224 vdd.n29248 vdd.n29245 0.002
R69225 vdd.n29214 vdd.n29213 0.002
R69226 vdd.n29214 vdd.n29211 0.002
R69227 vdd.n29266 vdd.n29265 0.002
R69228 vdd.n29266 vdd.n29263 0.002
R69229 vdd.n29346 vdd.n29344 0.002
R69230 vdd.n29346 vdd.n29342 0.002
R69231 vdd.n29367 vdd.n29365 0.002
R69232 vdd.n29367 vdd.n29363 0.002
R69233 vdd.n29389 vdd.n29388 0.002
R69234 vdd.n29389 vdd.n29386 0.002
R69235 vdd.n29405 vdd.n29404 0.002
R69236 vdd.n29405 vdd.n29402 0.002
R69237 vdd.n29472 vdd.n29471 0.002
R69238 vdd.n29472 vdd.n29469 0.002
R69239 vdd.n29491 vdd.n29490 0.002
R69240 vdd.n29491 vdd.n29488 0.002
R69241 vdd.n7218 vdd.n7216 0.002
R69242 vdd.n29561 vdd.n29559 0.002
R69243 vdd.n29561 vdd.n29557 0.002
R69244 vdd.n29588 vdd.n29586 0.002
R69245 vdd.n29588 vdd.n29584 0.002
R69246 vdd.n29610 vdd.n29608 0.002
R69247 vdd.n29610 vdd.n29606 0.002
R69248 vdd.n29628 vdd.n29627 0.002
R69249 vdd.n29628 vdd.n29626 0.002
R69250 vdd.n32731 vdd.n32729 0.002
R69251 vdd.n32731 vdd.n32727 0.002
R69252 vdd.n32711 vdd.n32709 0.002
R69253 vdd.n32711 vdd.n32708 0.002
R69254 vdd.n32634 vdd.n32632 0.002
R69255 vdd.n32634 vdd.n32630 0.002
R69256 vdd.n29679 vdd.n29677 0.002
R69257 vdd.n29679 vdd.n29676 0.002
R69258 vdd.n30035 vdd.n30033 0.002
R69259 vdd.n30035 vdd.n30031 0.002
R69260 vdd.n30004 vdd.n30002 0.002
R69261 vdd.n30004 vdd.n30001 0.002
R69262 vdd.n30068 vdd.n30066 0.002
R69263 vdd.n30068 vdd.n30064 0.002
R69264 vdd.n30133 vdd.n30131 0.002
R69265 vdd.n30133 vdd.n30130 0.002
R69266 vdd.n30155 vdd.n30153 0.002
R69267 vdd.n30155 vdd.n30151 0.002
R69268 vdd.n32613 vdd.n32611 0.002
R69269 vdd.n32613 vdd.n32610 0.002
R69270 vdd.n32593 vdd.n32591 0.002
R69271 vdd.n32593 vdd.n32589 0.002
R69272 vdd.n32571 vdd.n32569 0.002
R69273 vdd.n32571 vdd.n32568 0.002
R69274 vdd.n30173 vdd.n30171 0.002
R69275 vdd.n30173 vdd.n30169 0.002
R69276 vdd.n30869 vdd.n30867 0.002
R69277 vdd.n30869 vdd.n30865 0.002
R69278 vdd.n30720 vdd.n30718 0.002
R69279 vdd.n30720 vdd.n30716 0.002
R69280 vdd.n30892 vdd.n30890 0.002
R69281 vdd.n30892 vdd.n30888 0.002
R69282 vdd.n30915 vdd.n30913 0.002
R69283 vdd.n30915 vdd.n30911 0.002
R69284 vdd.n30936 vdd.n30934 0.002
R69285 vdd.n30936 vdd.n30933 0.002
R69286 vdd.n31400 vdd.n31398 0.002
R69287 vdd.n31400 vdd.n31396 0.002
R69288 vdd.n31364 vdd.n31362 0.002
R69289 vdd.n31364 vdd.n31361 0.002
R69290 vdd.n31347 vdd.n31345 0.002
R69291 vdd.n31347 vdd.n31343 0.002
R69292 vdd.n30984 vdd.n30978 0.002
R69293 vdd.n30984 vdd.n30977 0.002
R69294 vdd.n31326 vdd.n31324 0.002
R69295 vdd.n30813 vdd.n30733 0.002
R69296 vdd.n27245 vdd.n26722 0.002
R69297 vdd.n26181 vdd.n26118 0.002
R69298 vdd.n26217 vdd.n26115 0.002
R69299 vdd.n26711 vdd.n26625 0.002
R69300 vdd.n26673 vdd.n26656 0.002
R69301 vdd.n26665 vdd.n26659 0.002
R69302 vdd.n26320 vdd.n26273 0.002
R69303 vdd.n26407 vdd.n26355 0.002
R69304 vdd.n26391 vdd.n26389 0.002
R69305 vdd.n26520 vdd.n26516 0.002
R69306 vdd.n26524 vdd.n26479 0.002
R69307 vdd.n26472 vdd.n26454 0.002
R69308 vdd.n26467 vdd.n26456 0.002
R69309 vdd.n29093 vdd.n29090 0.002
R69310 vdd.n29097 vdd.n29066 0.002
R69311 vdd.n29101 vdd.n29047 0.002
R69312 vdd.n29136 vdd.n29121 0.002
R69313 vdd.n29165 vdd.n29162 0.002
R69314 vdd.n29240 vdd.n29236 0.002
R69315 vdd.n29206 vdd.n29182 0.002
R69316 vdd.n29281 vdd.n29274 0.002
R69317 vdd.n29336 vdd.n29273 0.002
R69318 vdd.n29311 vdd.n29285 0.002
R69319 vdd.n29294 vdd.n29287 0.002
R69320 vdd.n29432 vdd.n29417 0.002
R69321 vdd.n29464 vdd.n29413 0.002
R69322 vdd.n7185 vdd.n7178 0.002
R69323 vdd.n29552 vdd.n29498 0.002
R69324 vdd.n29530 vdd.n29499 0.002
R69325 vdd.n29513 vdd.n29501 0.002
R69326 vdd.n32664 vdd.n32651 0.002
R69327 vdd.n32678 vdd.n32648 0.002
R69328 vdd.n32703 vdd.n32641 0.002
R69329 vdd.n29641 vdd.n29635 0.002
R69330 vdd.n29671 vdd.n29633 0.002
R69331 vdd.n29973 vdd.n29962 0.002
R69332 vdd.n29995 vdd.n29959 0.002
R69333 vdd.n30059 vdd.n30041 0.002
R69334 vdd.n30125 vdd.n30075 0.002
R69335 vdd.n30104 vdd.n30078 0.002
R69336 vdd.n30087 vdd.n30080 0.002
R69337 vdd.n31428 vdd.n31413 0.002
R69338 vdd.n32563 vdd.n31410 0.002
R69339 vdd.n31441 vdd.n31432 0.002
R69340 vdd.n30860 vdd.n30727 0.002
R69341 vdd.n30831 vdd.n30729 0.002
R69342 vdd.n30813 vdd.n30730 0.002
R69343 vdd.n30767 vdd.n30734 0.002
R69344 vdd.n31225 vdd.n31191 0.002
R69345 vdd.n27710 vdd.n27709 0.002
R69346 vdd.n29616 vdd.n29615 0.002
R69347 vdd.n30921 vdd.n30920 0.002
R69348 vdd.n32077 vdd.n32056 0.002
R69349 vdd.n30962 vdd.n30961 0.002
R69350 vdd.n29948 vdd.n29947 0.001
R69351 vdd.n30584 vdd.n30583 0.001
R69352 vdd.n26133 vdd.n26132 0.001
R69353 vdd.n30966 vdd.n30965 0.001
R69354 vdd.n30740 vdd.n30737 0.001
R69355 vdd.n3887 vdd.n3803 0.001
R69356 vdd.n30944 vdd.n30943 0.001
R69357 vdd.n6404 vdd.n6402 0.001
R69358 vdd.n25272 vdd.n7901 0.001
R69359 vdd.n25278 vdd.n7844 0.001
R69360 vdd.n25284 vdd.n7787 0.001
R69361 vdd.n25288 vdd.n7730 0.001
R69362 vdd.n25293 vdd.n7673 0.001
R69363 vdd.n25298 vdd.n7616 0.001
R69364 vdd.n25303 vdd.n7558 0.001
R69365 vdd.n25309 vdd.n7501 0.001
R69366 vdd.n25315 vdd.n7447 0.001
R69367 vdd.n25320 vdd.n7390 0.001
R69368 vdd.n25326 vdd.n7332 0.001
R69369 vdd.n25332 vdd.n7278 0.001
R69370 vdd.n32737 vdd.n7220 0.001
R69371 vdd.n32742 vdd.n7109 0.001
R69372 vdd.n32748 vdd.n7054 0.001
R69373 vdd.n32754 vdd.n6998 0.001
R69374 vdd.n32760 vdd.n6941 0.001
R69375 vdd.n32766 vdd.n6884 0.001
R69376 vdd.n32772 vdd.n6829 0.001
R69377 vdd.n32778 vdd.n6770 0.001
R69378 vdd.n32782 vdd.n6713 0.001
R69379 vdd.n32788 vdd.n6659 0.001
R69380 vdd.n32793 vdd.n6600 0.001
R69381 vdd.n32799 vdd.n6546 0.001
R69382 vdd.n32804 vdd.n6488 0.001
R69383 vdd.n32809 vdd.n6433 0.001
R69384 vdd.n6404 vdd.n6401 0.001
R69385 vdd.n32739 vdd.n7147 0.001
R69386 vdd.n25298 vdd.n7608 0.001
R69387 vdd.n25296 vdd.n7636 0.001
R69388 vdd.n32751 vdd.n7017 0.001
R69389 vdd.n32748 vdd.n7045 0.001
R69390 vdd.n32745 vdd.n7071 0.001
R69391 vdd.n32788 vdd.n6650 0.001
R69392 vdd.n32799 vdd.n6538 0.001
R69393 vdd.n32796 vdd.n6566 0.001
R69394 vdd.n32812 vdd.n6385 0.001
R69395 vdd.n32809 vdd.n6426 0.001
R69396 vdd.n32809 vdd.n6424 0.001
R69397 vdd.n32807 vdd.n6456 0.001
R69398 vdd.n32807 vdd.n6454 0.001
R69399 vdd.n32804 vdd.n6481 0.001
R69400 vdd.n32804 vdd.n6480 0.001
R69401 vdd.n32802 vdd.n6511 0.001
R69402 vdd.n32802 vdd.n6509 0.001
R69403 vdd.n32799 vdd.n6540 0.001
R69404 vdd.n32799 vdd.n6536 0.001
R69405 vdd.n32796 vdd.n6568 0.001
R69406 vdd.n32796 vdd.n6564 0.001
R69407 vdd.n32793 vdd.n6594 0.001
R69408 vdd.n32793 vdd.n6592 0.001
R69409 vdd.n32790 vdd.n6624 0.001
R69410 vdd.n32790 vdd.n6622 0.001
R69411 vdd.n32788 vdd.n6651 0.001
R69412 vdd.n32788 vdd.n6649 0.001
R69413 vdd.n32785 vdd.n6684 0.001
R69414 vdd.n32785 vdd.n6682 0.001
R69415 vdd.n32782 vdd.n6706 0.001
R69416 vdd.n32782 vdd.n6705 0.001
R69417 vdd.n32780 vdd.n6735 0.001
R69418 vdd.n32780 vdd.n6733 0.001
R69419 vdd.n32778 vdd.n6763 0.001
R69420 vdd.n32778 vdd.n6761 0.001
R69421 vdd.n32775 vdd.n6795 0.001
R69422 vdd.n32775 vdd.n6793 0.001
R69423 vdd.n32772 vdd.n6823 0.001
R69424 vdd.n32772 vdd.n6821 0.001
R69425 vdd.n32769 vdd.n6850 0.001
R69426 vdd.n32769 vdd.n6848 0.001
R69427 vdd.n32766 vdd.n6879 0.001
R69428 vdd.n32766 vdd.n6877 0.001
R69429 vdd.n32763 vdd.n6906 0.001
R69430 vdd.n32763 vdd.n6904 0.001
R69431 vdd.n32760 vdd.n6935 0.001
R69432 vdd.n32760 vdd.n6933 0.001
R69433 vdd.n32757 vdd.n6963 0.001
R69434 vdd.n32757 vdd.n6961 0.001
R69435 vdd.n32754 vdd.n6992 0.001
R69436 vdd.n32754 vdd.n6990 0.001
R69437 vdd.n32751 vdd.n7019 0.001
R69438 vdd.n32751 vdd.n7016 0.001
R69439 vdd.n32748 vdd.n7047 0.001
R69440 vdd.n32748 vdd.n7043 0.001
R69441 vdd.n32745 vdd.n7073 0.001
R69442 vdd.n32745 vdd.n7069 0.001
R69443 vdd.n32742 vdd.n7103 0.001
R69444 vdd.n32742 vdd.n7101 0.001
R69445 vdd.n32739 vdd.n7136 0.001
R69446 vdd.n32739 vdd.n7134 0.001
R69447 vdd.n32737 vdd.n7202 0.001
R69448 vdd.n25335 vdd.n7242 0.001
R69449 vdd.n25335 vdd.n7240 0.001
R69450 vdd.n25332 vdd.n7271 0.001
R69451 vdd.n25332 vdd.n7270 0.001
R69452 vdd.n25329 vdd.n7300 0.001
R69453 vdd.n25329 vdd.n7298 0.001
R69454 vdd.n25326 vdd.n7326 0.001
R69455 vdd.n25326 vdd.n7325 0.001
R69456 vdd.n25323 vdd.n7354 0.001
R69457 vdd.n25323 vdd.n7352 0.001
R69458 vdd.n25320 vdd.n7383 0.001
R69459 vdd.n25320 vdd.n7382 0.001
R69460 vdd.n25318 vdd.n7411 0.001
R69461 vdd.n25318 vdd.n7409 0.001
R69462 vdd.n25315 vdd.n7440 0.001
R69463 vdd.n25315 vdd.n7439 0.001
R69464 vdd.n25312 vdd.n7467 0.001
R69465 vdd.n25312 vdd.n7465 0.001
R69466 vdd.n25309 vdd.n7492 0.001
R69467 vdd.n25309 vdd.n7490 0.001
R69468 vdd.n25306 vdd.n7524 0.001
R69469 vdd.n25306 vdd.n7522 0.001
R69470 vdd.n25303 vdd.n7552 0.001
R69471 vdd.n25303 vdd.n7551 0.001
R69472 vdd.n25301 vdd.n7580 0.001
R69473 vdd.n25301 vdd.n7578 0.001
R69474 vdd.n25298 vdd.n7609 0.001
R69475 vdd.n25298 vdd.n7607 0.001
R69476 vdd.n25296 vdd.n7638 0.001
R69477 vdd.n25296 vdd.n7634 0.001
R69478 vdd.n25293 vdd.n7666 0.001
R69479 vdd.n25293 vdd.n7665 0.001
R69480 vdd.n25291 vdd.n7695 0.001
R69481 vdd.n25291 vdd.n7693 0.001
R69482 vdd.n25288 vdd.n7723 0.001
R69483 vdd.n25288 vdd.n7722 0.001
R69484 vdd.n25286 vdd.n7750 0.001
R69485 vdd.n25286 vdd.n7748 0.001
R69486 vdd.n25284 vdd.n7780 0.001
R69487 vdd.n25284 vdd.n7779 0.001
R69488 vdd.n25281 vdd.n7810 0.001
R69489 vdd.n25281 vdd.n7808 0.001
R69490 vdd.n25278 vdd.n7838 0.001
R69491 vdd.n25278 vdd.n7837 0.001
R69492 vdd.n25275 vdd.n7866 0.001
R69493 vdd.n25275 vdd.n7864 0.001
R69494 vdd.n25272 vdd.n7894 0.001
R69495 vdd.n25272 vdd.n7893 0.001
R69496 vdd.n25269 vdd.n7922 0.001
R69497 vdd.n25269 vdd.n7920 0.001
R69498 vdd.n25266 vdd.n7951 0.001
R69499 vdd.n25266 vdd.n7950 0.001
R69500 vdd.n25264 vdd.n7970 0.001
R69501 vdd.n32812 vdd.n6383 0.001
R69502 vdd.n6372 vdd.n6367 0.001
R69503 vdd.n32812 vdd.n6384 0.001
R69504 vdd.n32812 vdd.n6378 0.001
R69505 vdd.n32809 vdd.n6422 0.001
R69506 vdd.n32807 vdd.n6452 0.001
R69507 vdd.n32807 vdd.n6451 0.001
R69508 vdd.n32804 vdd.n6479 0.001
R69509 vdd.n32802 vdd.n6508 0.001
R69510 vdd.n32802 vdd.n6506 0.001
R69511 vdd.n32796 vdd.n6563 0.001
R69512 vdd.n32793 vdd.n6591 0.001
R69513 vdd.n32790 vdd.n6620 0.001
R69514 vdd.n32790 vdd.n6617 0.001
R69515 vdd.n32785 vdd.n6680 0.001
R69516 vdd.n32785 vdd.n6677 0.001
R69517 vdd.n32782 vdd.n6704 0.001
R69518 vdd.n32780 vdd.n6731 0.001
R69519 vdd.n32780 vdd.n6728 0.001
R69520 vdd.n32778 vdd.n6760 0.001
R69521 vdd.n32775 vdd.n6792 0.001
R69522 vdd.n32775 vdd.n6790 0.001
R69523 vdd.n32772 vdd.n6820 0.001
R69524 vdd.n32769 vdd.n6847 0.001
R69525 vdd.n32769 vdd.n6845 0.001
R69526 vdd.n32766 vdd.n6876 0.001
R69527 vdd.n32763 vdd.n6903 0.001
R69528 vdd.n32763 vdd.n6901 0.001
R69529 vdd.n32760 vdd.n6932 0.001
R69530 vdd.n32757 vdd.n6960 0.001
R69531 vdd.n32757 vdd.n6958 0.001
R69532 vdd.n32754 vdd.n6988 0.001
R69533 vdd.n32751 vdd.n7015 0.001
R69534 vdd.n32745 vdd.n7068 0.001
R69535 vdd.n32742 vdd.n7099 0.001
R69536 vdd.n32739 vdd.n7131 0.001
R69537 vdd.n32739 vdd.n7129 0.001
R69538 vdd.n25335 vdd.n7238 0.001
R69539 vdd.n25335 vdd.n7236 0.001
R69540 vdd.n25332 vdd.n7268 0.001
R69541 vdd.n25329 vdd.n7296 0.001
R69542 vdd.n25329 vdd.n7294 0.001
R69543 vdd.n25326 vdd.n7323 0.001
R69544 vdd.n25323 vdd.n7350 0.001
R69545 vdd.n25323 vdd.n7348 0.001
R69546 vdd.n25320 vdd.n7380 0.001
R69547 vdd.n25318 vdd.n7407 0.001
R69548 vdd.n25318 vdd.n7405 0.001
R69549 vdd.n25315 vdd.n7437 0.001
R69550 vdd.n25312 vdd.n7464 0.001
R69551 vdd.n25312 vdd.n7462 0.001
R69552 vdd.n25309 vdd.n7489 0.001
R69553 vdd.n25306 vdd.n7521 0.001
R69554 vdd.n25306 vdd.n7518 0.001
R69555 vdd.n25303 vdd.n7549 0.001
R69556 vdd.n25301 vdd.n7576 0.001
R69557 vdd.n25301 vdd.n7574 0.001
R69558 vdd.n25296 vdd.n7632 0.001
R69559 vdd.n25293 vdd.n7663 0.001
R69560 vdd.n25291 vdd.n7691 0.001
R69561 vdd.n25291 vdd.n7689 0.001
R69562 vdd.n25288 vdd.n7720 0.001
R69563 vdd.n25286 vdd.n7747 0.001
R69564 vdd.n25286 vdd.n7745 0.001
R69565 vdd.n25284 vdd.n7777 0.001
R69566 vdd.n25281 vdd.n7806 0.001
R69567 vdd.n25281 vdd.n7804 0.001
R69568 vdd.n25278 vdd.n7835 0.001
R69569 vdd.n25275 vdd.n7862 0.001
R69570 vdd.n25275 vdd.n7860 0.001
R69571 vdd.n25272 vdd.n7891 0.001
R69572 vdd.n25269 vdd.n7918 0.001
R69573 vdd.n25269 vdd.n7916 0.001
R69574 vdd.n25266 vdd.n7947 0.001
R69575 vdd.n25266 vdd.n7946 0.001
R69576 vdd.n32812 vdd.n6380 0.001
R69577 vdd.n32812 vdd.n6381 0.001
R69578 vdd.n32809 vdd.n6417 0.001
R69579 vdd.n32809 vdd.n6419 0.001
R69580 vdd.n32807 vdd.n6447 0.001
R69581 vdd.n32807 vdd.n6449 0.001
R69582 vdd.n32804 vdd.n6475 0.001
R69583 vdd.n32804 vdd.n6477 0.001
R69584 vdd.n32802 vdd.n6504 0.001
R69585 vdd.n32802 vdd.n6505 0.001
R69586 vdd.n32799 vdd.n6532 0.001
R69587 vdd.n32799 vdd.n6534 0.001
R69588 vdd.n32796 vdd.n6561 0.001
R69589 vdd.n32796 vdd.n6562 0.001
R69590 vdd.n32793 vdd.n6587 0.001
R69591 vdd.n32793 vdd.n6589 0.001
R69592 vdd.n32790 vdd.n6613 0.001
R69593 vdd.n32790 vdd.n6615 0.001
R69594 vdd.n32788 vdd.n6646 0.001
R69595 vdd.n32788 vdd.n6648 0.001
R69596 vdd.n32785 vdd.n6673 0.001
R69597 vdd.n32785 vdd.n6675 0.001
R69598 vdd.n32782 vdd.n6701 0.001
R69599 vdd.n32782 vdd.n6703 0.001
R69600 vdd.n32780 vdd.n6726 0.001
R69601 vdd.n32780 vdd.n6727 0.001
R69602 vdd.n32778 vdd.n6756 0.001
R69603 vdd.n32778 vdd.n6758 0.001
R69604 vdd.n32775 vdd.n6787 0.001
R69605 vdd.n32775 vdd.n6788 0.001
R69606 vdd.n32772 vdd.n6815 0.001
R69607 vdd.n32772 vdd.n6817 0.001
R69608 vdd.n32769 vdd.n6843 0.001
R69609 vdd.n32769 vdd.n6844 0.001
R69610 vdd.n32766 vdd.n6871 0.001
R69611 vdd.n32766 vdd.n6873 0.001
R69612 vdd.n32763 vdd.n6898 0.001
R69613 vdd.n32763 vdd.n6900 0.001
R69614 vdd.n32760 vdd.n6927 0.001
R69615 vdd.n32760 vdd.n6929 0.001
R69616 vdd.n32757 vdd.n6955 0.001
R69617 vdd.n32757 vdd.n6956 0.001
R69618 vdd.n32754 vdd.n6983 0.001
R69619 vdd.n32754 vdd.n6985 0.001
R69620 vdd.n32751 vdd.n7012 0.001
R69621 vdd.n32751 vdd.n7014 0.001
R69622 vdd.n32748 vdd.n7039 0.001
R69623 vdd.n32748 vdd.n7041 0.001
R69624 vdd.n32745 vdd.n7066 0.001
R69625 vdd.n32745 vdd.n7067 0.001
R69626 vdd.n32742 vdd.n7095 0.001
R69627 vdd.n32742 vdd.n7097 0.001
R69628 vdd.n32739 vdd.n7123 0.001
R69629 vdd.n32739 vdd.n7126 0.001
R69630 vdd.n32737 vdd.n7198 0.001
R69631 vdd.n25335 vdd.n7232 0.001
R69632 vdd.n25335 vdd.n7234 0.001
R69633 vdd.n25332 vdd.n7265 0.001
R69634 vdd.n25332 vdd.n7267 0.001
R69635 vdd.n25329 vdd.n7290 0.001
R69636 vdd.n25329 vdd.n7292 0.001
R69637 vdd.n25326 vdd.n7320 0.001
R69638 vdd.n25326 vdd.n7322 0.001
R69639 vdd.n25323 vdd.n7344 0.001
R69640 vdd.n25323 vdd.n7346 0.001
R69641 vdd.n25320 vdd.n7377 0.001
R69642 vdd.n25320 vdd.n7379 0.001
R69643 vdd.n25318 vdd.n7402 0.001
R69644 vdd.n25318 vdd.n7403 0.001
R69645 vdd.n25315 vdd.n7434 0.001
R69646 vdd.n25315 vdd.n7436 0.001
R69647 vdd.n25312 vdd.n7459 0.001
R69648 vdd.n25312 vdd.n7460 0.001
R69649 vdd.n25309 vdd.n7485 0.001
R69650 vdd.n25309 vdd.n7487 0.001
R69651 vdd.n25306 vdd.n7514 0.001
R69652 vdd.n25306 vdd.n7516 0.001
R69653 vdd.n25303 vdd.n7545 0.001
R69654 vdd.n25303 vdd.n7547 0.001
R69655 vdd.n25301 vdd.n7570 0.001
R69656 vdd.n25301 vdd.n7572 0.001
R69657 vdd.n25298 vdd.n7603 0.001
R69658 vdd.n25298 vdd.n7605 0.001
R69659 vdd.n25296 vdd.n7628 0.001
R69660 vdd.n25296 vdd.n7630 0.001
R69661 vdd.n25293 vdd.n7660 0.001
R69662 vdd.n25293 vdd.n7662 0.001
R69663 vdd.n25291 vdd.n7685 0.001
R69664 vdd.n25291 vdd.n7687 0.001
R69665 vdd.n25288 vdd.n7717 0.001
R69666 vdd.n25288 vdd.n7719 0.001
R69667 vdd.n25286 vdd.n7742 0.001
R69668 vdd.n25286 vdd.n7743 0.001
R69669 vdd.n25284 vdd.n7773 0.001
R69670 vdd.n25284 vdd.n7775 0.001
R69671 vdd.n25281 vdd.n7800 0.001
R69672 vdd.n25281 vdd.n7802 0.001
R69673 vdd.n25278 vdd.n7832 0.001
R69674 vdd.n25278 vdd.n7834 0.001
R69675 vdd.n25275 vdd.n7856 0.001
R69676 vdd.n25275 vdd.n7858 0.001
R69677 vdd.n25272 vdd.n7888 0.001
R69678 vdd.n25272 vdd.n7890 0.001
R69679 vdd.n25269 vdd.n7913 0.001
R69680 vdd.n25269 vdd.n7914 0.001
R69681 vdd.n25266 vdd.n7943 0.001
R69682 vdd.n25264 vdd.n7967 0.001
R69683 vdd.n25264 vdd.n7966 0.001
R69684 vdd.n6372 vdd.n6368 0.001
R69685 vdd.n32812 vdd.n6377 0.001
R69686 vdd.n32809 vdd.n6415 0.001
R69687 vdd.n32809 vdd.n6413 0.001
R69688 vdd.n32807 vdd.n6444 0.001
R69689 vdd.n32804 vdd.n6474 0.001
R69690 vdd.n32804 vdd.n6473 0.001
R69691 vdd.n32802 vdd.n6501 0.001
R69692 vdd.n32799 vdd.n6530 0.001
R69693 vdd.n32799 vdd.n6528 0.001
R69694 vdd.n32796 vdd.n6558 0.001
R69695 vdd.n32793 vdd.n6585 0.001
R69696 vdd.n32793 vdd.n6583 0.001
R69697 vdd.n32790 vdd.n6610 0.001
R69698 vdd.n32788 vdd.n6645 0.001
R69699 vdd.n32788 vdd.n6644 0.001
R69700 vdd.n32785 vdd.n6671 0.001
R69701 vdd.n32782 vdd.n6700 0.001
R69702 vdd.n32782 vdd.n6699 0.001
R69703 vdd.n32780 vdd.n6724 0.001
R69704 vdd.n32778 vdd.n6754 0.001
R69705 vdd.n32778 vdd.n6752 0.001
R69706 vdd.n32775 vdd.n6784 0.001
R69707 vdd.n32772 vdd.n6814 0.001
R69708 vdd.n32772 vdd.n6812 0.001
R69709 vdd.n32769 vdd.n6841 0.001
R69710 vdd.n32766 vdd.n6869 0.001
R69711 vdd.n32766 vdd.n6867 0.001
R69712 vdd.n32763 vdd.n6896 0.001
R69713 vdd.n32760 vdd.n6925 0.001
R69714 vdd.n32760 vdd.n6924 0.001
R69715 vdd.n32757 vdd.n6953 0.001
R69716 vdd.n32754 vdd.n6982 0.001
R69717 vdd.n32754 vdd.n6980 0.001
R69718 vdd.n32751 vdd.n7010 0.001
R69719 vdd.n32748 vdd.n7037 0.001
R69720 vdd.n32748 vdd.n7036 0.001
R69721 vdd.n32745 vdd.n7064 0.001
R69722 vdd.n32742 vdd.n7093 0.001
R69723 vdd.n32742 vdd.n7091 0.001
R69724 vdd.n32739 vdd.n7121 0.001
R69725 vdd.n32737 vdd.n7192 0.001
R69726 vdd.n25335 vdd.n7230 0.001
R69727 vdd.n25332 vdd.n7264 0.001
R69728 vdd.n25332 vdd.n7263 0.001
R69729 vdd.n25329 vdd.n7288 0.001
R69730 vdd.n25326 vdd.n7319 0.001
R69731 vdd.n25326 vdd.n7318 0.001
R69732 vdd.n25323 vdd.n7342 0.001
R69733 vdd.n25320 vdd.n7376 0.001
R69734 vdd.n25320 vdd.n7375 0.001
R69735 vdd.n25318 vdd.n7400 0.001
R69736 vdd.n25315 vdd.n7433 0.001
R69737 vdd.n25315 vdd.n7431 0.001
R69738 vdd.n25312 vdd.n7457 0.001
R69739 vdd.n25309 vdd.n7484 0.001
R69740 vdd.n25309 vdd.n7482 0.001
R69741 vdd.n25306 vdd.n7512 0.001
R69742 vdd.n25303 vdd.n7544 0.001
R69743 vdd.n25303 vdd.n7543 0.001
R69744 vdd.n25301 vdd.n7568 0.001
R69745 vdd.n25298 vdd.n7602 0.001
R69746 vdd.n25298 vdd.n7601 0.001
R69747 vdd.n25296 vdd.n7626 0.001
R69748 vdd.n25293 vdd.n7659 0.001
R69749 vdd.n25293 vdd.n7658 0.001
R69750 vdd.n25291 vdd.n7683 0.001
R69751 vdd.n25288 vdd.n7716 0.001
R69752 vdd.n25288 vdd.n7715 0.001
R69753 vdd.n25286 vdd.n7740 0.001
R69754 vdd.n25284 vdd.n7772 0.001
R69755 vdd.n25284 vdd.n7770 0.001
R69756 vdd.n25281 vdd.n7798 0.001
R69757 vdd.n25278 vdd.n7831 0.001
R69758 vdd.n25278 vdd.n7830 0.001
R69759 vdd.n25275 vdd.n7854 0.001
R69760 vdd.n25272 vdd.n7887 0.001
R69761 vdd.n25272 vdd.n7886 0.001
R69762 vdd.n25269 vdd.n7911 0.001
R69763 vdd.n25266 vdd.n7945 0.001
R69764 vdd.n25266 vdd.n7941 0.001
R69765 vdd.n25266 vdd.n7956 0.001
R69766 vdd.n25266 vdd.n7960 0.001
R69767 vdd.n32812 vdd.n6395 0.001
R69768 vdd.n32812 vdd.n6393 0.001
R69769 vdd.n32809 vdd.n6431 0.001
R69770 vdd.n32807 vdd.n6462 0.001
R69771 vdd.n32807 vdd.n6460 0.001
R69772 vdd.n32804 vdd.n6486 0.001
R69773 vdd.n32802 vdd.n6516 0.001
R69774 vdd.n32802 vdd.n6515 0.001
R69775 vdd.n32799 vdd.n6544 0.001
R69776 vdd.n32796 vdd.n6573 0.001
R69777 vdd.n32796 vdd.n6572 0.001
R69778 vdd.n32793 vdd.n6598 0.001
R69779 vdd.n32790 vdd.n6630 0.001
R69780 vdd.n32790 vdd.n6629 0.001
R69781 vdd.n32788 vdd.n6657 0.001
R69782 vdd.n32785 vdd.n6688 0.001
R69783 vdd.n32785 vdd.n6687 0.001
R69784 vdd.n32782 vdd.n6712 0.001
R69785 vdd.n32780 vdd.n6739 0.001
R69786 vdd.n32780 vdd.n6737 0.001
R69787 vdd.n32778 vdd.n6768 0.001
R69788 vdd.n32775 vdd.n6801 0.001
R69789 vdd.n32775 vdd.n6799 0.001
R69790 vdd.n32772 vdd.n6827 0.001
R69791 vdd.n32769 vdd.n6855 0.001
R69792 vdd.n32769 vdd.n6854 0.001
R69793 vdd.n32766 vdd.n6883 0.001
R69794 vdd.n32763 vdd.n6910 0.001
R69795 vdd.n32763 vdd.n6909 0.001
R69796 vdd.n32760 vdd.n6939 0.001
R69797 vdd.n32757 vdd.n6969 0.001
R69798 vdd.n32757 vdd.n6967 0.001
R69799 vdd.n32754 vdd.n6996 0.001
R69800 vdd.n32751 vdd.n7025 0.001
R69801 vdd.n32751 vdd.n7023 0.001
R69802 vdd.n32748 vdd.n7052 0.001
R69803 vdd.n32745 vdd.n7078 0.001
R69804 vdd.n32745 vdd.n7077 0.001
R69805 vdd.n32742 vdd.n7108 0.001
R69806 vdd.n32739 vdd.n7144 0.001
R69807 vdd.n32739 vdd.n7143 0.001
R69808 vdd.n25335 vdd.n7247 0.001
R69809 vdd.n25335 vdd.n7245 0.001
R69810 vdd.n25332 vdd.n7277 0.001
R69811 vdd.n25329 vdd.n7304 0.001
R69812 vdd.n25329 vdd.n7303 0.001
R69813 vdd.n25326 vdd.n7331 0.001
R69814 vdd.n25323 vdd.n7360 0.001
R69815 vdd.n25323 vdd.n7358 0.001
R69816 vdd.n25320 vdd.n7388 0.001
R69817 vdd.n25318 vdd.n7416 0.001
R69818 vdd.n25318 vdd.n7415 0.001
R69819 vdd.n25315 vdd.n7445 0.001
R69820 vdd.n25312 vdd.n7470 0.001
R69821 vdd.n25312 vdd.n7469 0.001
R69822 vdd.n25309 vdd.n7499 0.001
R69823 vdd.n25306 vdd.n7529 0.001
R69824 vdd.n25306 vdd.n7528 0.001
R69825 vdd.n25303 vdd.n7556 0.001
R69826 vdd.n25301 vdd.n7586 0.001
R69827 vdd.n25301 vdd.n7584 0.001
R69828 vdd.n25298 vdd.n7614 0.001
R69829 vdd.n25296 vdd.n7643 0.001
R69830 vdd.n25296 vdd.n7642 0.001
R69831 vdd.n25293 vdd.n7671 0.001
R69832 vdd.n25291 vdd.n7700 0.001
R69833 vdd.n25291 vdd.n7699 0.001
R69834 vdd.n25288 vdd.n7728 0.001
R69835 vdd.n25286 vdd.n7755 0.001
R69836 vdd.n25286 vdd.n7754 0.001
R69837 vdd.n25284 vdd.n7785 0.001
R69838 vdd.n25281 vdd.n7815 0.001
R69839 vdd.n25281 vdd.n7814 0.001
R69840 vdd.n25278 vdd.n7842 0.001
R69841 vdd.n25275 vdd.n7872 0.001
R69842 vdd.n25275 vdd.n7870 0.001
R69843 vdd.n25272 vdd.n7899 0.001
R69844 vdd.n25269 vdd.n7927 0.001
R69845 vdd.n25269 vdd.n7926 0.001
R69846 vdd.n25264 vdd.n7976 0.001
R69847 vdd.n25264 vdd.n7977 0.001
R69848 vdd.n32812 vdd.n6399 0.001
R69849 vdd.n32812 vdd.n6400 0.001
R69850 vdd.n32809 vdd.n6434 0.001
R69851 vdd.n32809 vdd.n6436 0.001
R69852 vdd.n32807 vdd.n6464 0.001
R69853 vdd.n32807 vdd.n6465 0.001
R69854 vdd.n32804 vdd.n6491 0.001
R69855 vdd.n32804 vdd.n6493 0.001
R69856 vdd.n32802 vdd.n6518 0.001
R69857 vdd.n32802 vdd.n6520 0.001
R69858 vdd.n32799 vdd.n6549 0.001
R69859 vdd.n32799 vdd.n6551 0.001
R69860 vdd.n32796 vdd.n6575 0.001
R69861 vdd.n32796 vdd.n6577 0.001
R69862 vdd.n32793 vdd.n6602 0.001
R69863 vdd.n32793 vdd.n6604 0.001
R69864 vdd.n32790 vdd.n6633 0.001
R69865 vdd.n32790 vdd.n6634 0.001
R69866 vdd.n32788 vdd.n6661 0.001
R69867 vdd.n32788 vdd.n6663 0.001
R69868 vdd.n32785 vdd.n6691 0.001
R69869 vdd.n32785 vdd.n6692 0.001
R69870 vdd.n32782 vdd.n6714 0.001
R69871 vdd.n32782 vdd.n6716 0.001
R69872 vdd.n32780 vdd.n6742 0.001
R69873 vdd.n32780 vdd.n6743 0.001
R69874 vdd.n32778 vdd.n6773 0.001
R69875 vdd.n32778 vdd.n6775 0.001
R69876 vdd.n32775 vdd.n6803 0.001
R69877 vdd.n32775 vdd.n6805 0.001
R69878 vdd.n32772 vdd.n6832 0.001
R69879 vdd.n32772 vdd.n6834 0.001
R69880 vdd.n32769 vdd.n6857 0.001
R69881 vdd.n32769 vdd.n6859 0.001
R69882 vdd.n32766 vdd.n6887 0.001
R69883 vdd.n32766 vdd.n6889 0.001
R69884 vdd.n32763 vdd.n6913 0.001
R69885 vdd.n32763 vdd.n6915 0.001
R69886 vdd.n32760 vdd.n6944 0.001
R69887 vdd.n32760 vdd.n6946 0.001
R69888 vdd.n32757 vdd.n6971 0.001
R69889 vdd.n32757 vdd.n6972 0.001
R69890 vdd.n32754 vdd.n7001 0.001
R69891 vdd.n32754 vdd.n7003 0.001
R69892 vdd.n32751 vdd.n7027 0.001
R69893 vdd.n32751 vdd.n7028 0.001
R69894 vdd.n32748 vdd.n7057 0.001
R69895 vdd.n32748 vdd.n7059 0.001
R69896 vdd.n32745 vdd.n7080 0.001
R69897 vdd.n32745 vdd.n7082 0.001
R69898 vdd.n32742 vdd.n7111 0.001
R69899 vdd.n32742 vdd.n7113 0.001
R69900 vdd.n32739 vdd.n7149 0.001
R69901 vdd.n32737 vdd.n7225 0.001
R69902 vdd.n25335 vdd.n7251 0.001
R69903 vdd.n25335 vdd.n7253 0.001
R69904 vdd.n25332 vdd.n7279 0.001
R69905 vdd.n25332 vdd.n7281 0.001
R69906 vdd.n25329 vdd.n7308 0.001
R69907 vdd.n25329 vdd.n7310 0.001
R69908 vdd.n25326 vdd.n7333 0.001
R69909 vdd.n25326 vdd.n7335 0.001
R69910 vdd.n25323 vdd.n7364 0.001
R69911 vdd.n25323 vdd.n7366 0.001
R69912 vdd.n25320 vdd.n7391 0.001
R69913 vdd.n25320 vdd.n7393 0.001
R69914 vdd.n25318 vdd.n7419 0.001
R69915 vdd.n25318 vdd.n7421 0.001
R69916 vdd.n25315 vdd.n7448 0.001
R69917 vdd.n25315 vdd.n7450 0.001
R69918 vdd.n25312 vdd.n7472 0.001
R69919 vdd.n25312 vdd.n7473 0.001
R69920 vdd.n25309 vdd.n7503 0.001
R69921 vdd.n25309 vdd.n7505 0.001
R69922 vdd.n25306 vdd.n7532 0.001
R69923 vdd.n25306 vdd.n7534 0.001
R69924 vdd.n25303 vdd.n7559 0.001
R69925 vdd.n25303 vdd.n7561 0.001
R69926 vdd.n25301 vdd.n7589 0.001
R69927 vdd.n25301 vdd.n7591 0.001
R69928 vdd.n25298 vdd.n7617 0.001
R69929 vdd.n25298 vdd.n7619 0.001
R69930 vdd.n25296 vdd.n7646 0.001
R69931 vdd.n25296 vdd.n7648 0.001
R69932 vdd.n25293 vdd.n7674 0.001
R69933 vdd.n25293 vdd.n7676 0.001
R69934 vdd.n25291 vdd.n7703 0.001
R69935 vdd.n25291 vdd.n7705 0.001
R69936 vdd.n25288 vdd.n7731 0.001
R69937 vdd.n25288 vdd.n7733 0.001
R69938 vdd.n25286 vdd.n7758 0.001
R69939 vdd.n25286 vdd.n7760 0.001
R69940 vdd.n25284 vdd.n7788 0.001
R69941 vdd.n25284 vdd.n7790 0.001
R69942 vdd.n25281 vdd.n7818 0.001
R69943 vdd.n25281 vdd.n7820 0.001
R69944 vdd.n25278 vdd.n7845 0.001
R69945 vdd.n25278 vdd.n7847 0.001
R69946 vdd.n25275 vdd.n7875 0.001
R69947 vdd.n25275 vdd.n7877 0.001
R69948 vdd.n25272 vdd.n7902 0.001
R69949 vdd.n25272 vdd.n7904 0.001
R69950 vdd.n25269 vdd.n7930 0.001
R69951 vdd.n25269 vdd.n7931 0.001
R69952 vdd.n25266 vdd.n7958 0.001
R69953 vdd.n25266 vdd.n7957 0.001
R69954 vdd.n32812 vdd.n6375 0.001
R69955 vdd.n32809 vdd.n6411 0.001
R69956 vdd.n32807 vdd.n6441 0.001
R69957 vdd.n32804 vdd.n6471 0.001
R69958 vdd.n32802 vdd.n6498 0.001
R69959 vdd.n32799 vdd.n6525 0.001
R69960 vdd.n32796 vdd.n6555 0.001
R69961 vdd.n32793 vdd.n6581 0.001
R69962 vdd.n32790 vdd.n6608 0.001
R69963 vdd.n32788 vdd.n6641 0.001
R69964 vdd.n32785 vdd.n6669 0.001
R69965 vdd.n32782 vdd.n6697 0.001
R69966 vdd.n32780 vdd.n6722 0.001
R69967 vdd.n32778 vdd.n6750 0.001
R69968 vdd.n32775 vdd.n6781 0.001
R69969 vdd.n32772 vdd.n6809 0.001
R69970 vdd.n32769 vdd.n6838 0.001
R69971 vdd.n32766 vdd.n6864 0.001
R69972 vdd.n32763 vdd.n6894 0.001
R69973 vdd.n32760 vdd.n6920 0.001
R69974 vdd.n32757 vdd.n6950 0.001
R69975 vdd.n32754 vdd.n6976 0.001
R69976 vdd.n32751 vdd.n7007 0.001
R69977 vdd.n32748 vdd.n7032 0.001
R69978 vdd.n32745 vdd.n7062 0.001
R69979 vdd.n32742 vdd.n7088 0.001
R69980 vdd.n32739 vdd.n7118 0.001
R69981 vdd.n25335 vdd.n7228 0.001
R69982 vdd.n25332 vdd.n7259 0.001
R69983 vdd.n25329 vdd.n7286 0.001
R69984 vdd.n25326 vdd.n7315 0.001
R69985 vdd.n25323 vdd.n7340 0.001
R69986 vdd.n25320 vdd.n7372 0.001
R69987 vdd.n25318 vdd.n7398 0.001
R69988 vdd.n25315 vdd.n7428 0.001
R69989 vdd.n25312 vdd.n7455 0.001
R69990 vdd.n25309 vdd.n7479 0.001
R69991 vdd.n25306 vdd.n7510 0.001
R69992 vdd.n25303 vdd.n7540 0.001
R69993 vdd.n25301 vdd.n7566 0.001
R69994 vdd.n25298 vdd.n7598 0.001
R69995 vdd.n25296 vdd.n7624 0.001
R69996 vdd.n25293 vdd.n7655 0.001
R69997 vdd.n25291 vdd.n7681 0.001
R69998 vdd.n25288 vdd.n7712 0.001
R69999 vdd.n25286 vdd.n7738 0.001
R70000 vdd.n25284 vdd.n7767 0.001
R70001 vdd.n25281 vdd.n7796 0.001
R70002 vdd.n25278 vdd.n7827 0.001
R70003 vdd.n25275 vdd.n7852 0.001
R70004 vdd.n25272 vdd.n7883 0.001
R70005 vdd.n25269 vdd.n7909 0.001
R70006 vdd.n25266 vdd.n7937 0.001
R70007 vdd.n25266 vdd.n7939 0.001
R70008 vdd.n25264 vdd.n7963 0.001
R70009 vdd.n31203 vdd.n31202 0.001
R70010 vdd.n32014 vdd.n31609 0.001
R70011 vdd.n32357 vdd.n31468 0.001
R70012 vdd.n6372 vdd.n6366 0.001
R70013 vdd.n6372 vdd.n6371 0.001
R70014 vdd.n2530 vdd.n2529 0.001
R70015 vdd.n32737 vdd.n31305 0.001
R70016 vdd.n3880 vdd.n3879 0.001
R70017 vdd.n1887 vdd.n1886 0.001
R70018 vdd.n1839 vdd.n1837 0.001
R70019 vdd.n32004 vdd.n32002 0.001
R70020 vdd.n32331 vdd.n32329 0.001
R70021 vdd.n32348 vdd.n32346 0.001
R70022 vdd.n25254 vdd.n25253 0.001
R70023 vdd.n30786 vdd.n30785 0.001
R70024 vdd.n29520 vdd.n29519 0.001
R70025 vdd.n30745 vdd.n30744 0.001
R70026 vdd.n32655 vdd.n32654 0.001
R70027 vdd.n2548 vdd.n2547 0.001
R70028 vdd.n26458 vdd.n26457 0.001
R70029 vdd.n1827 vdd.n1826 0.001
R70030 vdd.n2250 vdd.n2249 0.001
R70031 vdd.n32739 vdd.n32738 0.001
R70032 vdd.n24932 vdd.n24931 0.001
R70033 vdd.n26141 vdd.n26140 0.001
R70034 vdd.n32807 vdd.n6468 0.001
R70035 vdd.n32802 vdd.n6522 0.001
R70036 vdd.n32796 vdd.n6578 0.001
R70037 vdd.n32790 vdd.n6636 0.001
R70038 vdd.n32785 vdd.n6693 0.001
R70039 vdd.n32780 vdd.n6746 0.001
R70040 vdd.n32775 vdd.n6806 0.001
R70041 vdd.n32769 vdd.n6860 0.001
R70042 vdd.n32763 vdd.n6916 0.001
R70043 vdd.n32757 vdd.n6973 0.001
R70044 vdd.n32751 vdd.n7029 0.001
R70045 vdd.n32745 vdd.n7083 0.001
R70046 vdd.n32739 vdd.n7151 0.001
R70047 vdd.n25335 vdd.n7255 0.001
R70048 vdd.n25329 vdd.n7312 0.001
R70049 vdd.n25323 vdd.n7368 0.001
R70050 vdd.n25318 vdd.n7424 0.001
R70051 vdd.n25312 vdd.n7475 0.001
R70052 vdd.n25306 vdd.n7536 0.001
R70053 vdd.n25301 vdd.n7594 0.001
R70054 vdd.n25296 vdd.n7651 0.001
R70055 vdd.n25291 vdd.n7708 0.001
R70056 vdd.n25286 vdd.n7763 0.001
R70057 vdd.n25281 vdd.n7822 0.001
R70058 vdd.n25275 vdd.n7879 0.001
R70059 vdd.n25269 vdd.n7933 0.001
R70060 vdd.n25272 vdd.n7898 0.001
R70061 vdd.n25278 vdd.n7841 0.001
R70062 vdd.n25284 vdd.n7784 0.001
R70063 vdd.n25288 vdd.n7727 0.001
R70064 vdd.n25293 vdd.n7670 0.001
R70065 vdd.n25298 vdd.n7613 0.001
R70066 vdd.n25303 vdd.n7555 0.001
R70067 vdd.n25309 vdd.n7497 0.001
R70068 vdd.n25315 vdd.n7444 0.001
R70069 vdd.n25320 vdd.n7387 0.001
R70070 vdd.n25326 vdd.n7330 0.001
R70071 vdd.n25332 vdd.n7276 0.001
R70072 vdd.n32737 vdd.n7209 0.001
R70073 vdd.n32742 vdd.n7107 0.001
R70074 vdd.n32748 vdd.n7050 0.001
R70075 vdd.n32754 vdd.n6994 0.001
R70076 vdd.n32760 vdd.n6938 0.001
R70077 vdd.n32766 vdd.n6882 0.001
R70078 vdd.n32772 vdd.n6826 0.001
R70079 vdd.n32778 vdd.n6766 0.001
R70080 vdd.n32782 vdd.n6710 0.001
R70081 vdd.n32788 vdd.n6655 0.001
R70082 vdd.n32793 vdd.n6597 0.001
R70083 vdd.n32799 vdd.n6543 0.001
R70084 vdd.n32804 vdd.n6484 0.001
R70085 vdd.n32809 vdd.n6429 0.001
R70086 vdd.n25266 vdd.n7954 0.001
R70087 vdd.n6405 vdd.n6404 0.001
R70088 vdd.n32812 vdd.n6397 0.001
R70089 vdd.n32809 vdd.n6437 0.001
R70090 vdd.n32807 vdd.n6463 0.001
R70091 vdd.n32804 vdd.n6494 0.001
R70092 vdd.n32802 vdd.n6517 0.001
R70093 vdd.n32799 vdd.n6552 0.001
R70094 vdd.n32796 vdd.n6574 0.001
R70095 vdd.n32793 vdd.n6605 0.001
R70096 vdd.n32790 vdd.n6632 0.001
R70097 vdd.n32788 vdd.n6665 0.001
R70098 vdd.n32785 vdd.n6690 0.001
R70099 vdd.n32782 vdd.n6717 0.001
R70100 vdd.n32780 vdd.n6740 0.001
R70101 vdd.n32778 vdd.n6777 0.001
R70102 vdd.n32775 vdd.n6802 0.001
R70103 vdd.n32772 vdd.n6835 0.001
R70104 vdd.n32769 vdd.n6856 0.001
R70105 vdd.n32766 vdd.n6890 0.001
R70106 vdd.n32763 vdd.n6911 0.001
R70107 vdd.n32760 vdd.n6947 0.001
R70108 vdd.n32757 vdd.n6970 0.001
R70109 vdd.n32754 vdd.n7004 0.001
R70110 vdd.n32751 vdd.n7026 0.001
R70111 vdd.n32748 vdd.n7060 0.001
R70112 vdd.n32745 vdd.n7079 0.001
R70113 vdd.n32742 vdd.n7114 0.001
R70114 vdd.n25335 vdd.n7249 0.001
R70115 vdd.n25332 vdd.n7282 0.001
R70116 vdd.n25329 vdd.n7306 0.001
R70117 vdd.n25326 vdd.n7336 0.001
R70118 vdd.n25323 vdd.n7362 0.001
R70119 vdd.n25320 vdd.n7394 0.001
R70120 vdd.n25318 vdd.n7418 0.001
R70121 vdd.n25315 vdd.n7451 0.001
R70122 vdd.n25312 vdd.n7471 0.001
R70123 vdd.n25309 vdd.n7506 0.001
R70124 vdd.n25306 vdd.n7531 0.001
R70125 vdd.n25303 vdd.n7562 0.001
R70126 vdd.n25301 vdd.n7588 0.001
R70127 vdd.n25298 vdd.n7620 0.001
R70128 vdd.n25296 vdd.n7645 0.001
R70129 vdd.n25293 vdd.n7677 0.001
R70130 vdd.n25291 vdd.n7702 0.001
R70131 vdd.n25288 vdd.n7734 0.001
R70132 vdd.n25286 vdd.n7757 0.001
R70133 vdd.n25284 vdd.n7792 0.001
R70134 vdd.n25281 vdd.n7817 0.001
R70135 vdd.n25278 vdd.n7848 0.001
R70136 vdd.n25275 vdd.n7874 0.001
R70137 vdd.n25272 vdd.n7905 0.001
R70138 vdd.n25269 vdd.n7929 0.001
R70139 vdd.n25266 vdd.n7961 0.001
R70140 vdd.n25264 vdd.n7980 0.001
R70141 vdd.n25269 vdd.n7924 0.001
R70142 vdd.n25275 vdd.n7868 0.001
R70143 vdd.n25281 vdd.n7812 0.001
R70144 vdd.n25286 vdd.n7752 0.001
R70145 vdd.n25291 vdd.n7697 0.001
R70146 vdd.n25296 vdd.n7640 0.001
R70147 vdd.n25301 vdd.n7582 0.001
R70148 vdd.n25306 vdd.n7526 0.001
R70149 vdd.n25312 vdd.n7468 0.001
R70150 vdd.n25318 vdd.n7413 0.001
R70151 vdd.n25323 vdd.n7356 0.001
R70152 vdd.n25329 vdd.n7302 0.001
R70153 vdd.n25335 vdd.n7244 0.001
R70154 vdd.n32745 vdd.n7074 0.001
R70155 vdd.n32751 vdd.n7020 0.001
R70156 vdd.n32757 vdd.n6964 0.001
R70157 vdd.n32763 vdd.n6907 0.001
R70158 vdd.n32769 vdd.n6851 0.001
R70159 vdd.n32775 vdd.n6796 0.001
R70160 vdd.n32780 vdd.n6736 0.001
R70161 vdd.n32785 vdd.n6686 0.001
R70162 vdd.n32790 vdd.n6626 0.001
R70163 vdd.n32796 vdd.n6569 0.001
R70164 vdd.n32802 vdd.n6512 0.001
R70165 vdd.n32807 vdd.n6458 0.001
R70166 vdd.n32812 vdd.n6387 0.001
R70167 vdd.n32812 vdd.n6390 0.001
R70168 vdd.n32809 vdd.n6427 0.001
R70169 vdd.n32804 vdd.n6482 0.001
R70170 vdd.n32799 vdd.n6541 0.001
R70171 vdd.n32793 vdd.n6595 0.001
R70172 vdd.n32788 vdd.n6652 0.001
R70173 vdd.n32782 vdd.n6708 0.001
R70174 vdd.n32778 vdd.n6765 0.001
R70175 vdd.n32772 vdd.n6824 0.001
R70176 vdd.n32766 vdd.n6880 0.001
R70177 vdd.n32760 vdd.n6937 0.001
R70178 vdd.n32754 vdd.n6993 0.001
R70179 vdd.n32748 vdd.n7048 0.001
R70180 vdd.n32742 vdd.n7104 0.001
R70181 vdd.n32739 vdd.n7140 0.001
R70182 vdd.n25332 vdd.n7273 0.001
R70183 vdd.n25326 vdd.n7328 0.001
R70184 vdd.n25320 vdd.n7384 0.001
R70185 vdd.n25315 vdd.n7441 0.001
R70186 vdd.n25309 vdd.n7494 0.001
R70187 vdd.n25303 vdd.n7553 0.001
R70188 vdd.n25298 vdd.n7610 0.001
R70189 vdd.n25293 vdd.n7667 0.001
R70190 vdd.n25288 vdd.n7724 0.001
R70191 vdd.n25284 vdd.n7781 0.001
R70192 vdd.n25278 vdd.n7839 0.001
R70193 vdd.n25272 vdd.n7895 0.001
R70194 vdd.n25266 vdd.n7952 0.001
R70195 vdd.n25264 vdd.n7974 0.001
R70196 vdd.n35617 vdd.n35616 0.001
R70197 vdd.n5777 vdd.n5776 0.001
R70198 vdd.n26126 vdd.n26125 0.001
R70199 vdd.n31391 vdd.n31390 0.001
R70200 vdd.n26123 vdd.n26122 0.001
R70201 vdd.n7219 vdd.n7218 0.001
R70202 vdd.n7177 vdd.n7173 0.001
R70203 vdd.n30578 vdd.n30577 0.001
R70204 vdd.n29725 vdd.n29714 0.001
R70205 vdd.n29424 vdd.n29423 0.001
R70206 vdd.n26278 vdd.n26277 0.001
R70207 vdd.n30807 vdd.n30805 0.001
R70208 vdd.n34345 vdd.n34233 0.001
R70209 vdd.n35024 vdd.n34875 0.001
R70210 vdd.n5771 vdd.n5622 0.001
R70211 vdd.n30960 vdd.n30959 0.001
R70212 vdd.n30948 vdd.n30947 0.001
R70213 vdd.n11681 vdd.n11680 0.001
R70214 vdd.n21762 vdd.n21761 0.001
R70215 vdd.n31211 vdd.n31207 0.001
R70216 vdd.n31214 vdd.n31200 0.001
R70217 vdd.n25264 vdd.n25263 0.001
R70218 vdd.n33451 vdd.n33448 0.001
R70219 vdd.n33379 vdd.n33377 0.001
R70220 vdd.n33389 vdd.n33387 0.001
R70221 vdd.n33379 vdd.n33378 0.001
R70222 vdd.n33389 vdd.n33388 0.001
R70223 vdd.n33360 vdd.n33357 0.001
R70224 vdd.n33305 vdd.n33304 0.001
R70225 vdd.n33312 vdd.n33311 0.001
R70226 vdd.n33695 vdd.n33692 0.001
R70227 vdd.n33691 vdd.n33689 0.001
R70228 vdd.n33628 vdd.n33627 0.001
R70229 vdd.n33636 vdd.n33635 0.001
R70230 vdd.n33778 vdd.n33774 0.001
R70231 vdd.n34337 vdd.n34334 0.001
R70232 vdd.n34230 vdd.n34227 0.001
R70233 vdd.n34226 vdd.n34224 0.001
R70234 vdd.n33931 vdd.n33930 0.001
R70235 vdd.n34071 vdd.n33973 0.001
R70236 vdd.n34054 vdd.n34051 0.001
R70237 vdd.n34056 vdd.n34054 0.001
R70238 vdd.n34060 vdd.n34057 0.001
R70239 vdd.n34023 vdd.n34022 0.001
R70240 vdd.n34025 vdd.n34024 0.001
R70241 vdd.n35603 vdd.n35600 0.001
R70242 vdd.n35423 vdd.n35421 0.001
R70243 vdd.n35423 vdd.n35422 0.001
R70244 vdd.n35215 vdd.n35212 0.001
R70245 vdd.n35217 vdd.n35215 0.001
R70246 vdd.n35221 vdd.n35218 0.001
R70247 vdd.n35185 vdd.n35184 0.001
R70248 vdd.n35187 vdd.n35186 0.001
R70249 vdd.n35351 vdd.n35348 0.001
R70250 vdd.n35347 vdd.n35345 0.001
R70251 vdd.n35015 vdd.n35012 0.001
R70252 vdd.n34767 vdd.n34764 0.001
R70253 vdd.n34763 vdd.n34761 0.001
R70254 vdd.n34827 vdd.n34825 0.001
R70255 vdd.n34827 vdd.n34826 0.001
R70256 vdd.n34646 vdd.n34545 0.001
R70257 vdd.n34628 vdd.n34625 0.001
R70258 vdd.n34630 vdd.n34628 0.001
R70259 vdd.n34634 vdd.n34631 0.001
R70260 vdd.n34594 vdd.n34593 0.001
R70261 vdd.n34609 vdd.n34608 0.001
R70262 vdd.n770 vdd.n767 0.001
R70263 vdd.n693 vdd.n691 0.001
R70264 vdd.n702 vdd.n700 0.001
R70265 vdd.n705 vdd.n704 0.001
R70266 vdd.n693 vdd.n692 0.001
R70267 vdd.n702 vdd.n701 0.001
R70268 vdd.n678 vdd.n675 0.001
R70269 vdd.n634 vdd.n633 0.001
R70270 vdd.n659 vdd.n658 0.001
R70271 vdd.n1161 vdd.n1158 0.001
R70272 vdd.n1157 vdd.n1155 0.001
R70273 vdd.n1085 vdd.n1084 0.001
R70274 vdd.n1130 vdd.n1129 0.001
R70275 vdd.n873 vdd.n869 0.001
R70276 vdd.n541 vdd.n540 0.001
R70277 vdd.n543 vdd.n542 0.001
R70278 vdd.n570 vdd.n567 0.001
R70279 vdd.n491 vdd.n489 0.001
R70280 vdd.n501 vdd.n499 0.001
R70281 vdd.n491 vdd.n490 0.001
R70282 vdd.n501 vdd.n500 0.001
R70283 vdd.n465 vdd.n462 0.001
R70284 vdd.n209 vdd.n208 0.001
R70285 vdd.n195 vdd.n192 0.001
R70286 vdd.n191 vdd.n189 0.001
R70287 vdd.n127 vdd.n126 0.001
R70288 vdd.n135 vdd.n134 0.001
R70289 vdd.n219 vdd.n215 0.001
R70290 vdd.n6038 vdd.n6035 0.001
R70291 vdd.n6214 vdd.n6203 0.001
R70292 vdd.n6215 vdd.n6214 0.001
R70293 vdd.n6339 vdd.n6336 0.001
R70294 vdd.n6341 vdd.n6339 0.001
R70295 vdd.n6345 vdd.n6342 0.001
R70296 vdd.n6305 vdd.n6304 0.001
R70297 vdd.n6320 vdd.n6319 0.001
R70298 vdd.n5857 vdd.n5854 0.001
R70299 vdd.n5853 vdd.n5851 0.001
R70300 vdd.n5762 vdd.n5759 0.001
R70301 vdd.n5514 vdd.n5511 0.001
R70302 vdd.n5510 vdd.n5508 0.001
R70303 vdd.n5574 vdd.n5572 0.001
R70304 vdd.n5574 vdd.n5573 0.001
R70305 vdd.n5393 vdd.n5291 0.001
R70306 vdd.n5375 vdd.n5372 0.001
R70307 vdd.n5377 vdd.n5375 0.001
R70308 vdd.n5381 vdd.n5378 0.001
R70309 vdd.n5341 vdd.n5340 0.001
R70310 vdd.n5356 vdd.n5355 0.001
R70311 vdd.n5107 vdd.n5106 0.001
R70312 vdd.n5115 vdd.n5114 0.001
R70313 vdd.n5175 vdd.n5172 0.001
R70314 vdd.n5171 vdd.n5169 0.001
R70315 vdd.n5169 vdd.n5166 0.001
R70316 vdd.n5011 vdd.n5010 0.001
R70317 vdd.n5010 vdd.n5009 0.001
R70318 vdd.n4702 vdd.n4699 0.001
R70319 vdd.n4945 vdd.n4942 0.001
R70320 vdd.n4941 vdd.n4939 0.001
R70321 vdd.n4592 vdd.n4589 0.001
R70322 vdd.n4341 vdd.n4338 0.001
R70323 vdd.n4337 vdd.n4335 0.001
R70324 vdd.n4400 vdd.n4398 0.001
R70325 vdd.n4400 vdd.n4399 0.001
R70326 vdd.n4205 vdd.n4202 0.001
R70327 vdd.n4207 vdd.n4205 0.001
R70328 vdd.n4211 vdd.n4208 0.001
R70329 vdd.n4172 vdd.n4171 0.001
R70330 vdd.n4187 vdd.n4186 0.001
R70331 vdd.n36978 vdd.n36975 0.001
R70332 vdd.n36986 vdd.n36981 0.001
R70333 vdd.n36992 vdd.n36989 0.001
R70334 vdd.n37000 vdd.n36995 0.001
R70335 vdd.n37009 vdd.n37007 0.001
R70336 vdd.n37014 vdd.n37011 0.001
R70337 vdd.n37024 vdd.n37022 0.001
R70338 vdd.n37029 vdd.n37026 0.001
R70339 vdd.n37034 vdd.n37032 0.001
R70340 vdd.n37062 vdd.n37048 0.001
R70341 vdd.n37076 vdd.n37075 0.001
R70342 vdd.n37075 vdd.n37072 0.001
R70343 vdd.n33252 vdd.n33251 0.001
R70344 vdd.n33251 vdd.n33240 0.001
R70345 vdd.n33240 vdd.n33237 0.001
R70346 vdd.n37098 vdd.n37088 0.001
R70347 vdd.n37085 vdd.n37083 0.001
R70348 vdd.n33225 vdd.n33223 0.001
R70349 vdd.n33221 vdd.n33211 0.001
R70350 vdd.n37119 vdd.n37118 0.001
R70351 vdd.n37118 vdd.n37116 0.001
R70352 vdd.n37114 vdd.n37107 0.001
R70353 vdd.n33200 vdd.n33198 0.001
R70354 vdd.n33185 vdd.n33177 0.001
R70355 vdd.n33162 vdd.n33161 0.001
R70356 vdd.n33161 vdd.n33159 0.001
R70357 vdd.n37168 vdd.n37166 0.001
R70358 vdd.n35633 vdd.n35631 0.001
R70359 vdd.n35629 vdd.n35627 0.001
R70360 vdd.n37187 vdd.n37185 0.001
R70361 vdd.n33139 vdd.n33138 0.001
R70362 vdd.n33138 vdd.n33128 0.001
R70363 vdd.n33126 vdd.n33124 0.001
R70364 vdd.n37207 vdd.n37197 0.001
R70365 vdd.n37221 vdd.n37213 0.001
R70366 vdd.n33098 vdd.n33096 0.001
R70367 vdd.n37239 vdd.n37238 0.001
R70368 vdd.n33087 vdd.n33084 0.001
R70369 vdd.n37261 vdd.n37250 0.001
R70370 vdd.n37250 vdd.n37247 0.001
R70371 vdd.n33060 vdd.n33050 0.001
R70372 vdd.n37285 vdd.n37284 0.001
R70373 vdd.n37284 vdd.n37282 0.001
R70374 vdd.n37280 vdd.n37270 0.001
R70375 vdd.n33029 vdd.n33026 0.001
R70376 vdd.n33040 vdd.n33038 0.001
R70377 vdd.n33014 vdd.n33007 0.001
R70378 vdd.n33019 vdd.n33014 0.001
R70379 vdd.n37314 vdd.n37307 0.001
R70380 vdd.n33004 vdd.n33003 0.001
R70381 vdd.n37339 vdd.n37337 0.001
R70382 vdd.n35650 vdd.n35648 0.001
R70383 vdd.n37363 vdd.n37361 0.001
R70384 vdd.n37375 vdd.n37370 0.001
R70385 vdd.n37389 vdd.n37379 0.001
R70386 vdd.n37398 vdd.n37395 0.001
R70387 vdd.n32943 vdd.n32941 0.001
R70388 vdd.n37425 vdd.n37423 0.001
R70389 vdd.n32937 vdd.n32931 0.001
R70390 vdd.n37456 vdd.n37453 0.001
R70391 vdd.n32915 vdd.n32905 0.001
R70392 vdd.n32905 vdd.n32902 0.001
R70393 vdd.n32889 vdd.n32886 0.001
R70394 vdd.n32893 vdd.n32891 0.001
R70395 vdd.n37488 vdd.n37483 0.001
R70396 vdd.n37494 vdd.n37491 0.001
R70397 vdd.n37497 vdd.n37494 0.001
R70398 vdd.n32874 vdd.n32869 0.001
R70399 vdd.n37510 vdd.n37503 0.001
R70400 vdd.n37515 vdd.n37510 0.001
R70401 vdd.n32850 vdd.n32840 0.001
R70402 vdd.n37538 vdd.n37529 0.001
R70403 vdd.n35660 vdd.n35658 0.001
R70404 vdd.n37551 vdd.n37550 0.001
R70405 vdd.n37562 vdd.n37557 0.001
R70406 vdd.n37579 vdd.n37576 0.001
R70407 vdd.n37587 vdd.n37582 0.001
R70408 vdd.n38215 vdd.n37587 0.001
R70409 vdd.n38214 vdd.n38204 0.001
R70410 vdd.n38202 vdd.n38200 0.001
R70411 vdd.n38197 vdd.n38190 0.001
R70412 vdd.n38188 vdd.n38186 0.001
R70413 vdd.n38176 vdd.n38174 0.001
R70414 vdd.n38159 vdd.n38157 0.001
R70415 vdd.n38157 vdd.n38155 0.001
R70416 vdd.n30636 vdd.n30209 0.001
R70417 vdd.n30692 vdd.n30690 0.001
R70418 vdd.n30698 vdd.n30697 0.001
R70419 vdd.n29767 vdd.n29751 0.001
R70420 vdd.n30008 vdd.n30007 0.001
R70421 vdd.n29943 vdd.n29873 0.001
R70422 vdd.n29904 vdd.n29887 0.001
R70423 vdd.n29882 vdd.n29878 0.001
R70424 vdd.n27890 vdd.n27886 0.001
R70425 vdd.n27941 vdd.n27940 0.001
R70426 vdd.n27957 vdd.n27884 0.001
R70427 vdd.n27988 vdd.n27976 0.001
R70428 vdd.n28027 vdd.n27824 0.001
R70429 vdd.n27754 vdd.n27753 0.001
R70430 vdd.n28976 vdd.n28972 0.001
R70431 vdd.n28068 vdd.n28067 0.001
R70432 vdd.n28934 vdd.n28068 0.001
R70433 vdd.n28097 vdd.n28093 0.001
R70434 vdd.n28919 vdd.n28099 0.001
R70435 vdd.n28918 vdd.n28917 0.001
R70436 vdd.n28865 vdd.n28120 0.001
R70437 vdd.n28104 vdd.n28103 0.001
R70438 vdd.n30201 vdd.n30196 0.001
R70439 vdd.n30603 vdd.n30263 0.001
R70440 vdd.n28838 vdd.n28837 0.001
R70441 vdd.n28846 vdd.n28843 0.001
R70442 vdd.n28903 vdd.n28900 0.001
R70443 vdd.n28916 vdd.n28913 0.001
R70444 vdd.n28941 vdd.n28938 0.001
R70445 vdd.n28953 vdd.n28950 0.001
R70446 vdd.n28991 vdd.n28958 0.001
R70447 vdd.n28037 vdd.n28035 0.001
R70448 vdd.n28013 vdd.n28010 0.001
R70449 vdd.n28006 vdd.n28005 0.001
R70450 vdd.n27997 vdd.n27996 0.001
R70451 vdd.n27961 vdd.n27959 0.001
R70452 vdd.n27953 vdd.n27951 0.001
R70453 vdd.n29898 vdd.n29895 0.001
R70454 vdd.n29904 vdd.n29903 0.001
R70455 vdd.n29911 vdd.n29908 0.001
R70456 vdd.n29810 vdd.n29805 0.001
R70457 vdd.n29741 vdd.n29738 0.001
R70458 vdd.n30649 vdd.n30647 0.001
R70459 vdd.n30640 vdd.n30638 0.001
R70460 vdd.n30629 vdd.n30628 0.001
R70461 vdd.n30628 vdd.n30627 0.001
R70462 vdd.n30621 vdd.n30620 0.001
R70463 vdd.n30619 vdd.n30617 0.001
R70464 vdd.n30610 vdd.n30608 0.001
R70465 vdd.n30594 vdd.n30593 0.001
R70466 vdd.n30593 vdd.n30592 0.001
R70467 vdd.n30588 vdd.n30587 0.001
R70468 vdd.n30587 vdd.n30584 0.001
R70469 vdd.n30575 vdd.n30571 0.001
R70470 vdd.n30570 vdd.n30569 0.001
R70471 vdd.n30553 vdd.n30550 0.001
R70472 vdd.n30550 vdd.n30549 0.001
R70473 vdd.n30549 vdd.n30548 0.001
R70474 vdd.n30535 vdd.n30533 0.001
R70475 vdd.n30521 vdd.n30519 0.001
R70476 vdd.n27606 vdd.n27603 0.001
R70477 vdd.n27601 vdd.n27600 0.001
R70478 vdd.n27463 vdd.n27460 0.001
R70479 vdd.n27357 vdd.n27354 0.001
R70480 vdd.n27353 vdd.n27352 0.001
R70481 vdd.n30989 vdd.n30988 0.001
R70482 vdd.n26022 vdd.n26019 0.001
R70483 vdd.n26017 vdd.n26016 0.001
R70484 vdd.n25909 vdd.n25906 0.001
R70485 vdd.n25809 vdd.n25806 0.001
R70486 vdd.n25805 vdd.n25804 0.001
R70487 vdd.n32737 vdd.n7207 0.001
R70488 vdd.n25607 vdd.n25604 0.001
R70489 vdd.n25530 vdd.n25526 0.001
R70490 vdd.n25492 vdd.n25489 0.001
R70491 vdd.n25488 vdd.n25485 0.001
R70492 vdd.n32599 vdd.n32598 0.001
R70493 vdd.n29374 vdd.n29373 0.001
R70494 vdd.n26235 vdd.n26234 0.001
R70495 vdd.n32737 vdd.n7204 0.001
R70496 vdd.n30797 vdd.n30793 0.001
R70497 vdd.n30987 vdd.n30986 0.001
R70498 vdd.n30801 vdd.n30800 0.001
R70499 vdd.n26139 vdd.n26138 0.001
R70500 vdd.n32737 vdd.n7201 0.001
R70501 vdd.n30810 vdd.n30808 0.001
R70502 vdd.n30995 vdd.n30994 0.001
R70503 vdd.n30996 vdd.n30995 0.001
R70504 vdd.n26665 vdd.n26661 0.001
R70505 vdd.n26520 vdd.n26511 0.001
R70506 vdd.n29097 vdd.n29070 0.001
R70507 vdd.n29281 vdd.n29276 0.001
R70508 vdd.n29294 vdd.n29290 0.001
R70509 vdd.n32678 vdd.n32670 0.001
R70510 vdd.n29973 vdd.n29967 0.001
R70511 vdd.n30087 vdd.n30083 0.001
R70512 vdd.n25344 vdd.n25343 0.001
R70513 vdd.n26568 vdd.n26566 0.001
R70514 vdd.n27715 vdd.n27714 0.001
R70515 vdd.n29359 vdd.n29356 0.001
R70516 vdd.n29621 vdd.n29620 0.001
R70517 vdd.n32624 vdd.n32622 0.001
R70518 vdd.n30145 vdd.n30142 0.001
R70519 vdd.n30927 vdd.n30925 0.001
R70520 vdd.n31356 vdd.n31353 0.001
R70521 vdd.n26092 vdd.n26083 0.001
R70522 vdd.n25360 vdd.n25359 0.001
R70523 vdd.n25354 vdd.n25344 0.001
R70524 vdd.n25339 vdd.n25338 0.001
R70525 vdd.n26226 vdd.n26217 0.001
R70526 vdd.n26094 vdd.n26093 0.001
R70527 vdd.n26718 vdd.n26711 0.001
R70528 vdd.n26584 vdd.n26583 0.001
R70529 vdd.n26578 vdd.n26568 0.001
R70530 vdd.n26561 vdd.n26560 0.001
R70531 vdd.n26250 vdd.n26241 0.001
R70532 vdd.n26231 vdd.n26230 0.001
R70533 vdd.n26267 vdd.n26258 0.001
R70534 vdd.n26252 vdd.n26251 0.001
R70535 vdd.n26415 vdd.n26407 0.001
R70536 vdd.n26270 vdd.n26269 0.001
R70537 vdd.n26557 vdd.n26549 0.001
R70538 vdd.n26540 vdd.n26539 0.001
R70539 vdd.n26438 vdd.n26429 0.001
R70540 vdd.n26419 vdd.n26418 0.001
R70541 vdd.n26534 vdd.n26524 0.001
R70542 vdd.n26442 vdd.n26441 0.001
R70543 vdd.n27681 vdd.n27673 0.001
R70544 vdd.n27664 vdd.n27663 0.001
R70545 vdd.n27704 vdd.n27695 0.001
R70546 vdd.n27685 vdd.n27684 0.001
R70547 vdd.n27723 vdd.n27715 0.001
R70548 vdd.n27708 vdd.n27707 0.001
R70549 vdd.n27743 vdd.n27735 0.001
R70550 vdd.n27727 vdd.n27726 0.001
R70551 vdd.n29110 vdd.n29101 0.001
R70552 vdd.n29042 vdd.n29041 0.001
R70553 vdd.n29144 vdd.n29136 0.001
R70554 vdd.n29116 vdd.n29115 0.001
R70555 vdd.n29172 vdd.n29165 0.001
R70556 vdd.n29147 vdd.n29146 0.001
R70557 vdd.n29248 vdd.n29240 0.001
R70558 vdd.n29219 vdd.n29218 0.001
R70559 vdd.n29214 vdd.n29206 0.001
R70560 vdd.n29179 vdd.n29178 0.001
R70561 vdd.n29266 vdd.n29258 0.001
R70562 vdd.n29253 vdd.n29252 0.001
R70563 vdd.n29346 vdd.n29336 0.001
R70564 vdd.n29270 vdd.n29269 0.001
R70565 vdd.n29367 vdd.n29359 0.001
R70566 vdd.n29351 vdd.n29350 0.001
R70567 vdd.n29389 vdd.n29380 0.001
R70568 vdd.n29371 vdd.n29370 0.001
R70569 vdd.n29405 vdd.n29398 0.001
R70570 vdd.n29472 vdd.n29464 0.001
R70571 vdd.n29491 vdd.n29481 0.001
R70572 vdd.n7206 vdd.n7205 0.001
R70573 vdd.n7213 vdd.n7212 0.001
R70574 vdd.n29561 vdd.n29552 0.001
R70575 vdd.n29497 vdd.n29496 0.001
R70576 vdd.n29588 vdd.n29578 0.001
R70577 vdd.n29569 vdd.n29568 0.001
R70578 vdd.n29610 vdd.n29601 0.001
R70579 vdd.n29592 vdd.n29591 0.001
R70580 vdd.n29628 vdd.n29621 0.001
R70581 vdd.n29614 vdd.n29613 0.001
R70582 vdd.n32731 vdd.n32721 0.001
R70583 vdd.n32714 vdd.n32713 0.001
R70584 vdd.n32711 vdd.n32703 0.001
R70585 vdd.n32638 vdd.n32637 0.001
R70586 vdd.n32634 vdd.n32624 0.001
R70587 vdd.n32620 vdd.n32619 0.001
R70588 vdd.n29679 vdd.n29671 0.001
R70589 vdd.n29630 vdd.n29629 0.001
R70590 vdd.n30035 vdd.n30025 0.001
R70591 vdd.n30017 vdd.n30016 0.001
R70592 vdd.n30004 vdd.n29995 0.001
R70593 vdd.n29956 vdd.n29955 0.001
R70594 vdd.n30068 vdd.n30059 0.001
R70595 vdd.n30039 vdd.n30038 0.001
R70596 vdd.n30133 vdd.n30125 0.001
R70597 vdd.n30072 vdd.n30071 0.001
R70598 vdd.n30155 vdd.n30145 0.001
R70599 vdd.n30137 vdd.n30136 0.001
R70600 vdd.n32613 vdd.n32605 0.001
R70601 vdd.n32596 vdd.n32595 0.001
R70602 vdd.n32593 vdd.n32583 0.001
R70603 vdd.n32575 vdd.n32574 0.001
R70604 vdd.n32571 vdd.n32563 0.001
R70605 vdd.n31407 vdd.n31406 0.001
R70606 vdd.n30173 vdd.n30164 0.001
R70607 vdd.n30157 vdd.n30156 0.001
R70608 vdd.n30869 vdd.n30860 0.001
R70609 vdd.n30724 vdd.n30723 0.001
R70610 vdd.n30720 vdd.n30711 0.001
R70611 vdd.n30702 vdd.n30701 0.001
R70612 vdd.n30892 vdd.n30883 0.001
R70613 vdd.n30873 vdd.n30872 0.001
R70614 vdd.n30915 vdd.n30905 0.001
R70615 vdd.n30936 vdd.n30927 0.001
R70616 vdd.n30919 vdd.n30918 0.001
R70617 vdd.n31400 vdd.n31391 0.001
R70618 vdd.n31367 vdd.n31366 0.001
R70619 vdd.n31364 vdd.n31356 0.001
R70620 vdd.n31351 vdd.n31350 0.001
R70621 vdd.n31347 vdd.n31337 0.001
R70622 vdd.n31331 vdd.n31330 0.001
R70623 vdd.n30984 vdd.n30975 0.001
R70624 vdd.n30938 vdd.n30937 0.001
R70625 vdd.n31326 vdd.n31319 0.001
R70626 vdd.n27660 vdd.n26092 0.001
R70627 vdd.n27660 vdd.n25354 0.001
R70628 vdd.n27660 vdd.n26226 0.001
R70629 vdd.n27660 vdd.n26718 0.001
R70630 vdd.n26580 vdd.n26579 0.001
R70631 vdd.n27660 vdd.n26578 0.001
R70632 vdd.n27660 vdd.n26250 0.001
R70633 vdd.n27660 vdd.n26267 0.001
R70634 vdd.n27660 vdd.n26415 0.001
R70635 vdd.n27660 vdd.n26557 0.001
R70636 vdd.n26440 vdd.n26439 0.001
R70637 vdd.n27660 vdd.n26438 0.001
R70638 vdd.n27660 vdd.n26534 0.001
R70639 vdd.n32737 vdd.n27681 0.001
R70640 vdd.n32737 vdd.n27704 0.001
R70641 vdd.n32737 vdd.n27723 0.001
R70642 vdd.n27745 vdd.n27744 0.001
R70643 vdd.n32737 vdd.n27743 0.001
R70644 vdd.n29112 vdd.n29111 0.001
R70645 vdd.n32737 vdd.n29110 0.001
R70646 vdd.n29114 vdd.n29113 0.001
R70647 vdd.n32737 vdd.n29144 0.001
R70648 vdd.n29174 vdd.n29173 0.001
R70649 vdd.n32737 vdd.n29172 0.001
R70650 vdd.n29217 vdd.n29216 0.001
R70651 vdd.n32737 vdd.n29248 0.001
R70652 vdd.n29177 vdd.n29176 0.001
R70653 vdd.n32737 vdd.n29214 0.001
R70654 vdd.n29251 vdd.n29250 0.001
R70655 vdd.n32737 vdd.n29266 0.001
R70656 vdd.n29348 vdd.n29347 0.001
R70657 vdd.n32737 vdd.n29346 0.001
R70658 vdd.n32737 vdd.n29367 0.001
R70659 vdd.n32737 vdd.n29389 0.001
R70660 vdd.n29407 vdd.n29406 0.001
R70661 vdd.n32737 vdd.n29405 0.001
R70662 vdd.n29409 vdd.n29408 0.001
R70663 vdd.n32737 vdd.n29472 0.001
R70664 vdd.n29493 vdd.n29492 0.001
R70665 vdd.n32737 vdd.n29491 0.001
R70666 vdd.n29565 vdd.n29564 0.001
R70667 vdd.n32737 vdd.n29561 0.001
R70668 vdd.n32737 vdd.n29588 0.001
R70669 vdd.n32737 vdd.n29610 0.001
R70670 vdd.n32737 vdd.n29628 0.001
R70671 vdd.n32733 vdd.n32732 0.001
R70672 vdd.n32737 vdd.n32731 0.001
R70673 vdd.n32737 vdd.n32711 0.001
R70674 vdd.n32737 vdd.n32634 0.001
R70675 vdd.n32737 vdd.n29679 0.001
R70676 vdd.n32737 vdd.n30035 0.001
R70677 vdd.n32737 vdd.n30004 0.001
R70678 vdd.n32737 vdd.n30068 0.001
R70679 vdd.n32737 vdd.n30133 0.001
R70680 vdd.n32737 vdd.n30155 0.001
R70681 vdd.n32737 vdd.n32613 0.001
R70682 vdd.n32737 vdd.n32593 0.001
R70683 vdd.n32737 vdd.n32571 0.001
R70684 vdd.n32737 vdd.n30173 0.001
R70685 vdd.n32737 vdd.n30869 0.001
R70686 vdd.n32737 vdd.n30720 0.001
R70687 vdd.n32737 vdd.n30892 0.001
R70688 vdd.n32737 vdd.n30915 0.001
R70689 vdd.n32737 vdd.n30936 0.001
R70690 vdd.n32737 vdd.n31400 0.001
R70691 vdd.n32737 vdd.n31364 0.001
R70692 vdd.n32737 vdd.n31347 0.001
R70693 vdd.n32737 vdd.n30984 0.001
R70694 vdd.n32737 vdd.n31326 0.001
R70695 vdd.n3680 vdd.n2713 0.001
R70696 vdd.n3982 vdd.n3762 0.001
R70697 vdd.n2602 vdd.n2594 0.001
R70698 vdd.n3679 vdd.n3676 0.001
R70699 vdd.n3682 vdd.n3681 0.001
R70700 vdd.n3684 vdd.n3683 0.001
R70701 vdd.n3694 vdd.n3693 0.001
R70702 vdd.n3700 vdd.n3695 0.001
R70703 vdd.n3703 vdd.n3700 0.001
R70704 vdd.n4016 vdd.n4015 0.001
R70705 vdd.n3999 vdd.n3998 0.001
R70706 vdd.n3984 vdd.n3983 0.001
R70707 vdd.n3974 vdd.n3972 0.001
R70708 vdd.n3963 vdd.n3961 0.001
R70709 vdd.n3940 vdd.n3938 0.001
R70710 vdd.n3924 vdd.n3921 0.001
R70711 vdd.n3916 vdd.n3914 0.001
R70712 vdd.n3891 vdd.n3889 0.001
R70713 vdd.n3866 vdd.n3865 0.001
R70714 vdd.n3861 vdd.n3859 0.001
R70715 vdd.n3859 vdd.n3858 0.001
R70716 vdd.n3855 vdd.n3846 0.001
R70717 vdd.n3841 vdd.n3837 0.001
R70718 vdd.n2233 vdd.n2228 0.001
R70719 vdd.n2256 vdd.n2253 0.001
R70720 vdd.n2259 vdd.n2258 0.001
R70721 vdd.n2261 vdd.n2260 0.001
R70722 vdd.n2267 vdd.n2266 0.001
R70723 vdd.n2273 vdd.n2268 0.001
R70724 vdd.n2276 vdd.n2273 0.001
R70725 vdd.n2297 vdd.n2294 0.001
R70726 vdd.n2317 vdd.n2316 0.001
R70727 vdd.n2336 vdd.n2335 0.001
R70728 vdd.n2352 vdd.n2349 0.001
R70729 vdd.n2367 vdd.n2364 0.001
R70730 vdd.n2556 vdd.n2554 0.001
R70731 vdd.n2544 vdd.n2542 0.001
R70732 vdd.n2518 vdd.n2516 0.001
R70733 vdd.n2511 vdd.n2506 0.001
R70734 vdd.n2501 vdd.n2500 0.001
R70735 vdd.n2486 vdd.n2484 0.001
R70736 vdd.n2484 vdd.n2483 0.001
R70737 vdd.n2480 vdd.n2472 0.001
R70738 vdd.n2467 vdd.n2463 0.001
R70739 vdd.n2616 vdd.n2611 0.001
R70740 vdd.n2648 vdd.n2645 0.001
R70741 vdd.n2659 vdd.n2658 0.001
R70742 vdd.n2661 vdd.n2660 0.001
R70743 vdd.n1962 vdd.n1961 0.001
R70744 vdd.n1970 vdd.n1967 0.001
R70745 vdd.n2084 vdd.n2083 0.001
R70746 vdd.n1952 vdd.n1951 0.001
R70747 vdd.n1946 vdd.n1944 0.001
R70748 vdd.n1919 vdd.n1917 0.001
R70749 vdd.n1893 vdd.n1892 0.001
R70750 vdd.n1889 vdd.n1888 0.001
R70751 vdd.n1888 vdd.n1887 0.001
R70752 vdd.n1872 vdd.n1866 0.001
R70753 vdd.n1866 vdd.n1861 0.001
R70754 vdd.n1858 vdd.n1856 0.001
R70755 vdd.n1854 vdd.n1851 0.001
R70756 vdd.n1846 vdd.n1845 0.001
R70757 vdd.n1843 vdd.n1841 0.001
R70758 vdd.n1807 vdd.n1805 0.001
R70759 vdd.n1805 vdd.n1802 0.001
R70760 vdd.n1799 vdd.n1791 0.001
R70761 vdd.n1786 vdd.n1784 0.001
R70762 vdd.n1775 vdd.n1774 0.001
R70763 vdd.n1799 vdd.n1261 0.001
R70764 vdd.n27241 vdd.n27229 0.001
R70765 vdd.n26193 vdd.n26190 0.001
R70766 vdd.n26595 vdd.n26591 0.001
R70767 vdd.n26620 vdd.n26601 0.001
R70768 vdd.n26612 vdd.n26609 0.001
R70769 vdd.n26609 vdd.n26608 0.001
R70770 vdd.n26686 vdd.n26683 0.001
R70771 vdd.n26337 vdd.n26330 0.001
R70772 vdd.n26336 vdd.n26334 0.001
R70773 vdd.n26349 vdd.n26348 0.001
R70774 vdd.n26348 vdd.n26343 0.001
R70775 vdd.n31785 vdd.n31767 0.001
R70776 vdd.n31794 vdd.n31791 0.001
R70777 vdd.n31805 vdd.n31804 0.001
R70778 vdd.n31814 vdd.n31811 0.001
R70779 vdd.n31826 vdd.n31825 0.001
R70780 vdd.n31851 vdd.n31850 0.001
R70781 vdd.n31905 vdd.n31900 0.001
R70782 vdd.n31907 vdd.n31906 0.001
R70783 vdd.n31936 vdd.n31916 0.001
R70784 vdd.n31938 vdd.n31937 0.001
R70785 vdd.n31950 vdd.n31942 0.001
R70786 vdd.n31973 vdd.n31972 0.001
R70787 vdd.n31988 vdd.n31986 0.001
R70788 vdd.n31996 vdd.n31994 0.001
R70789 vdd.n32007 vdd.n32004 0.001
R70790 vdd.n32031 vdd.n32024 0.001
R70791 vdd.n32040 vdd.n32037 0.001
R70792 vdd.n32053 vdd.n32050 0.001
R70793 vdd.n32107 vdd.n32106 0.001
R70794 vdd.n32133 vdd.n32117 0.001
R70795 vdd.n32134 vdd.n32133 0.001
R70796 vdd.n32144 vdd.n32141 0.001
R70797 vdd.n32172 vdd.n32169 0.001
R70798 vdd.n32187 vdd.n32186 0.001
R70799 vdd.n32206 vdd.n32205 0.001
R70800 vdd.n32245 vdd.n32236 0.001
R70801 vdd.n32270 vdd.n32265 0.001
R70802 vdd.n32277 vdd.n32270 0.001
R70803 vdd.n32279 vdd.n32278 0.001
R70804 vdd.n32296 vdd.n32288 0.001
R70805 vdd.n32298 vdd.n32297 0.001
R70806 vdd.n32306 vdd.n32303 0.001
R70807 vdd.n32356 vdd.n32354 0.001
R70808 vdd.n32362 vdd.n32359 0.001
R70809 vdd.n32533 vdd.n32531 0.001
R70810 vdd.n32517 vdd.n32515 0.001
R70811 vdd.n32511 vdd.n32507 0.001
R70812 vdd.n32507 vdd.n32502 0.001
R70813 vdd.n32502 vdd.n32500 0.001
R70814 vdd.n32486 vdd.n32480 0.001
R70815 vdd.n32480 vdd.n32478 0.001
R70816 vdd.n32461 vdd.n32459 0.001
R70817 vdd.n31058 vdd.n31055 0.001
R70818 vdd.n31073 vdd.n31072 0.001
R70819 vdd.n31099 vdd.n31098 0.001
R70820 vdd.n31187 vdd.n31124 0.001
R70821 vdd.n31981 vdd.n31980 0.001
R70822 vdd.n32087 vdd.n32086 0.001
R70823 vdd.n32243 vdd.n32242 0.001
R70824 vdd.n32323 vdd.n32322 0.001
R70825 vdd.n29206 vdd.n29187 0.001
R70826 vdd.n29283 vdd.n29282 0.001
R70827 vdd.n29311 vdd.n29297 0.001
R70828 vdd.n29295 vdd.n29294 0.001
R70829 vdd.n29435 vdd.n29434 0.001
R70830 vdd.n29438 vdd.n29437 0.001
R70831 vdd.n29552 vdd.n29535 0.001
R70832 vdd.n29517 vdd.n29516 0.001
R70833 vdd.n29516 vdd.n29515 0.001
R70834 vdd.n29515 vdd.n29514 0.001
R70835 vdd.n32665 vdd.n32664 0.001
R70836 vdd.n32678 vdd.n32667 0.001
R70837 vdd.n32643 vdd.n32642 0.001
R70838 vdd.n29643 vdd.n29642 0.001
R70839 vdd.n29671 vdd.n29646 0.001
R70840 vdd.n29973 vdd.n29963 0.001
R70841 vdd.n29974 vdd.n29973 0.001
R70842 vdd.n29995 vdd.n29976 0.001
R70843 vdd.n30104 vdd.n30090 0.001
R70844 vdd.n30088 vdd.n30087 0.001
R70845 vdd.n31431 vdd.n31430 0.001
R70846 vdd.n30860 vdd.n30834 0.001
R70847 vdd.n30832 vdd.n30831 0.001
R70848 vdd.n30779 vdd.n30778 0.001
R70849 vdd.n30767 vdd.n30743 0.001
R70850 vdd.n30741 vdd.n30740 0.001
R70851 vdd.n31228 vdd.n31227 0.001
R70852 vdd.n31238 vdd.n31237 0.001
R70853 vdd.n31248 vdd.n31247 0.001
R70854 vdd.n31302 vdd.n31290 0.001
R70855 vdd.n31303 vdd.n31302 0.001
R70856 vdd.n31236 vdd.n31235 0.001
R70857 vdd.n27245 vdd.n27244 0.001
R70858 vdd.n26162 vdd.n26157 0.001
R70859 vdd.n26163 vdd.n26162 0.001
R70860 vdd.n26181 vdd.n26180 0.001
R70861 vdd.n26673 vdd.n26672 0.001
R70862 vdd.n26670 vdd.n26665 0.001
R70863 vdd.n26351 vdd.n26322 0.001
R70864 vdd.n26406 vdd.n26405 0.001
R70865 vdd.n26520 vdd.n26519 0.001
R70866 vdd.n26524 vdd.n26523 0.001
R70867 vdd.n26471 vdd.n26470 0.001
R70868 vdd.n26470 vdd.n26469 0.001
R70869 vdd.n26469 vdd.n26468 0.001
R70870 vdd.n29094 vdd.n29093 0.001
R70871 vdd.n29097 vdd.n29096 0.001
R70872 vdd.n29118 vdd.n29117 0.001
R70873 vdd.n29165 vdd.n29164 0.001
R70874 vdd.n29240 vdd.n29238 0.001
R70875 vdd.n29240 vdd.n29239 0.001
R70876 vdd.n12572 vdd.n10257 0.001
R70877 vdd.n10601 vdd.n10589 0.001
R70878 vdd.n12478 vdd.n12477 0.001
R70879 vdd.n12377 vdd.n12376 0.001
R70880 vdd.n12375 vdd.n10752 0.001
R70881 vdd.n10945 vdd.n10944 0.001
R70882 vdd.n10948 vdd.n10946 0.001
R70883 vdd.n11091 vdd.n11089 0.001
R70884 vdd.n11113 vdd.n11111 0.001
R70885 vdd.n12078 vdd.n12077 0.001
R70886 vdd.n11293 vdd.n11267 0.001
R70887 vdd.n11497 vdd.n11464 0.001
R70888 vdd.n11521 vdd.n11460 0.001
R70889 vdd.n11538 vdd.n11453 0.001
R70890 vdd.n11941 vdd.n11553 0.001
R70891 vdd.n11939 vdd.n11554 0.001
R70892 vdd.n13860 vdd.n8704 0.001
R70893 vdd.n14102 vdd.n8495 0.001
R70894 vdd.n14149 vdd.n8481 0.001
R70895 vdd.n14412 vdd.n8292 0.001
R70896 vdd.n14415 vdd.n8266 0.001
R70897 vdd.n13815 vdd.n8717 0.001
R70898 vdd.n9197 vdd.n9183 0.001
R70899 vdd.n13281 vdd.n13280 0.001
R70900 vdd.n8975 vdd.n8962 0.001
R70901 vdd.n13573 vdd.n13572 0.001
R70902 vdd.n12600 vdd.n10082 0.001
R70903 vdd.n10449 vdd.n10448 0.001
R70904 vdd.n10302 vdd.n10293 0.001
R70905 vdd.n9349 vdd.n9334 0.001
R70906 vdd.n13038 vdd.n13037 0.001
R70907 vdd.n12941 vdd.n12940 0.001
R70908 vdd.n9534 vdd.n9533 0.001
R70909 vdd.n9709 vdd.n9694 0.001
R70910 vdd.n12830 vdd.n12829 0.001
R70911 vdd.n12733 vdd.n12732 0.001
R70912 vdd.n9895 vdd.n9894 0.001
R70913 vdd.n10162 vdd.n10147 0.001
R70914 vdd.n12621 vdd.n12620 0.001
R70915 vdd.n11686 vdd.n11682 0.001
R70916 vdd.n11869 vdd.n11809 0.001
R70917 vdd.n11919 vdd.n9284 0.001
R70918 vdd.n13182 vdd.n13181 0.001
R70919 vdd.n13210 vdd.n9205 0.001
R70920 vdd.n13251 vdd.n9176 0.001
R70921 vdd.n13272 vdd.n13271 0.001
R70922 vdd.n13298 vdd.n13297 0.001
R70923 vdd.n13297 vdd.n13296 0.001
R70924 vdd.n13342 vdd.n13341 0.001
R70925 vdd.n13415 vdd.n9039 0.001
R70926 vdd.n13419 vdd.n13418 0.001
R70927 vdd.n13418 vdd.n8998 0.001
R70928 vdd.n13487 vdd.n13486 0.001
R70929 vdd.n13476 vdd.n8985 0.001
R70930 vdd.n13564 vdd.n13563 0.001
R70931 vdd.n13584 vdd.n8926 0.001
R70932 vdd.n13590 vdd.n13589 0.001
R70933 vdd.n13589 vdd.n13588 0.001
R70934 vdd.n13634 vdd.n13633 0.001
R70935 vdd.n13691 vdd.n13690 0.001
R70936 vdd.n13709 vdd.n8818 0.001
R70937 vdd.n13712 vdd.n13711 0.001
R70938 vdd.n13711 vdd.n8781 0.001
R70939 vdd.n13767 vdd.n13766 0.001
R70940 vdd.n13756 vdd.n8770 0.001
R70941 vdd.n13846 vdd.n13845 0.001
R70942 vdd.n13852 vdd.n13847 0.001
R70943 vdd.n13894 vdd.n13893 0.001
R70944 vdd.n13893 vdd.n13892 0.001
R70945 vdd.n13909 vdd.n8673 0.001
R70946 vdd.n8670 vdd.n8669 0.001
R70947 vdd.n13986 vdd.n13985 0.001
R70948 vdd.n14058 vdd.n14057 0.001
R70949 vdd.n14057 vdd.n14056 0.001
R70950 vdd.n14046 vdd.n14045 0.001
R70951 vdd.n14074 vdd.n8556 0.001
R70952 vdd.n14135 vdd.n14134 0.001
R70953 vdd.n14141 vdd.n14136 0.001
R70954 vdd.n14183 vdd.n14182 0.001
R70955 vdd.n14182 vdd.n14181 0.001
R70956 vdd.n14199 vdd.n8449 0.001
R70957 vdd.n14276 vdd.n14275 0.001
R70958 vdd.n14333 vdd.n14332 0.001
R70959 vdd.n14332 vdd.n14331 0.001
R70960 vdd.n14351 vdd.n14350 0.001
R70961 vdd.n14352 vdd.n8300 0.001
R70962 vdd.n14425 vdd.n14424 0.001
R70963 vdd.n8280 vdd.n8246 0.001
R70964 vdd.n14652 vdd.n14651 0.001
R70965 vdd.n14690 vdd.n14689 0.001
R70966 vdd.n14719 vdd.n8110 0.001
R70967 vdd.n14766 vdd.n14765 0.001
R70968 vdd.n14767 vdd.n8068 0.001
R70969 vdd.n8062 vdd.n8060 0.001
R70970 vdd.n14824 vdd.n14823 0.001
R70971 vdd.n14864 vdd.n14863 0.001
R70972 vdd.n14901 vdd.n14900 0.001
R70973 vdd.n14937 vdd.n7982 0.001
R70974 vdd.n22323 vdd.n22322 0.001
R70975 vdd.n24327 vdd.n24324 0.001
R70976 vdd.n24295 vdd.n24294 0.001
R70977 vdd.n24210 vdd.n24207 0.001
R70978 vdd.n24202 vdd.n24192 0.001
R70979 vdd.n23982 vdd.n23980 0.001
R70980 vdd.n23970 vdd.n23960 0.001
R70981 vdd.n23750 vdd.n23748 0.001
R70982 vdd.n23738 vdd.n23728 0.001
R70983 vdd.n23062 vdd.n23060 0.001
R70984 vdd.n23282 vdd.n23272 0.001
R70985 vdd.n23294 vdd.n23292 0.001
R70986 vdd.n23514 vdd.n23504 0.001
R70987 vdd.n23526 vdd.n23524 0.001
R70988 vdd.n22483 vdd.n22481 0.001
R70989 vdd.n22703 vdd.n22693 0.001
R70990 vdd.n22715 vdd.n22713 0.001
R70991 vdd.n22935 vdd.n22925 0.001
R70992 vdd.n22947 vdd.n22945 0.001
R70993 vdd.n22467 vdd.n22466 0.001
R70994 vdd.n22382 vdd.n22379 0.001
R70995 vdd.n15122 vdd.n15120 0.001
R70996 vdd.n16981 vdd.n16980 0.001
R70997 vdd.n16996 vdd.n16982 0.001
R70998 vdd.n17253 vdd.n17252 0.001
R70999 vdd.n17268 vdd.n17254 0.001
R71000 vdd.n17525 vdd.n17524 0.001
R71001 vdd.n17540 vdd.n17526 0.001
R71002 vdd.n17783 vdd.n17782 0.001
R71003 vdd.n17798 vdd.n17784 0.001
R71004 vdd.n18054 vdd.n18053 0.001
R71005 vdd.n18069 vdd.n18055 0.001
R71006 vdd.n18316 vdd.n18315 0.001
R71007 vdd.n18349 vdd.n18348 0.001
R71008 vdd.n18376 vdd.n18373 0.001
R71009 vdd.n18392 vdd.n18391 0.001
R71010 vdd.n18404 vdd.n18403 0.001
R71011 vdd.n19140 vdd.n19134 0.001
R71012 vdd.n18908 vdd.n18906 0.001
R71013 vdd.n18888 vdd.n18876 0.001
R71014 vdd.n18649 vdd.n18647 0.001
R71015 vdd.n18629 vdd.n18617 0.001
R71016 vdd.n21017 vdd.n21015 0.001
R71017 vdd.n21533 vdd.n21531 0.001
R71018 vdd.n21513 vdd.n21501 0.001
R71019 vdd.n21274 vdd.n21272 0.001
R71020 vdd.n21254 vdd.n21242 0.001
R71021 vdd.n16743 vdd.n16717 0.001
R71022 vdd.n15309 vdd.n15308 0.001
R71023 vdd.n15328 vdd.n15314 0.001
R71024 vdd.n15537 vdd.n15536 0.001
R71025 vdd.n15562 vdd.n15542 0.001
R71026 vdd.n15793 vdd.n15792 0.001
R71027 vdd.n15818 vdd.n15798 0.001
R71028 vdd.n16049 vdd.n16048 0.001
R71029 vdd.n16074 vdd.n16054 0.001
R71030 vdd.n16305 vdd.n16304 0.001
R71031 vdd.n16330 vdd.n16310 0.001
R71032 vdd.n16577 vdd.n16576 0.001
R71033 vdd.n16754 vdd.n16753 0.001
R71034 vdd.n20664 vdd.n20662 0.001
R71035 vdd.n20648 vdd.n20646 0.001
R71036 vdd.n20615 vdd.n20613 0.001
R71037 vdd.n20599 vdd.n20597 0.001
R71038 vdd.n20467 vdd.n20466 0.001
R71039 vdd.n20411 vdd.n20409 0.001
R71040 vdd.n20369 vdd.n20367 0.001
R71041 vdd.n20303 vdd.n20301 0.001
R71042 vdd.n20287 vdd.n20285 0.001
R71043 vdd.n20267 vdd.n20255 0.001
R71044 vdd.n20251 vdd.n20239 0.001
R71045 vdd.n20175 vdd.n20173 0.001
R71046 vdd.n20133 vdd.n20131 0.001
R71047 vdd.n20067 vdd.n20065 0.001
R71048 vdd.n19487 vdd.n19485 0.001
R71049 vdd.n19499 vdd.n19487 0.001
R71050 vdd.n19514 vdd.n19502 0.001
R71051 vdd.n19546 vdd.n19544 0.001
R71052 vdd.n19562 vdd.n19560 0.001
R71053 vdd.n19564 vdd.n19562 0.001
R71054 vdd.n19580 vdd.n19578 0.001
R71055 vdd.n19596 vdd.n19594 0.001
R71056 vdd.n19655 vdd.n19653 0.001
R71057 vdd.n19671 vdd.n19669 0.001
R71058 vdd.n19687 vdd.n19685 0.001
R71059 vdd.n19699 vdd.n19687 0.001
R71060 vdd.n19715 vdd.n19703 0.001
R71061 vdd.n19731 vdd.n19730 0.001
R71062 vdd.n19748 vdd.n19746 0.001
R71063 vdd.n19764 vdd.n19762 0.001
R71064 vdd.n19766 vdd.n19764 0.001
R71065 vdd.n19782 vdd.n19780 0.001
R71066 vdd.n19798 vdd.n19796 0.001
R71067 vdd.n20995 vdd.n20993 0.001
R71068 vdd.n20979 vdd.n20977 0.001
R71069 vdd.n20963 vdd.n20961 0.001
R71070 vdd.n20961 vdd.n20959 0.001
R71071 vdd.n20945 vdd.n20943 0.001
R71072 vdd.n20928 vdd.n20927 0.001
R71073 vdd.n20912 vdd.n20900 0.001
R71074 vdd.n20896 vdd.n20884 0.001
R71075 vdd.n20884 vdd.n20882 0.001
R71076 vdd.n20868 vdd.n20866 0.001
R71077 vdd.n20863 vdd.n20861 0.001
R71078 vdd.n20804 vdd.n20802 0.001
R71079 vdd.n20788 vdd.n20786 0.001
R71080 vdd.n20772 vdd.n20770 0.001
R71081 vdd.n20770 vdd.n20769 0.001
R71082 vdd.n20755 vdd.n20753 0.001
R71083 vdd.n20723 vdd.n20711 0.001
R71084 vdd.n20708 vdd.n20696 0.001
R71085 vdd.n20696 vdd.n20694 0.001
R71086 vdd.n19390 vdd.n19388 0.001
R71087 vdd.n19406 vdd.n19404 0.001
R71088 vdd.n19439 vdd.n19437 0.001
R71089 vdd.n19455 vdd.n19453 0.001
R71090 vdd.n21798 vdd.n21771 0.001
R71091 vdd.n21960 vdd.n21900 0.001
R71092 vdd.n21747 vdd.n21746 0.001
R71093 vdd.n24734 vdd.n24732 0.001
R71094 vdd.n24762 vdd.n24760 0.001
R71095 vdd.n24830 vdd.n24822 0.001
R71096 vdd.n25248 vdd.n25240 0.001
R71097 vdd.n25180 vdd.n25178 0.001
R71098 vdd.n25152 vdd.n25150 0.001
R71099 vdd.n30558 vdd.n30557 0.001
R71100 vdd.n4019 vdd.n4016 0.001
R71101 vdd.n4019 vdd.n4018 0.001
R71102 vdd.n24837 vdd.n24836 0.001
R71103 vdd.n25363 vdd.n25362 0.001
R71104 vdd.n25263 vdd.n25262 0.001
R71105 vdd.n31206 vdd.n31205 0.001
R71106 vdd.n32390 vdd.n31446 0.001
R71107 vdd.n24863 vdd.n24862 0.001
R71108 vdd.n24836 vdd.n24835 0.001
R71109 vdd.n24835 vdd.n24834 0.001
R71110 vdd.n24879 vdd.n24878 0.001
R71111 vdd.n24878 vdd.n24877 0.001
R71112 vdd.n31221 vdd.n31220 0.001
R71113 vdd.n26292 vdd.n26291 0.001
R71114 vdd.n31214 vdd.n31213 0.001
R71115 vdd.n31383 vdd.n31382 0.001
R71116 vdd.n30971 vdd.n30970 0.001
R71117 vdd.n30763 vdd.n30762 0.001
R71118 vdd.n29206 vdd.n29185 0.001
R71119 vdd.n29294 vdd.n29288 0.001
R71120 vdd.n29433 vdd.n29432 0.001
R71121 vdd.n7186 vdd.n7185 0.001
R71122 vdd.n29552 vdd.n29534 0.001
R71123 vdd.n32679 vdd.n32678 0.001
R71124 vdd.n32703 vdd.n32645 0.001
R71125 vdd.n29995 vdd.n29961 0.001
R71126 vdd.n30087 vdd.n30081 0.001
R71127 vdd.n31429 vdd.n31428 0.001
R71128 vdd.n32563 vdd.n32538 0.001
R71129 vdd.n31441 vdd.n31433 0.001
R71130 vdd.n30831 vdd.n30816 0.001
R71131 vdd.n30740 vdd.n30736 0.001
R71132 vdd.n31226 vdd.n31225 0.001
R71133 vdd.n29136 vdd.n29119 0.001
R71134 vdd.n29098 vdd.n29097 0.001
R71135 vdd.n26524 vdd.n26476 0.001
R71136 vdd.n26391 vdd.n26390 0.001
R71137 vdd.n26321 vdd.n26320 0.001
R71138 vdd.n26182 vdd.n26181 0.001
R71139 vdd.n26665 vdd.n26658 0.001
R71140 vdd.n29101 vdd.n29044 0.001
R71141 vdd.n32106 vdd.n32090 0.001
R71142 vdd.n32513 vdd.n32511 0.001
R71143 vdd.n31225 vdd.n31216 0.001
R71144 vdd.n26724 vdd.n26723 0.001
R71145 vdd.n3886 vdd.n3885 0.001
R71146 vdd.n30577 vdd.n30576 0.001
R71147 vdd.n7173 vdd.n7155 0.001
R71148 vdd.n30860 vdd.n30833 0.001
R71149 vdd.n29336 vdd.n29315 0.001
R71150 vdd.n29513 vdd.n29502 0.001
R71151 vdd.n30125 vdd.n30108 0.001
R71152 vdd.n30776 vdd.n30771 0.001
R71153 vdd.n26521 vdd.n26520 0.001
R71154 vdd.n26711 vdd.n26710 0.001
R71155 vdd.n26467 vdd.n26466 0.001
R71156 vdd.n32737 vdd.n29566 0.001
R71157 vdd.n32738 vdd.n32737 0.001
R71158 vdd.n1826 vdd.n1825 0.001
R71159 vdd.n1837 vdd.n1249 0.001
R71160 vdd.n32002 vdd.n32001 0.001
R71161 vdd.n32329 vdd.n32328 0.001
R71162 vdd.n32346 vdd.n32345 0.001
R71163 vdd.n32737 vdd.n7219 0.001
R71164 vdd.n32737 vdd.n7177 0.001
R71165 vdd.n32812 vdd.n6373 0.001
R71166 vdd.n32812 vdd.n6364 0.001
R71167 vdd.n32807 vdd.n6439 0.001
R71168 vdd.n32802 vdd.n6496 0.001
R71169 vdd.n32796 vdd.n6554 0.001
R71170 vdd.n32790 vdd.n6606 0.001
R71171 vdd.n32785 vdd.n6667 0.001
R71172 vdd.n32780 vdd.n6719 0.001
R71173 vdd.n32775 vdd.n6779 0.001
R71174 vdd.n32769 vdd.n6836 0.001
R71175 vdd.n32760 vdd.n6918 0.001
R71176 vdd.n32757 vdd.n6949 0.001
R71177 vdd.n32754 vdd.n6975 0.001
R71178 vdd.n32751 vdd.n7006 0.001
R71179 vdd.n32748 vdd.n7031 0.001
R71180 vdd.n32745 vdd.n7061 0.001
R71181 vdd.n32742 vdd.n7085 0.001
R71182 vdd.n32737 vdd.n7188 0.001
R71183 vdd.n25335 vdd.n7226 0.001
R71184 vdd.n25332 vdd.n7256 0.001
R71185 vdd.n25329 vdd.n7284 0.001
R71186 vdd.n25326 vdd.n7313 0.001
R71187 vdd.n25323 vdd.n7337 0.001
R71188 vdd.n25320 vdd.n7369 0.001
R71189 vdd.n25318 vdd.n7395 0.001
R71190 vdd.n25315 vdd.n7425 0.001
R71191 vdd.n25312 vdd.n7452 0.001
R71192 vdd.n25309 vdd.n7476 0.001
R71193 vdd.n25306 vdd.n7507 0.001
R71194 vdd.n25303 vdd.n7537 0.001
R71195 vdd.n25301 vdd.n7563 0.001
R71196 vdd.n25298 vdd.n7595 0.001
R71197 vdd.n25296 vdd.n7621 0.001
R71198 vdd.n25293 vdd.n7652 0.001
R71199 vdd.n25291 vdd.n7678 0.001
R71200 vdd.n25288 vdd.n7709 0.001
R71201 vdd.n25286 vdd.n7735 0.001
R71202 vdd.n25284 vdd.n7764 0.001
R71203 vdd.n25281 vdd.n7793 0.001
R71204 vdd.n25278 vdd.n7824 0.001
R71205 vdd.n25275 vdd.n7850 0.001
R71206 vdd.n25272 vdd.n7881 0.001
R71207 vdd.n25269 vdd.n7907 0.001
R71208 vdd.n25266 vdd.n7935 0.001
R71209 vdd.n26136 vdd.n26135 0.001
R71210 vdd.n31379 vdd.n31378 0.001
R71211 vdd.n29655 vdd.n29654 0.001
R71212 vdd.n27732 vdd.n27730 0.001
R71213 vdd.n31233 vdd.n31232 0.001
R71214 vdd.n35619 vdd.n35618 0.001
R71215 vdd.n35029 vdd.n34444 0.001
R71216 vdd.n35615 vdd.n35030 0.001
R71217 vdd.n6362 vdd.n6361 0.001
R71218 vdd.n5191 vdd.n5190 0.001
R71219 vdd.n4607 vdd.n4606 0.001
R71220 vdd.n31202 vdd.n31201 0.001
R71221 vdd.n30140 vdd.n30138 0.001
R71222 vdd.n29354 vdd.n29352 0.001
R71223 vdd.n29192 vdd.n29191 0.001
R71224 vdd.n26564 vdd.n26562 0.001
R71225 vdd.n6404 vdd.n6403 0.001
R71226 vdd.n6372 vdd.n6370 0.001
R71227 vdd.n3803 vdd.n3802 0.001
R71228 vdd.n24368 vdd.n22043 0.001
R71229 vdd.n32811 vdd.n32809 0.001
R71230 vdd.n32808 vdd.n32807 0.001
R71231 vdd.n32806 vdd.n32804 0.001
R71232 vdd.n32803 vdd.n32802 0.001
R71233 vdd.n32801 vdd.n32799 0.001
R71234 vdd.n32798 vdd.n32796 0.001
R71235 vdd.n32795 vdd.n32793 0.001
R71236 vdd.n32792 vdd.n32790 0.001
R71237 vdd.n32789 vdd.n32788 0.001
R71238 vdd.n32787 vdd.n32785 0.001
R71239 vdd.n32784 vdd.n32782 0.001
R71240 vdd.n32781 vdd.n32780 0.001
R71241 vdd.n32779 vdd.n32778 0.001
R71242 vdd.n32777 vdd.n32775 0.001
R71243 vdd.n32774 vdd.n32772 0.001
R71244 vdd.n32771 vdd.n32769 0.001
R71245 vdd.n32768 vdd.n32766 0.001
R71246 vdd.n32765 vdd.n32763 0.001
R71247 vdd.n32762 vdd.n32760 0.001
R71248 vdd.n32759 vdd.n32757 0.001
R71249 vdd.n32756 vdd.n32754 0.001
R71250 vdd.n32753 vdd.n32751 0.001
R71251 vdd.n32750 vdd.n32748 0.001
R71252 vdd.n32747 vdd.n32745 0.001
R71253 vdd.n32744 vdd.n32742 0.001
R71254 vdd.n32741 vdd.n32739 0.001
R71255 vdd.n25336 vdd.n25335 0.001
R71256 vdd.n25334 vdd.n25332 0.001
R71257 vdd.n25331 vdd.n25329 0.001
R71258 vdd.n25328 vdd.n25326 0.001
R71259 vdd.n25325 vdd.n25323 0.001
R71260 vdd.n25322 vdd.n25320 0.001
R71261 vdd.n25319 vdd.n25318 0.001
R71262 vdd.n25317 vdd.n25315 0.001
R71263 vdd.n25314 vdd.n25312 0.001
R71264 vdd.n25311 vdd.n25309 0.001
R71265 vdd.n25308 vdd.n25306 0.001
R71266 vdd.n25305 vdd.n25303 0.001
R71267 vdd.n25302 vdd.n25301 0.001
R71268 vdd.n25300 vdd.n25298 0.001
R71269 vdd.n25297 vdd.n25296 0.001
R71270 vdd.n25295 vdd.n25293 0.001
R71271 vdd.n25292 vdd.n25291 0.001
R71272 vdd.n25290 vdd.n25288 0.001
R71273 vdd.n25287 vdd.n25286 0.001
R71274 vdd.n25285 vdd.n25284 0.001
R71275 vdd.n25283 vdd.n25281 0.001
R71276 vdd.n25280 vdd.n25278 0.001
R71277 vdd.n25277 vdd.n25275 0.001
R71278 vdd.n25274 vdd.n25272 0.001
R71279 vdd.n25271 vdd.n25269 0.001
R71280 vdd.n25268 vdd.n25266 0.001
R71281 vdd.n25265 vdd.n25264 0.001
R71282 vdd.n32737 vdd.n27661 0.001
R71283 vdd.n27661 vdd.n27660 0.001
R71284 vdd.n33862 vdd.n33861 0.001
R71285 vdd.n34442 vdd.n34441 0.001
R71286 vdd.n35614 vdd.n35613 0.001
R71287 vdd.n35028 vdd.n35027 0.001
R71288 vdd.n1175 vdd.n1174 0.001
R71289 vdd.n589 vdd.n588 0.001
R71290 vdd.n6360 vdd.n6359 0.001
R71291 vdd.n5774 vdd.n5773 0.001
R71292 vdd.n5188 vdd.n5187 0.001
R71293 vdd.n4604 vdd.n4603 0.001
R71294 vdd.n4020 vdd.n2676 0.001
R71295 vdd.n2676 vdd.n2563 0.001
R71296 vdd.n4605 vdd.n4604 0.001
R71297 vdd.n5189 vdd.n5188 0.001
R71298 vdd.n5775 vdd.n5774 0.001
R71299 vdd.n6359 vdd.n6358 0.001
R71300 vdd.n588 vdd.n587 0.001
R71301 vdd.n1174 vdd.n1173 0.001
R71302 vdd.n35027 vdd.n35026 0.001
R71303 vdd.n35613 vdd.n35612 0.001
R71304 vdd.n34443 vdd.n34442 0.001
R71305 vdd.n33863 vdd.n33862 0.001
R71306 vdd.n2547 vdd.n2546 0.001
R71307 vdd.n32812 vdd.n32811 0.001
R71308 vdd.n32809 vdd.n32808 0.001
R71309 vdd.n32807 vdd.n32806 0.001
R71310 vdd.n32804 vdd.n32803 0.001
R71311 vdd.n32802 vdd.n32801 0.001
R71312 vdd.n32799 vdd.n32798 0.001
R71313 vdd.n32796 vdd.n32795 0.001
R71314 vdd.n32793 vdd.n32792 0.001
R71315 vdd.n32790 vdd.n32789 0.001
R71316 vdd.n32788 vdd.n32787 0.001
R71317 vdd.n32785 vdd.n32784 0.001
R71318 vdd.n32782 vdd.n32781 0.001
R71319 vdd.n32780 vdd.n32779 0.001
R71320 vdd.n32778 vdd.n32777 0.001
R71321 vdd.n32775 vdd.n32774 0.001
R71322 vdd.n32772 vdd.n32771 0.001
R71323 vdd.n32769 vdd.n32768 0.001
R71324 vdd.n32766 vdd.n32765 0.001
R71325 vdd.n32763 vdd.n32762 0.001
R71326 vdd.n32760 vdd.n32759 0.001
R71327 vdd.n32757 vdd.n32756 0.001
R71328 vdd.n32754 vdd.n32753 0.001
R71329 vdd.n32751 vdd.n32750 0.001
R71330 vdd.n32748 vdd.n32747 0.001
R71331 vdd.n32745 vdd.n32744 0.001
R71332 vdd.n32742 vdd.n32741 0.001
R71333 vdd.n32737 vdd.n25336 0.001
R71334 vdd.n25335 vdd.n25334 0.001
R71335 vdd.n25332 vdd.n25331 0.001
R71336 vdd.n25329 vdd.n25328 0.001
R71337 vdd.n25326 vdd.n25325 0.001
R71338 vdd.n25323 vdd.n25322 0.001
R71339 vdd.n25320 vdd.n25319 0.001
R71340 vdd.n25318 vdd.n25317 0.001
R71341 vdd.n25315 vdd.n25314 0.001
R71342 vdd.n25312 vdd.n25311 0.001
R71343 vdd.n25309 vdd.n25308 0.001
R71344 vdd.n25306 vdd.n25305 0.001
R71345 vdd.n25303 vdd.n25302 0.001
R71346 vdd.n25301 vdd.n25300 0.001
R71347 vdd.n25298 vdd.n25297 0.001
R71348 vdd.n25296 vdd.n25295 0.001
R71349 vdd.n25293 vdd.n25292 0.001
R71350 vdd.n25291 vdd.n25290 0.001
R71351 vdd.n25288 vdd.n25287 0.001
R71352 vdd.n25286 vdd.n25285 0.001
R71353 vdd.n25284 vdd.n25283 0.001
R71354 vdd.n25281 vdd.n25280 0.001
R71355 vdd.n25278 vdd.n25277 0.001
R71356 vdd.n25275 vdd.n25274 0.001
R71357 vdd.n25272 vdd.n25271 0.001
R71358 vdd.n25269 vdd.n25268 0.001
R71359 vdd.n25266 vdd.n25265 0.001
R71360 vdd.n24864 vdd.n24863 0.001
R71361 vdd.n24880 vdd.n24879 0.001
R71362 out.n5394 out.n5392 19.587
R71363 out.n6453 out.n6451 19.587
R71364 out.n7255 out.n7253 19.587
R71365 out.n1366 out.n1365 15.024
R71366 out.n2142 out.n2141 15.024
R71367 out.n2210 out.n2209 15.024
R71368 out.n13030 out.n13029 14.919
R71369 out.n13145 out.n13144 14.919
R71370 out.n12606 out.n12605 14.919
R71371 out.n12726 out.n12725 14.919
R71372 out.n12165 out.n12164 14.919
R71373 out.n12280 out.n12279 14.919
R71374 out.n13439 out.n13438 14.919
R71375 out.n13560 out.n13559 14.919
R71376 out.n11339 out.n11338 14.919
R71377 out.n11449 out.n11448 14.919
R71378 out.n10912 out.n10911 14.919
R71379 out.n11022 out.n11021 14.919
R71380 out.n11745 out.n11744 14.919
R71381 out.n11860 out.n11859 14.919
R71382 out.n13894 out.n13893 14.919
R71383 out.n14015 out.n14014 14.919
R71384 out.n10478 out.n10477 14.919
R71385 out.n10593 out.n10592 14.919
R71386 out.n14399 out.n14398 14.919
R71387 out.n14454 out.n14453 14.919
R71388 out.n14243 out.n14242 14.919
R71389 out.n1041 out.n1040 14.919
R71390 out.n5128 out.n5127 14.919
R71391 out.n5308 out.n5307 14.919
R71392 out.n5885 out.n5884 14.919
R71393 out.n10070 out.n10069 13.423
R71394 out.n12892 out.n12890 13.423
R71395 out.n12874 out.n12872 13.423
R71396 out.n12857 out.n12855 13.423
R71397 out.n12455 out.n12453 13.423
R71398 out.n12440 out.n12439 13.423
R71399 out.n12419 out.n12417 13.423
R71400 out.n12025 out.n12023 13.423
R71401 out.n12007 out.n12005 13.423
R71402 out.n11992 out.n11990 13.423
R71403 out.n13299 out.n13297 13.423
R71404 out.n13284 out.n13283 13.423
R71405 out.n13266 out.n13264 13.423
R71406 out.n11193 out.n11191 13.423
R71407 out.n11172 out.n11170 13.423
R71408 out.n11152 out.n11150 13.423
R71409 out.n10767 out.n10765 13.423
R71410 out.n10749 out.n10747 13.423
R71411 out.n10729 out.n10727 13.423
R71412 out.n11607 out.n11605 13.423
R71413 out.n11587 out.n11585 13.423
R71414 out.n11572 out.n11570 13.423
R71415 out.n13754 out.n13752 13.423
R71416 out.n13737 out.n13736 13.423
R71417 out.n13719 out.n13717 13.423
R71418 out.n10340 out.n10338 13.423
R71419 out.n10320 out.n10318 13.423
R71420 out.n10305 out.n10303 13.423
R71421 out.n14365 out.n14363 13.423
R71422 out.n14273 out.n14271 13.423
R71423 out.n14190 out.n14188 13.423
R71424 out.n979 out.n977 13.423
R71425 out.n5054 out.n5052 13.423
R71426 out.n4961 out.n4959 13.423
R71427 out.n5399 out.n5397 13.423
R71428 out.n5370 out.n5368 13.423
R71429 out.n6458 out.n6456 13.423
R71430 out.n6177 out.n6175 13.423
R71431 out.n5904 out.n5902 13.423
R71432 out.n7260 out.n7258 13.423
R71433 out.n10250 out.n10249 13.176
R71434 out.n5836 out.n5835 13.176
R71435 out.n6408 out.n6407 13.176
R71436 out.n6970 out.n6969 13.176
R71437 out.n7791 out.n7790 13.176
R71438 out.n5194 out.n5193 12.92
R71439 out.n7027 out.n7026 12.92
R71440 out.n1584 out.n1583 12.808
R71441 out.n2803 out.n2801 12.313
R71442 out.n1927 out.n1925 12.313
R71443 out.n1707 out.n1705 12.313
R71444 out.n7590 out.n7588 12.313
R71445 out.n2448 out.n2446 11.955
R71446 out.n5458 out.n5457 11.693
R71447 out.n6623 out.n6622 11.693
R71448 out.n7316 out.n7315 11.693
R71449 out.n5698 out.n5696 11.67
R71450 out.n6275 out.n6273 11.67
R71451 out.n6832 out.n6830 11.67
R71452 out.n7679 out.n7677 11.67
R71453 out.n5952 out.n5950 11.636
R71454 out.n12892 out.n12891 11.609
R71455 out.n12874 out.n12873 11.609
R71456 out.n12871 out.n12870 11.609
R71457 out.n12859 out.n12858 11.609
R71458 out.n12857 out.n12856 11.609
R71459 out.n12455 out.n12454 11.609
R71460 out.n12440 out.n12438 11.609
R71461 out.n12437 out.n12436 11.609
R71462 out.n12421 out.n12420 11.609
R71463 out.n12419 out.n12418 11.609
R71464 out.n12025 out.n12024 11.609
R71465 out.n12007 out.n12006 11.609
R71466 out.n12004 out.n12003 11.609
R71467 out.n11992 out.n11991 11.609
R71468 out.n11989 out.n11988 11.609
R71469 out.n13299 out.n13298 11.609
R71470 out.n13284 out.n13282 11.609
R71471 out.n13281 out.n13280 11.609
R71472 out.n13266 out.n13265 11.609
R71473 out.n13263 out.n13262 11.609
R71474 out.n11193 out.n11192 11.609
R71475 out.n11172 out.n11171 11.609
R71476 out.n11169 out.n11168 11.609
R71477 out.n11152 out.n11151 11.609
R71478 out.n11149 out.n11148 11.609
R71479 out.n10767 out.n10766 11.609
R71480 out.n10749 out.n10748 11.609
R71481 out.n10746 out.n10745 11.609
R71482 out.n10729 out.n10728 11.609
R71483 out.n10726 out.n10725 11.609
R71484 out.n11607 out.n11606 11.609
R71485 out.n11589 out.n11588 11.609
R71486 out.n11587 out.n11586 11.609
R71487 out.n11574 out.n11573 11.609
R71488 out.n11572 out.n11571 11.609
R71489 out.n13754 out.n13753 11.609
R71490 out.n13739 out.n13738 11.609
R71491 out.n13737 out.n13735 11.609
R71492 out.n13721 out.n13720 11.609
R71493 out.n13719 out.n13718 11.609
R71494 out.n10340 out.n10339 11.609
R71495 out.n10322 out.n10321 11.609
R71496 out.n10320 out.n10319 11.609
R71497 out.n10307 out.n10306 11.609
R71498 out.n10305 out.n10304 11.609
R71499 out.n14365 out.n14364 11.609
R71500 out.n14367 out.n14366 11.609
R71501 out.n14273 out.n14272 11.609
R71502 out.n14275 out.n14274 11.609
R71503 out.n14190 out.n14189 11.609
R71504 out.n979 out.n978 11.609
R71505 out.n5056 out.n5055 11.609
R71506 out.n5054 out.n5053 11.609
R71507 out.n4961 out.n4960 11.609
R71508 out.n4958 out.n4957 11.609
R71509 out.n5641 out.n5640 11.609
R71510 out.n5399 out.n5398 11.609
R71511 out.n5370 out.n5369 11.609
R71512 out.n5367 out.n5366 11.609
R71513 out.n5192 out.n5191 11.609
R71514 out.n6458 out.n6457 11.609
R71515 out.n6213 out.n6212 11.609
R71516 out.n6174 out.n6173 11.609
R71517 out.n6177 out.n6176 11.609
R71518 out.n5904 out.n5903 11.609
R71519 out.n6775 out.n6774 11.609
R71520 out.n7260 out.n7259 11.609
R71521 out.n7025 out.n7024 11.609
R71522 out.n7486 out.n7485 11.609
R71523 out.n12951 out.n12947 11.482
R71524 out.n12086 out.n12082 11.482
R71525 out.n11263 out.n11259 11.482
R71526 out.n10833 out.n10829 11.482
R71527 out.n11666 out.n11662 11.482
R71528 out.n10399 out.n10395 11.482
R71529 out.n975 out.n971 11.482
R71530 out.n6048 out.n6044 11.482
R71531 out.n5952 out.n5951 11.378
R71532 out.n5458 out.n5456 11.31
R71533 out.n6623 out.n6621 11.31
R71534 out.n7316 out.n7314 11.31
R71535 out.n1280 out.n1278 11.294
R71536 out.n7094 out.n7092 11.294
R71537 out.n5705 out.n5703 11.112
R71538 out.n6282 out.n6280 11.112
R71539 out.n6839 out.n6837 11.112
R71540 out.n7686 out.n7684 11.112
R71541 out.n5682 out.n5678 11.106
R71542 out.n6259 out.n6255 11.106
R71543 out.n6816 out.n6812 11.106
R71544 out.n7663 out.n7659 11.106
R71545 out.n2800 out.n2799 11.058
R71546 out.n1924 out.n1923 11.058
R71547 out.n1704 out.n1703 11.058
R71548 out.n7587 out.n7586 11.058
R71549 out.n1395 out.n1393 11.031
R71550 out.n2114 out.n2112 11.031
R71551 out.n2239 out.n2237 11.031
R71552 out.n5460 out.n5459 10.879
R71553 out.n6625 out.n6624 10.879
R71554 out.n7318 out.n7317 10.879
R71555 out.n1273 out.n1271 10.736
R71556 out.n7101 out.n7099 10.736
R71557 out.n2445 out.n2444 10.735
R71558 out.n1185 out.n1184 10.729
R71559 out.n7078 out.n7077 10.729
R71560 out.n5428 out.n5424 10.353
R71561 out.n6614 out.n6610 10.353
R71562 out.n7289 out.n7285 10.353
R71563 out.n1395 out.n1394 9.654
R71564 out.n2114 out.n2113 9.654
R71565 out.n2239 out.n2238 9.654
R71566 out.t1 out.n9428 9.362
R71567 out.n1323 out.n1141 9.312
R71568 out.n1607 out.n1539 9.307
R71569 out.n2932 out.n2731 9.305
R71570 out.n1836 out.n1635 9.305
R71571 out.n2061 out.n1860 9.305
R71572 out.n2708 out.n2622 9.305
R71573 out.n2584 out.n2389 9.303
R71574 out.n9436 out.n9433 9.3
R71575 out.n9436 out.n9426 9.3
R71576 out.n9437 out.n9436 9.3
R71577 out.n9442 out.n9436 9.3
R71578 out.n9455 out.n9454 9.3
R71579 out.n10105 out.n10104 9.3
R71580 out.n10118 out.n10117 9.3
R71581 out.n10144 out.n10143 9.3
R71582 out.n10142 out.n10141 9.3
R71583 out.n10199 out.n10198 9.3
R71584 out.n10196 out.n10195 9.3
R71585 out.n10201 out.n10200 9.3
R71586 out.n10233 out.n10232 9.3
R71587 out.n10242 out.n10241 9.3
R71588 out.n10235 out.n10234 9.3
R71589 out.n10256 out.n10255 9.3
R71590 out.n10259 out.n10258 9.3
R71591 out.n12897 out.n12896 9.3
R71592 out.n12906 out.n12905 9.3
R71593 out.n12913 out.n12912 9.3
R71594 out.n12920 out.n12919 9.3
R71595 out.n12929 out.n12928 9.3
R71596 out.n12927 out.n12926 9.3
R71597 out.n12963 out.n12962 9.3
R71598 out.n12956 out.n12955 9.3
R71599 out.n13019 out.n13018 9.3
R71600 out.n13021 out.n13020 9.3
R71601 out.n13031 out.n13030 9.3
R71602 out.n13038 out.n13037 9.3
R71603 out.n13047 out.n13046 9.3
R71604 out.n13045 out.n13044 9.3
R71605 out.n13072 out.n13071 9.3
R71606 out.n13074 out.n13073 9.3
R71607 out.n13095 out.n13094 9.3
R71608 out.n13101 out.n13100 9.3
R71609 out.n13136 out.n13135 9.3
R71610 out.n13146 out.n13145 9.3
R71611 out.n13155 out.n13154 9.3
R71612 out.n13153 out.n13152 9.3
R71613 out.n13196 out.n13195 9.3
R71614 out.n13184 out.n13183 9.3
R71615 out.n13186 out.n13185 9.3
R71616 out.n13198 out.n13197 9.3
R71617 out.n13226 out.n13225 9.3
R71618 out.n13229 out.n13228 9.3
R71619 out.n12473 out.n12472 9.3
R71620 out.n12482 out.n12481 9.3
R71621 out.n12489 out.n12488 9.3
R71622 out.n12496 out.n12495 9.3
R71623 out.n12505 out.n12504 9.3
R71624 out.n12503 out.n12502 9.3
R71625 out.n12530 out.n12529 9.3
R71626 out.n12595 out.n12594 9.3
R71627 out.n12597 out.n12596 9.3
R71628 out.n12607 out.n12606 9.3
R71629 out.n12614 out.n12613 9.3
R71630 out.n12623 out.n12622 9.3
R71631 out.n12621 out.n12620 9.3
R71632 out.n12650 out.n12649 9.3
R71633 out.n12652 out.n12651 9.3
R71634 out.n12677 out.n12676 9.3
R71635 out.n12673 out.n12672 9.3
R71636 out.n12670 out.n12669 9.3
R71637 out.n12680 out.n12679 9.3
R71638 out.n12708 out.n12707 9.3
R71639 out.n12711 out.n12710 9.3
R71640 out.n12717 out.n12716 9.3
R71641 out.n12727 out.n12726 9.3
R71642 out.n12773 out.n12772 9.3
R71643 out.n12763 out.n12762 9.3
R71644 out.n12800 out.n12799 9.3
R71645 out.n12803 out.n12802 9.3
R71646 out.n12032 out.n12031 9.3
R71647 out.n12041 out.n12040 9.3
R71648 out.n12048 out.n12047 9.3
R71649 out.n12055 out.n12054 9.3
R71650 out.n12064 out.n12063 9.3
R71651 out.n12062 out.n12061 9.3
R71652 out.n12098 out.n12097 9.3
R71653 out.n12091 out.n12090 9.3
R71654 out.n12154 out.n12153 9.3
R71655 out.n12156 out.n12155 9.3
R71656 out.n12166 out.n12165 9.3
R71657 out.n12173 out.n12172 9.3
R71658 out.n12182 out.n12181 9.3
R71659 out.n12180 out.n12179 9.3
R71660 out.n12207 out.n12206 9.3
R71661 out.n12209 out.n12208 9.3
R71662 out.n12230 out.n12229 9.3
R71663 out.n12236 out.n12235 9.3
R71664 out.n12271 out.n12270 9.3
R71665 out.n12281 out.n12280 9.3
R71666 out.n12290 out.n12289 9.3
R71667 out.n12288 out.n12287 9.3
R71668 out.n12331 out.n12330 9.3
R71669 out.n12319 out.n12318 9.3
R71670 out.n12321 out.n12320 9.3
R71671 out.n12333 out.n12332 9.3
R71672 out.n12361 out.n12360 9.3
R71673 out.n12364 out.n12363 9.3
R71674 out.n13306 out.n13305 9.3
R71675 out.n13315 out.n13314 9.3
R71676 out.n13322 out.n13321 9.3
R71677 out.n13329 out.n13328 9.3
R71678 out.n13338 out.n13337 9.3
R71679 out.n13336 out.n13335 9.3
R71680 out.n13363 out.n13362 9.3
R71681 out.n13428 out.n13427 9.3
R71682 out.n13430 out.n13429 9.3
R71683 out.n13440 out.n13439 9.3
R71684 out.n13447 out.n13446 9.3
R71685 out.n13456 out.n13455 9.3
R71686 out.n13454 out.n13453 9.3
R71687 out.n13483 out.n13482 9.3
R71688 out.n13485 out.n13484 9.3
R71689 out.n13511 out.n13510 9.3
R71690 out.n13506 out.n13505 9.3
R71691 out.n13503 out.n13502 9.3
R71692 out.n13514 out.n13513 9.3
R71693 out.n13542 out.n13541 9.3
R71694 out.n13545 out.n13544 9.3
R71695 out.n13551 out.n13550 9.3
R71696 out.n13561 out.n13560 9.3
R71697 out.n13607 out.n13606 9.3
R71698 out.n13597 out.n13596 9.3
R71699 out.n13634 out.n13633 9.3
R71700 out.n13637 out.n13636 9.3
R71701 out.n11209 out.n11208 9.3
R71702 out.n11218 out.n11217 9.3
R71703 out.n11225 out.n11224 9.3
R71704 out.n11232 out.n11231 9.3
R71705 out.n11241 out.n11240 9.3
R71706 out.n11239 out.n11238 9.3
R71707 out.n11275 out.n11274 9.3
R71708 out.n11268 out.n11267 9.3
R71709 out.n11328 out.n11327 9.3
R71710 out.n11330 out.n11329 9.3
R71711 out.n11340 out.n11339 9.3
R71712 out.n11347 out.n11346 9.3
R71713 out.n11356 out.n11355 9.3
R71714 out.n11354 out.n11353 9.3
R71715 out.n11381 out.n11380 9.3
R71716 out.n11383 out.n11382 9.3
R71717 out.n11404 out.n11403 9.3
R71718 out.n11410 out.n11409 9.3
R71719 out.n11440 out.n11439 9.3
R71720 out.n11450 out.n11449 9.3
R71721 out.n11459 out.n11458 9.3
R71722 out.n11457 out.n11456 9.3
R71723 out.n11500 out.n11499 9.3
R71724 out.n11488 out.n11487 9.3
R71725 out.n11490 out.n11489 9.3
R71726 out.n11502 out.n11501 9.3
R71727 out.n11530 out.n11529 9.3
R71728 out.n11533 out.n11532 9.3
R71729 out.n10779 out.n10778 9.3
R71730 out.n10788 out.n10787 9.3
R71731 out.n10795 out.n10794 9.3
R71732 out.n10802 out.n10801 9.3
R71733 out.n10811 out.n10810 9.3
R71734 out.n10809 out.n10808 9.3
R71735 out.n10845 out.n10844 9.3
R71736 out.n10838 out.n10837 9.3
R71737 out.n10901 out.n10900 9.3
R71738 out.n10903 out.n10902 9.3
R71739 out.n10913 out.n10912 9.3
R71740 out.n10920 out.n10919 9.3
R71741 out.n10929 out.n10928 9.3
R71742 out.n10927 out.n10926 9.3
R71743 out.n10954 out.n10953 9.3
R71744 out.n10956 out.n10955 9.3
R71745 out.n10977 out.n10976 9.3
R71746 out.n10983 out.n10982 9.3
R71747 out.n11013 out.n11012 9.3
R71748 out.n11023 out.n11022 9.3
R71749 out.n11032 out.n11031 9.3
R71750 out.n11030 out.n11029 9.3
R71751 out.n11073 out.n11072 9.3
R71752 out.n11061 out.n11060 9.3
R71753 out.n11063 out.n11062 9.3
R71754 out.n11075 out.n11074 9.3
R71755 out.n11103 out.n11102 9.3
R71756 out.n11106 out.n11105 9.3
R71757 out.n11612 out.n11611 9.3
R71758 out.n11621 out.n11620 9.3
R71759 out.n11628 out.n11627 9.3
R71760 out.n11635 out.n11634 9.3
R71761 out.n11644 out.n11643 9.3
R71762 out.n11642 out.n11641 9.3
R71763 out.n11678 out.n11677 9.3
R71764 out.n11671 out.n11670 9.3
R71765 out.n11734 out.n11733 9.3
R71766 out.n11736 out.n11735 9.3
R71767 out.n11746 out.n11745 9.3
R71768 out.n11753 out.n11752 9.3
R71769 out.n11762 out.n11761 9.3
R71770 out.n11760 out.n11759 9.3
R71771 out.n11787 out.n11786 9.3
R71772 out.n11789 out.n11788 9.3
R71773 out.n11810 out.n11809 9.3
R71774 out.n11816 out.n11815 9.3
R71775 out.n11851 out.n11850 9.3
R71776 out.n11861 out.n11860 9.3
R71777 out.n11870 out.n11869 9.3
R71778 out.n11868 out.n11867 9.3
R71779 out.n11911 out.n11910 9.3
R71780 out.n11899 out.n11898 9.3
R71781 out.n11901 out.n11900 9.3
R71782 out.n11913 out.n11912 9.3
R71783 out.n11941 out.n11940 9.3
R71784 out.n11944 out.n11943 9.3
R71785 out.n13761 out.n13760 9.3
R71786 out.n13770 out.n13769 9.3
R71787 out.n13777 out.n13776 9.3
R71788 out.n13784 out.n13783 9.3
R71789 out.n13793 out.n13792 9.3
R71790 out.n13791 out.n13790 9.3
R71791 out.n13818 out.n13817 9.3
R71792 out.n13883 out.n13882 9.3
R71793 out.n13885 out.n13884 9.3
R71794 out.n13895 out.n13894 9.3
R71795 out.n13902 out.n13901 9.3
R71796 out.n13911 out.n13910 9.3
R71797 out.n13909 out.n13908 9.3
R71798 out.n13938 out.n13937 9.3
R71799 out.n13940 out.n13939 9.3
R71800 out.n13966 out.n13965 9.3
R71801 out.n13961 out.n13960 9.3
R71802 out.n13958 out.n13957 9.3
R71803 out.n13969 out.n13968 9.3
R71804 out.n13997 out.n13996 9.3
R71805 out.n14000 out.n13999 9.3
R71806 out.n14006 out.n14005 9.3
R71807 out.n14016 out.n14015 9.3
R71808 out.n14062 out.n14061 9.3
R71809 out.n14052 out.n14051 9.3
R71810 out.n14089 out.n14088 9.3
R71811 out.n14092 out.n14091 9.3
R71812 out.n10345 out.n10344 9.3
R71813 out.n10354 out.n10353 9.3
R71814 out.n10361 out.n10360 9.3
R71815 out.n10368 out.n10367 9.3
R71816 out.n10377 out.n10376 9.3
R71817 out.n10375 out.n10374 9.3
R71818 out.n10411 out.n10410 9.3
R71819 out.n10404 out.n10403 9.3
R71820 out.n10467 out.n10466 9.3
R71821 out.n10469 out.n10468 9.3
R71822 out.n10479 out.n10478 9.3
R71823 out.n10486 out.n10485 9.3
R71824 out.n10495 out.n10494 9.3
R71825 out.n10493 out.n10492 9.3
R71826 out.n10520 out.n10519 9.3
R71827 out.n10522 out.n10521 9.3
R71828 out.n10543 out.n10542 9.3
R71829 out.n10549 out.n10548 9.3
R71830 out.n10584 out.n10583 9.3
R71831 out.n10594 out.n10593 9.3
R71832 out.n10603 out.n10602 9.3
R71833 out.n10601 out.n10600 9.3
R71834 out.n10644 out.n10643 9.3
R71835 out.n10632 out.n10631 9.3
R71836 out.n10634 out.n10633 9.3
R71837 out.n10646 out.n10645 9.3
R71838 out.n10674 out.n10673 9.3
R71839 out.n10677 out.n10676 9.3
R71840 out.n14169 out.n14168 9.3
R71841 out.n14171 out.n14170 9.3
R71842 out.n14400 out.n14399 9.3
R71843 out.n14407 out.n14406 9.3
R71844 out.n14393 out.n14392 9.3
R71845 out.n14391 out.n14390 9.3
R71846 out.n14418 out.n14417 9.3
R71847 out.n14354 out.n14353 9.3
R71848 out.n14178 out.n14152 9.3
R71849 out.n14445 out.n14444 9.3
R71850 out.n14455 out.n14454 9.3
R71851 out.n14464 out.n14463 9.3
R71852 out.n14462 out.n14461 9.3
R71853 out.n14286 out.n14285 9.3
R71854 out.n14288 out.n14287 9.3
R71855 out.n14297 out.n14296 9.3
R71856 out.n14299 out.n14298 9.3
R71857 out.n14488 out.n14487 9.3
R71858 out.n14491 out.n14490 9.3
R71859 out.n14250 out.n14249 9.3
R71860 out.n14247 out.n14246 9.3
R71861 out.n14501 out.n14500 9.3
R71862 out.n14244 out.n14243 9.3
R71863 out.n14513 out.n14512 9.3
R71864 out.n14515 out.n14514 9.3
R71865 out.n14545 out.n14544 9.3
R71866 out.n14548 out.n14547 9.3
R71867 out.n14536 out.n14535 9.3
R71868 out.n14539 out.n14538 9.3
R71869 out.n1107 out.n1106 9.3
R71870 out.n946 out.n945 9.3
R71871 out.n1097 out.n1096 9.3
R71872 out.n1090 out.n1089 9.3
R71873 out.n949 out.n948 9.3
R71874 out.n952 out.n951 9.3
R71875 out.n955 out.n954 9.3
R71876 out.n1077 out.n1076 9.3
R71877 out.n1069 out.n1068 9.3
R71878 out.n1071 out.n1070 9.3
R71879 out.n1030 out.n1029 9.3
R71880 out.n1032 out.n1031 9.3
R71881 out.n1042 out.n1041 9.3
R71882 out.n1035 out.n1034 9.3
R71883 out.n5082 out.n5081 9.3
R71884 out.n5080 out.n5079 9.3
R71885 out.n5092 out.n5091 9.3
R71886 out.n5043 out.n5042 9.3
R71887 out.n5119 out.n5118 9.3
R71888 out.n5129 out.n5128 9.3
R71889 out.n5138 out.n5137 9.3
R71890 out.n5136 out.n5135 9.3
R71891 out.n4986 out.n4985 9.3
R71892 out.n4972 out.n4971 9.3
R71893 out.n4984 out.n4983 9.3
R71894 out.n4974 out.n4973 9.3
R71895 out.n5165 out.n5164 9.3
R71896 out.n5162 out.n5161 9.3
R71897 out.n2738 out.n2737 9.3
R71898 out.n2735 out.n2734 9.3
R71899 out.n5818 out.n5817 9.3
R71900 out.n5827 out.n5826 9.3
R71901 out.n5825 out.n5824 9.3
R71902 out.n5802 out.n5801 9.3
R71903 out.n5800 out.n5799 9.3
R71904 out.n5793 out.n5792 9.3
R71905 out.n5791 out.n5790 9.3
R71906 out.n5784 out.n5783 9.3
R71907 out.n5777 out.n5776 9.3
R71908 out.n5768 out.n5767 9.3
R71909 out.n5762 out.n5761 9.3
R71910 out.n5759 out.n5758 9.3
R71911 out.n5687 out.n5686 9.3
R71912 out.n5694 out.n5693 9.3
R71913 out.n5701 out.n5700 9.3
R71914 out.n5671 out.n5670 9.3
R71915 out.n5669 out.n5668 9.3
R71916 out.n5662 out.n5661 9.3
R71917 out.n5660 out.n5659 9.3
R71918 out.n2877 out.n2876 9.3
R71919 out.n2872 out.n2871 9.3
R71920 out.n2865 out.n2864 9.3
R71921 out.n2869 out.n2868 9.3
R71922 out.n2863 out.n2862 9.3
R71923 out.n2815 out.n2814 9.3
R71924 out.n2755 out.n2754 9.3
R71925 out.n2762 out.n2761 9.3
R71926 out.n2752 out.n2751 9.3
R71927 out.n2758 out.n2757 9.3
R71928 out.n2766 out.n2765 9.3
R71929 out.n2771 out.n2770 9.3
R71930 out.n2775 out.n2774 9.3
R71931 out.n2784 out.n2783 9.3
R71932 out.n2934 out.n2933 9.3
R71933 out.n1346 out.n1345 9.3
R71934 out.n1343 out.n1342 9.3
R71935 out.n1352 out.n1351 9.3
R71936 out.n1352 out.n1349 9.3
R71937 out.n5574 out.n5573 9.3
R71938 out.n5583 out.n5582 9.3
R71939 out.n5572 out.n5571 9.3
R71940 out.n5581 out.n5580 9.3
R71941 out.n5547 out.n5546 9.3
R71942 out.n5545 out.n5544 9.3
R71943 out.n5538 out.n5537 9.3
R71944 out.n5531 out.n5530 9.3
R71945 out.n5524 out.n5523 9.3
R71946 out.n5515 out.n5514 9.3
R71947 out.n5436 out.n5435 9.3
R71948 out.n5434 out.n5433 9.3
R71949 out.n5439 out.n5438 9.3
R71950 out.n1462 out.n1461 9.3
R71951 out.n1457 out.n1456 9.3
R71952 out.n1449 out.n1448 9.3
R71953 out.n1453 out.n1452 9.3
R71954 out.n1476 out.n1475 9.3
R71955 out.n1430 out.n1429 9.3
R71956 out.n1433 out.n1432 9.3
R71957 out.n1425 out.n1424 9.3
R71958 out.n1406 out.n1405 9.3
R71959 out.n1357 out.n1356 9.3
R71960 out.n1363 out.n1362 9.3
R71961 out.n1355 out.n1354 9.3
R71962 out.n1359 out.n1358 9.3
R71963 out.n1367 out.n1366 9.3
R71964 out.n1392 out.n1391 9.3
R71965 out.n5376 out.n5375 9.3
R71966 out.n5352 out.n5351 9.3
R71967 out.n5336 out.n5335 9.3
R71968 out.n5334 out.n5333 9.3
R71969 out.n5327 out.n5326 9.3
R71970 out.n5325 out.n5324 9.3
R71971 out.n5318 out.n5317 9.3
R71972 out.n5302 out.n5301 9.3
R71973 out.n5299 out.n5298 9.3
R71974 out.n5274 out.n5273 9.3
R71975 out.n5282 out.n5281 9.3
R71976 out.n5235 out.n5234 9.3
R71977 out.n5242 out.n5241 9.3
R71978 out.n5219 out.n5218 9.3
R71979 out.n5217 out.n5216 9.3
R71980 out.n5210 out.n5209 9.3
R71981 out.n5208 out.n5207 9.3
R71982 out.n5201 out.n5200 9.3
R71983 out.n1243 out.n1242 9.3
R71984 out.n1239 out.n1238 9.3
R71985 out.n1234 out.n1233 9.3
R71986 out.n1236 out.n1235 9.3
R71987 out.n1156 out.n1155 9.3
R71988 out.n1163 out.n1162 9.3
R71989 out.n1159 out.n1158 9.3
R71990 out.n1309 out.n1308 9.3
R71991 out.n1302 out.n1301 9.3
R71992 out.n1166 out.n1165 9.3
R71993 out.n1169 out.n1168 9.3
R71994 out.n1173 out.n1172 9.3
R71995 out.n1176 out.n1175 9.3
R71996 out.n1292 out.n1291 9.3
R71997 out.n1284 out.n1283 9.3
R71998 out.n1277 out.n1276 9.3
R71999 out.n1286 out.n1285 9.3
R72000 out.n1325 out.n1324 9.3
R72001 out.n2082 out.n2081 9.3
R72002 out.n2079 out.n2078 9.3
R72003 out.n2086 out.n2085 9.3
R72004 out.n6728 out.n6727 9.3
R72005 out.n6737 out.n6736 9.3
R72006 out.n6726 out.n6725 9.3
R72007 out.n6735 out.n6734 9.3
R72008 out.n6701 out.n6700 9.3
R72009 out.n6699 out.n6698 9.3
R72010 out.n6692 out.n6691 9.3
R72011 out.n6463 out.n6462 9.3
R72012 out.n6468 out.n6467 9.3
R72013 out.n6679 out.n6678 9.3
R72014 out.n6603 out.n6602 9.3
R72015 out.n6601 out.n6600 9.3
R72016 out.n6594 out.n6593 9.3
R72017 out.n6587 out.n6586 9.3
R72018 out.n6580 out.n6579 9.3
R72019 out.n6504 out.n6503 9.3
R72020 out.n6501 out.n6500 9.3
R72021 out.n6570 out.n6569 9.3
R72022 out.n6518 out.n6517 9.3
R72023 out.n6513 out.n6512 9.3
R72024 out.n6551 out.n6550 9.3
R72025 out.n6532 out.n6531 9.3
R72026 out.n2091 out.n2090 9.3
R72027 out.n2097 out.n2096 9.3
R72028 out.n2089 out.n2088 9.3
R72029 out.n2093 out.n2092 9.3
R72030 out.n2143 out.n2142 9.3
R72031 out.n2126 out.n2125 9.3
R72032 out.n1867 out.n1866 9.3
R72033 out.n1864 out.n1863 9.3
R72034 out.n6390 out.n6389 9.3
R72035 out.n6399 out.n6398 9.3
R72036 out.n6397 out.n6396 9.3
R72037 out.n6374 out.n6373 9.3
R72038 out.n6372 out.n6371 9.3
R72039 out.n6365 out.n6364 9.3
R72040 out.n6363 out.n6362 9.3
R72041 out.n6356 out.n6355 9.3
R72042 out.n6218 out.n6217 9.3
R72043 out.n6345 out.n6344 9.3
R72044 out.n6339 out.n6338 9.3
R72045 out.n6336 out.n6335 9.3
R72046 out.n6264 out.n6263 9.3
R72047 out.n6271 out.n6270 9.3
R72048 out.n6278 out.n6277 9.3
R72049 out.n6248 out.n6247 9.3
R72050 out.n6246 out.n6245 9.3
R72051 out.n6239 out.n6238 9.3
R72052 out.n6237 out.n6236 9.3
R72053 out.n2001 out.n2000 9.3
R72054 out.n1996 out.n1995 9.3
R72055 out.n1989 out.n1988 9.3
R72056 out.n1993 out.n1992 9.3
R72057 out.n1987 out.n1986 9.3
R72058 out.n1939 out.n1938 9.3
R72059 out.n1884 out.n1883 9.3
R72060 out.n1891 out.n1890 9.3
R72061 out.n1881 out.n1880 9.3
R72062 out.n1887 out.n1886 9.3
R72063 out.n2046 out.n2045 9.3
R72064 out.n1895 out.n1894 9.3
R72065 out.n1899 out.n1898 9.3
R72066 out.n1908 out.n1907 9.3
R72067 out.n2063 out.n2062 9.3
R72068 out.n1544 out.n1543 9.3
R72069 out.n1542 out.n1541 9.3
R72070 out.n6188 out.n6187 9.3
R72071 out.n6185 out.n6184 9.3
R72072 out.n6166 out.n6165 9.3
R72073 out.n6164 out.n6163 9.3
R72074 out.n6139 out.n6138 9.3
R72075 out.n6137 out.n6136 9.3
R72076 out.n6130 out.n6129 9.3
R72077 out.n5886 out.n5885 9.3
R72078 out.n6118 out.n6117 9.3
R72079 out.n6116 out.n6115 9.3
R72080 out.n6099 out.n6098 9.3
R72081 out.n6053 out.n6052 9.3
R72082 out.n6061 out.n6060 9.3
R72083 out.n6059 out.n6058 9.3
R72084 out.n6026 out.n6025 9.3
R72085 out.n6024 out.n6023 9.3
R72086 out.n6017 out.n6016 9.3
R72087 out.n5909 out.n5908 9.3
R72088 out.n5914 out.n5913 9.3
R72089 out.n6004 out.n6003 9.3
R72090 out.n1595 out.n1594 9.3
R72091 out.n1550 out.n1549 9.3
R72092 out.n1546 out.n1545 9.3
R72093 out.n1585 out.n1584 9.3
R72094 out.n1578 out.n1577 9.3
R72095 out.n1553 out.n1552 9.3
R72096 out.n1642 out.n1641 9.3
R72097 out.n1639 out.n1638 9.3
R72098 out.n6952 out.n6951 9.3
R72099 out.n6961 out.n6960 9.3
R72100 out.n6959 out.n6958 9.3
R72101 out.n6936 out.n6935 9.3
R72102 out.n6934 out.n6933 9.3
R72103 out.n6927 out.n6926 9.3
R72104 out.n6925 out.n6924 9.3
R72105 out.n6918 out.n6917 9.3
R72106 out.n6911 out.n6910 9.3
R72107 out.n6902 out.n6901 9.3
R72108 out.n6896 out.n6895 9.3
R72109 out.n6893 out.n6892 9.3
R72110 out.n6821 out.n6820 9.3
R72111 out.n6828 out.n6827 9.3
R72112 out.n6835 out.n6834 9.3
R72113 out.n6805 out.n6804 9.3
R72114 out.n6803 out.n6802 9.3
R72115 out.n6796 out.n6795 9.3
R72116 out.n6794 out.n6793 9.3
R72117 out.n1781 out.n1780 9.3
R72118 out.n1776 out.n1775 9.3
R72119 out.n1769 out.n1768 9.3
R72120 out.n1773 out.n1772 9.3
R72121 out.n1767 out.n1766 9.3
R72122 out.n1719 out.n1718 9.3
R72123 out.n1659 out.n1658 9.3
R72124 out.n1666 out.n1665 9.3
R72125 out.n1656 out.n1655 9.3
R72126 out.n1662 out.n1661 9.3
R72127 out.n1670 out.n1669 9.3
R72128 out.n1675 out.n1674 9.3
R72129 out.n1679 out.n1678 9.3
R72130 out.n1688 out.n1687 9.3
R72131 out.n1838 out.n1837 9.3
R72132 out.n2190 out.n2189 9.3
R72133 out.n2187 out.n2186 9.3
R72134 out.n2196 out.n2195 9.3
R72135 out.n2196 out.n2193 9.3
R72136 out.n7432 out.n7431 9.3
R72137 out.n7441 out.n7440 9.3
R72138 out.n7430 out.n7429 9.3
R72139 out.n7439 out.n7438 9.3
R72140 out.n7405 out.n7404 9.3
R72141 out.n7403 out.n7402 9.3
R72142 out.n7396 out.n7395 9.3
R72143 out.n7389 out.n7388 9.3
R72144 out.n7382 out.n7381 9.3
R72145 out.n7373 out.n7372 9.3
R72146 out.n7297 out.n7296 9.3
R72147 out.n7295 out.n7294 9.3
R72148 out.n2311 out.n2310 9.3
R72149 out.n2306 out.n2305 9.3
R72150 out.n2301 out.n2300 9.3
R72151 out.n2293 out.n2292 9.3
R72152 out.n2297 out.n2296 9.3
R72153 out.n2323 out.n2322 9.3
R72154 out.n2274 out.n2273 9.3
R72155 out.n2277 out.n2276 9.3
R72156 out.n2269 out.n2268 9.3
R72157 out.n2250 out.n2249 9.3
R72158 out.n2201 out.n2200 9.3
R72159 out.n2207 out.n2206 9.3
R72160 out.n2199 out.n2198 9.3
R72161 out.n2203 out.n2202 9.3
R72162 out.n2211 out.n2210 9.3
R72163 out.n2236 out.n2235 9.3
R72164 out.n2396 out.n2395 9.3
R72165 out.n2393 out.n2392 9.3
R72166 out.n2404 out.n2403 9.3
R72167 out.n2402 out.n2401 9.3
R72168 out.n2402 out.n2399 9.3
R72169 out.n7202 out.n7201 9.3
R72170 out.n7211 out.n7210 9.3
R72171 out.n7209 out.n7208 9.3
R72172 out.n7186 out.n7185 9.3
R72173 out.n7184 out.n7183 9.3
R72174 out.n7177 out.n7176 9.3
R72175 out.n7175 out.n7174 9.3
R72176 out.n7034 out.n7033 9.3
R72177 out.n7039 out.n7038 9.3
R72178 out.n7162 out.n7161 9.3
R72179 out.n7156 out.n7155 9.3
R72180 out.n7153 out.n7152 9.3
R72181 out.n7083 out.n7082 9.3
R72182 out.n7090 out.n7089 9.3
R72183 out.n7097 out.n7096 9.3
R72184 out.n7069 out.n7068 9.3
R72185 out.n7067 out.n7066 9.3
R72186 out.n7060 out.n7059 9.3
R72187 out.n7058 out.n7057 9.3
R72188 out.n2511 out.n2510 9.3
R72189 out.n2518 out.n2517 9.3
R72190 out.n2504 out.n2503 9.3
R72191 out.n2508 out.n2507 9.3
R72192 out.n2502 out.n2501 9.3
R72193 out.n2485 out.n2484 9.3
R72194 out.n2479 out.n2478 9.3
R72195 out.n2488 out.n2487 9.3
R72196 out.n2482 out.n2481 9.3
R72197 out.n2462 out.n2461 9.3
R72198 out.n2412 out.n2411 9.3
R72199 out.n2419 out.n2418 9.3
R72200 out.n2409 out.n2408 9.3
R72201 out.n2415 out.n2414 9.3
R72202 out.n2567 out.n2566 9.3
R72203 out.n2560 out.n2559 9.3
R72204 out.n2422 out.n2421 9.3
R72205 out.n2430 out.n2429 9.3
R72206 out.n2586 out.n2585 9.3
R72207 out.n2628 out.n2627 9.3
R72208 out.n2625 out.n2624 9.3
R72209 out.n7802 out.n7801 9.3
R72210 out.n7773 out.n7772 9.3
R72211 out.n7782 out.n7781 9.3
R72212 out.n7780 out.n7779 9.3
R72213 out.n7757 out.n7756 9.3
R72214 out.n7755 out.n7754 9.3
R72215 out.n7748 out.n7747 9.3
R72216 out.n7746 out.n7745 9.3
R72217 out.n7739 out.n7738 9.3
R72218 out.n7491 out.n7490 9.3
R72219 out.n7728 out.n7727 9.3
R72220 out.n7722 out.n7721 9.3
R72221 out.n7719 out.n7718 9.3
R72222 out.n7668 out.n7667 9.3
R72223 out.n7675 out.n7674 9.3
R72224 out.n7682 out.n7681 9.3
R72225 out.n7652 out.n7651 9.3
R72226 out.n7650 out.n7649 9.3
R72227 out.n7643 out.n7642 9.3
R72228 out.n7641 out.n7640 9.3
R72229 out.n7530 out.n7529 9.3
R72230 out.n7535 out.n7534 9.3
R72231 out.n7542 out.n7541 9.3
R72232 out.n7539 out.n7538 9.3
R72233 out.n7626 out.n7625 9.3
R72234 out.n7584 out.n7583 9.3
R72235 out.n2633 out.n2632 9.3
R72236 out.n2637 out.n2636 9.3
R72237 out.n2630 out.n2629 9.3
R72238 out.n2681 out.n2680 9.3
R72239 out.n2674 out.n2673 9.3
R72240 out.n2639 out.n2638 9.3
R72241 out.n2647 out.n2646 9.3
R72242 out.n1397 out.n1396 9.199
R72243 out.n2116 out.n2115 9.199
R72244 out.n2241 out.n2240 9.199
R72245 out.n6750 out.n6749 9.143
R72246 out.n5872 out.n5871 9.132
R72247 out.n12851 out.n12830 9.114
R72248 out.n12390 out.n12371 9.114
R72249 out.n11552 out.n11542 9.114
R72250 out.n11129 out.n11115 9.114
R72251 out.n11972 out.n11951 9.114
R72252 out.n10705 out.n10684 9.114
R72253 out.n1124 out.n1122 9.114
R72254 out.n1330 out.n1329 9.091
R72255 out.n14178 out.n14151 8.908
R72256 out.n14178 out.n14157 8.897
R72257 out.n1124 out.n1120 8.897
R72258 out.n14178 out.n14155 8.885
R72259 out.n1124 out.n1118 8.885
R72260 out.n12887 out.n12885 8.868
R72261 out.n12867 out.n12865 8.868
R72262 out.n13210 out.n13209 8.868
R72263 out.n12450 out.n12448 8.868
R72264 out.n12433 out.n12431 8.868
R72265 out.n12787 out.n12786 8.868
R72266 out.n12020 out.n12018 8.868
R72267 out.n12000 out.n11998 8.868
R72268 out.n12345 out.n12344 8.868
R72269 out.n13294 out.n13292 8.868
R72270 out.n13277 out.n13275 8.868
R72271 out.n13621 out.n13620 8.868
R72272 out.n11188 out.n11186 8.868
R72273 out.n11165 out.n11163 8.868
R72274 out.n11514 out.n11513 8.868
R72275 out.n10762 out.n10760 8.868
R72276 out.n10742 out.n10740 8.868
R72277 out.n11087 out.n11086 8.868
R72278 out.n11602 out.n11600 8.868
R72279 out.n11582 out.n11580 8.868
R72280 out.n11925 out.n11924 8.868
R72281 out.n13749 out.n13747 8.868
R72282 out.n13732 out.n13730 8.868
R72283 out.n14076 out.n14075 8.868
R72284 out.n10335 out.n10333 8.868
R72285 out.n10315 out.n10313 8.868
R72286 out.n10658 out.n10657 8.868
R72287 out.n14359 out.n14357 8.868
R72288 out.n14280 out.n14279 8.868
R72289 out.n14195 out.n14194 8.868
R72290 out.n983 out.n981 8.868
R72291 out.n5048 out.n5046 8.868
R72292 out.n4966 out.n4965 8.868
R72293 out.n5637 out.n5635 8.868
R72294 out.n5712 out.n5710 8.868
R72295 out.n5468 out.n5466 8.868
R72296 out.n5188 out.n5186 8.868
R72297 out.n1190 out.n1188 8.868
R72298 out.n6632 out.n6630 8.868
R72299 out.n6209 out.n6207 8.868
R72300 out.n6289 out.n6287 8.868
R72301 out.n6071 out.n6069 8.868
R72302 out.n5961 out.n5959 8.868
R72303 out.n6771 out.n6769 8.868
R72304 out.n6846 out.n6844 8.868
R72305 out.n7326 out.n7324 8.868
R72306 out.n7021 out.n7019 8.868
R72307 out.n7108 out.n7106 8.868
R72308 out.n7482 out.n7480 8.868
R72309 out.n7692 out.n7690 8.868
R72310 out.n12820 out.n12812 8.865
R72311 out.n13667 out.n13648 8.865
R72312 out.n13700 out.n13681 8.865
R72313 out.n1330 out.n1328 8.843
R72314 out.n12851 out.n12832 8.833
R72315 out.n12820 out.n12810 8.833
R72316 out.n12390 out.n12373 8.833
R72317 out.n13667 out.n13646 8.833
R72318 out.n11552 out.n11544 8.833
R72319 out.n11129 out.n11117 8.833
R72320 out.n11972 out.n11953 8.833
R72321 out.n13700 out.n13679 8.833
R72322 out.n10705 out.n10686 8.833
R72323 out.n1124 out.n1123 8.833
R72324 out.n1330 out.n1326 8.833
R72325 out.n5872 out.n5869 8.833
R72326 out.n7807 out.n7806 8.833
R72327 out.n2937 out.n2936 8.832
R72328 out.n2066 out.n2065 8.832
R72329 out.n1841 out.n1840 8.832
R72330 out.n2589 out.n2588 8.832
R72331 out.n2448 out.n2447 8.812
R72332 out.n2811 out.n2809 8.491
R72333 out.n1935 out.n1933 8.491
R72334 out.n1715 out.n1713 8.491
R72335 out.n7580 out.n7578 8.491
R72336 out.n2803 out.n2802 8.419
R72337 out.n1927 out.n1926 8.419
R72338 out.n1707 out.n1706 8.419
R72339 out.n7590 out.n7589 8.419
R72340 out.n5426 out.n5425 8.128
R72341 out.n1180 out.n1179 8.128
R72342 out.n6612 out.n6611 8.128
R72343 out.n7287 out.n7286 8.128
R72344 out.n7075 out.n7074 8.128
R72345 out.n2458 out.n2456 8.115
R72346 out.n5954 out.n5953 8.02
R72347 out.n1402 out.n1400 7.738
R72348 out.n6537 out.n6535 7.738
R72349 out.n2246 out.n2244 7.738
R72350 out.n10014 out.n10013 7.623
R72351 out.n5680 out.n5679 7.375
R72352 out.n6257 out.n6256 7.375
R72353 out.n6814 out.n6813 7.375
R72354 out.n7661 out.n7660 7.375
R72355 out.n10099 out.n10098 7.041
R72356 out.n12949 out.n12948 6.622
R72357 out.n12084 out.n12083 6.622
R72358 out.n11261 out.n11260 6.622
R72359 out.n10831 out.n10830 6.622
R72360 out.n11664 out.n11663 6.622
R72361 out.n10397 out.n10396 6.622
R72362 out.n973 out.n972 6.622
R72363 out.n6046 out.n6045 6.622
R72364 out.n12937 out.n12936 6.259
R72365 out.n12511 out.n12510 6.259
R72366 out.n12072 out.n12071 6.259
R72367 out.n13344 out.n13343 6.259
R72368 out.n11249 out.n11248 6.259
R72369 out.n10819 out.n10818 6.259
R72370 out.n11652 out.n11651 6.259
R72371 out.n13799 out.n13798 6.259
R72372 out.n10385 out.n10384 6.259
R72373 out.n967 out.n966 6.259
R72374 out.n5668 out.n5667 6.259
R72375 out.n5553 out.n5552 6.259
R72376 out.n5433 out.n5432 6.259
R72377 out.n1175 out.n1174 6.259
R72378 out.n6707 out.n6706 6.259
R72379 out.n6600 out.n6599 6.259
R72380 out.n6245 out.n6244 6.259
R72381 out.n6034 out.n6033 6.259
R72382 out.n6802 out.n6801 6.259
R72383 out.n7411 out.n7410 6.259
R72384 out.n7294 out.n7293 6.259
R72385 out.n7066 out.n7065 6.259
R72386 out.n7649 out.n7648 6.259
R72387 out.n12881 out.n12879 6.246
R72388 out.n12444 out.n12442 6.246
R72389 out.n12014 out.n12012 6.246
R72390 out.n13288 out.n13286 6.246
R72391 out.n11182 out.n11180 6.246
R72392 out.n10756 out.n10754 6.246
R72393 out.n11596 out.n11594 6.246
R72394 out.n13743 out.n13741 6.246
R72395 out.n10329 out.n10327 6.246
R72396 out.n14202 out.n14201 6.246
R72397 out.n990 out.n988 6.246
R72398 out.n5652 out.n5650 6.246
R72399 out.n2820 out.n2818 6.246
R72400 out.n5417 out.n5415 6.246
R72401 out.n1411 out.n1409 6.246
R72402 out.n1197 out.n1195 6.246
R72403 out.n6486 out.n6484 6.246
R72404 out.n6528 out.n6526 6.246
R72405 out.n6229 out.n6227 6.246
R72406 out.n1944 out.n1942 6.246
R72407 out.n5898 out.n5896 6.246
R72408 out.n5969 out.n5967 6.246
R72409 out.n6786 out.n6784 6.246
R72410 out.n1724 out.n1722 6.246
R72411 out.n7278 out.n7276 6.246
R72412 out.n2255 out.n2253 6.246
R72413 out.n7050 out.n7048 6.246
R72414 out.n2467 out.n2465 6.246
R72415 out.n7522 out.n7520 6.246
R72416 out.n7600 out.n7598 6.246
R72417 out.n10073 out.n10072 6.143
R72418 out.n10055 out.n10054 6.143
R72419 out.n12926 out.n12925 6.088
R72420 out.n13053 out.n13052 6.088
R72421 out.n12502 out.n12501 6.088
R72422 out.n12061 out.n12060 6.088
R72423 out.n12188 out.n12187 6.088
R72424 out.n13335 out.n13334 6.088
R72425 out.n11238 out.n11237 6.088
R72426 out.n11362 out.n11361 6.088
R72427 out.n10808 out.n10807 6.088
R72428 out.n10935 out.n10934 6.088
R72429 out.n11641 out.n11640 6.088
R72430 out.n11768 out.n11767 6.088
R72431 out.n13790 out.n13789 6.088
R72432 out.n10374 out.n10373 6.088
R72433 out.n10501 out.n10500 6.088
R72434 out.n14383 out.n14382 6.088
R72435 out.n954 out.n953 6.088
R72436 out.n5072 out.n5071 6.088
R72437 out.n5799 out.n5798 6.088
R72438 out.n5659 out.n5658 6.088
R72439 out.n2770 out.n2769 6.088
R72440 out.n5544 out.n5543 6.088
R72441 out.n5438 out.n5437 6.088
R72442 out.n1424 out.n1423 6.088
R72443 out.n5216 out.n5215 6.088
R72444 out.n1168 out.n1167 6.088
R72445 out.n6698 out.n6697 6.088
R72446 out.n6593 out.n6592 6.088
R72447 out.n6550 out.n6549 6.088
R72448 out.n6371 out.n6370 6.088
R72449 out.n6236 out.n6235 6.088
R72450 out.n1894 out.n1893 6.088
R72451 out.n6145 out.n6144 6.088
R72452 out.n6023 out.n6022 6.088
R72453 out.n1577 out.n1576 6.088
R72454 out.n6933 out.n6932 6.088
R72455 out.n6793 out.n6792 6.088
R72456 out.n1674 out.n1673 6.088
R72457 out.n7402 out.n7401 6.088
R72458 out.n2310 out.n2309 6.088
R72459 out.n2268 out.n2267 6.088
R72460 out.n7183 out.n7182 6.088
R72461 out.n7057 out.n7056 6.088
R72462 out.n2559 out.n2558 6.088
R72463 out.n7754 out.n7753 6.088
R72464 out.n7640 out.n7639 6.088
R72465 out.n2673 out.n2672 6.088
R72466 out.n12861 out.n12860 6.023
R72467 out.n12766 out.n12765 6.023
R72468 out.n11994 out.n11993 6.023
R72469 out.n13600 out.n13599 6.023
R72470 out.n11159 out.n11158 6.023
R72471 out.n10736 out.n10735 6.023
R72472 out.n11576 out.n11575 6.023
R72473 out.n14055 out.n14054 6.023
R72474 out.n10309 out.n10308 6.023
R72475 out.n5032 out.n5031 6.023
R72476 out.n12522 out.n12521 5.869
R72477 out.n13355 out.n13354 5.869
R72478 out.n13810 out.n13809 5.869
R72479 out.n14182 out.n14181 5.869
R72480 out.n5564 out.n5563 5.869
R72481 out.n6718 out.n6717 5.869
R72482 out.n7422 out.n7421 5.869
R72483 out.n5234 out.n5233 5.862
R72484 out.n7201 out.n7200 5.862
R72485 out.n1387 out.n1386 5.856
R72486 out.n2109 out.n2108 5.856
R72487 out.n2231 out.n2230 5.856
R72488 out.n5817 out.n5816 5.855
R72489 out.n6389 out.n6388 5.855
R72490 out.n6951 out.n6950 5.855
R72491 out.n7772 out.n7771 5.855
R72492 out.n10077 out.n10076 5.643
R72493 out.n5180 out.n5179 5.643
R72494 out.n5227 out.n5226 5.506
R72495 out.n7194 out.n7193 5.506
R72496 out.n2440 out.n2439 5.479
R72497 out.n12993 out.n12992 5.461
R72498 out.n12128 out.n12127 5.461
R72499 out.n11305 out.n11304 5.461
R72500 out.n10875 out.n10874 5.461
R72501 out.n11708 out.n11707 5.461
R72502 out.n10441 out.n10440 5.461
R72503 out.n1005 out.n1004 5.461
R72504 out.n5889 out.n5888 5.461
R72505 out.n10177 out.n10176 5.443
R72506 out.n12631 out.n12630 5.335
R72507 out.n13464 out.n13463 5.335
R72508 out.n13919 out.n13918 5.335
R72509 out.n14254 out.n14253 5.335
R72510 out.n10150 out.n10149 5.327
R72511 out.n5344 out.n5343 5.327
R72512 out.n10063 out.n10062 5.32
R72513 out.n13174 out.n13173 5.313
R72514 out.n12686 out.n12685 5.313
R72515 out.n12309 out.n12308 5.313
R72516 out.n13520 out.n13519 5.313
R72517 out.n11478 out.n11477 5.313
R72518 out.n11051 out.n11050 5.313
R72519 out.n11889 out.n11888 5.313
R72520 out.n13975 out.n13974 5.313
R72521 out.n10622 out.n10621 5.313
R72522 out.n14309 out.n14308 5.313
R72523 out.n4996 out.n4995 5.313
R72524 out.n13107 out.n13106 5.305
R72525 out.n12753 out.n12752 5.305
R72526 out.n12242 out.n12241 5.305
R72527 out.n13587 out.n13586 5.305
R72528 out.n11154 out.n11153 5.305
R72529 out.n10731 out.n10730 5.305
R72530 out.n11822 out.n11821 5.305
R72531 out.n14042 out.n14041 5.305
R72532 out.n10555 out.n10554 5.305
R72533 out.n14332 out.n14331 5.305
R72534 out.n5019 out.n5018 5.305
R72535 out.n5278 out.n5277 5.27
R72536 out.n2795 out.n2794 5.103
R72537 out.n1919 out.n1918 5.103
R72538 out.n1699 out.n1698 5.103
R72539 out.n2657 out.n2656 5.103
R72540 out.n5375 out.n5374 5.081
R72541 out.n13195 out.n13194 5.081
R72542 out.n12672 out.n12671 5.081
R72543 out.n12330 out.n12329 5.081
R72544 out.n13505 out.n13504 5.081
R72545 out.n11499 out.n11498 5.081
R72546 out.n11072 out.n11071 5.081
R72547 out.n11910 out.n11909 5.081
R72548 out.n13960 out.n13959 5.081
R72549 out.n10643 out.n10642 5.081
R72550 out.n14285 out.n14284 5.081
R72551 out.n4971 out.n4970 5.081
R72552 out.n10059 out.n10057 4.888
R72553 out.n10061 out.n10060 4.764
R72554 out.n5810 out.n5809 4.753
R72555 out.n6382 out.n6381 4.753
R72556 out.n6944 out.n6943 4.753
R72557 out.n7765 out.n7764 4.753
R72558 out.n13064 out.n13063 4.746
R72559 out.n12199 out.n12198 4.746
R72560 out.n11373 out.n11372 4.746
R72561 out.n10946 out.n10945 4.746
R72562 out.n11779 out.n11778 4.746
R72563 out.n10512 out.n10511 4.746
R72564 out.n14376 out.n14375 4.746
R72565 out.n5065 out.n5064 4.746
R72566 out.n6156 out.n6155 4.746
R72567 out.n1380 out.n1379 4.74
R72568 out.n2102 out.n2101 4.74
R72569 out.n2224 out.n2223 4.74
R72570 out.n12642 out.n12641 4.738
R72571 out.n13475 out.n13474 4.738
R72572 out.n13930 out.n13929 4.738
R72573 out.n14263 out.n14262 4.738
R72574 out.n5351 out.n5350 4.731
R72575 out.n5940 out.n5939 4.727
R72576 out.n10269 out.n10266 4.704
R72577 out.n13094 out.n13093 4.704
R72578 out.n12772 out.n12771 4.704
R72579 out.n12229 out.n12228 4.704
R72580 out.n13606 out.n13605 4.704
R72581 out.n11403 out.n11402 4.704
R72582 out.n10976 out.n10975 4.704
R72583 out.n11809 out.n11808 4.704
R72584 out.n14061 out.n14060 4.704
R72585 out.n10542 out.n10541 4.704
R72586 out.n14353 out.n14352 4.704
R72587 out.n5042 out.n5041 4.704
R72588 out.n6187 out.n6186 4.704
R72589 out.n10131 out.n10091 4.65
R72590 out.n10191 out.n10190 4.65
R72591 out.n10254 out.n10253 4.65
R72592 out.n13054 out.n13053 4.65
R72593 out.n13130 out.n13129 4.65
R72594 out.n13220 out.n13219 4.65
R72595 out.n12512 out.n12511 4.65
R72596 out.n12659 out.n12658 4.65
R72597 out.n12734 out.n12733 4.65
R72598 out.n12189 out.n12188 4.65
R72599 out.n12265 out.n12264 4.65
R72600 out.n12355 out.n12354 4.65
R72601 out.n13345 out.n13344 4.65
R72602 out.n13492 out.n13491 4.65
R72603 out.n13568 out.n13567 4.65
R72604 out.n11363 out.n11362 4.65
R72605 out.n11434 out.n11433 4.65
R72606 out.n11524 out.n11523 4.65
R72607 out.n10936 out.n10935 4.65
R72608 out.n11007 out.n11006 4.65
R72609 out.n11097 out.n11096 4.65
R72610 out.n11769 out.n11768 4.65
R72611 out.n11845 out.n11844 4.65
R72612 out.n11935 out.n11934 4.65
R72613 out.n13800 out.n13799 4.65
R72614 out.n13947 out.n13946 4.65
R72615 out.n14023 out.n14022 4.65
R72616 out.n10502 out.n10501 4.65
R72617 out.n10578 out.n10577 4.65
R72618 out.n10668 out.n10667 4.65
R72619 out.n14384 out.n14383 4.65
R72620 out.n14439 out.n14438 4.65
R72621 out.n14482 out.n14481 4.65
R72622 out.n14557 out.n14556 4.65
R72623 out.n5073 out.n5072 4.65
R72624 out.n5113 out.n5112 4.65
R72625 out.n5156 out.n5155 4.65
R72626 out.n5834 out.n5833 4.65
R72627 out.n2793 out.n2792 4.65
R72628 out.n5554 out.n5553 4.65
R72629 out.n5381 out.n5380 4.65
R72630 out.n5309 out.n5308 4.65
R72631 out.n1181 out.n1180 4.65
R72632 out.n6708 out.n6707 4.65
R72633 out.n6406 out.n6405 4.65
R72634 out.n1917 out.n1916 4.65
R72635 out.n6146 out.n6145 4.65
R72636 out.n6968 out.n6967 4.65
R72637 out.n1697 out.n1696 4.65
R72638 out.n7412 out.n7411 4.65
R72639 out.n7076 out.n7075 4.65
R72640 out.n7789 out.n7788 4.65
R72641 out.n2655 out.n2654 4.65
R72642 out.n12919 out.n12918 4.596
R72643 out.n13044 out.n13043 4.596
R72644 out.n12495 out.n12494 4.596
R72645 out.n12620 out.n12619 4.596
R72646 out.n12054 out.n12053 4.596
R72647 out.n12179 out.n12178 4.596
R72648 out.n13328 out.n13327 4.596
R72649 out.n13453 out.n13452 4.596
R72650 out.n11231 out.n11230 4.596
R72651 out.n11353 out.n11352 4.596
R72652 out.n10801 out.n10800 4.596
R72653 out.n10926 out.n10925 4.596
R72654 out.n11634 out.n11633 4.596
R72655 out.n11759 out.n11758 4.596
R72656 out.n13783 out.n13782 4.596
R72657 out.n13908 out.n13907 4.596
R72658 out.n10367 out.n10366 4.596
R72659 out.n10492 out.n10491 4.596
R72660 out.n14390 out.n14389 4.596
R72661 out.n14249 out.n14248 4.596
R72662 out.n948 out.n947 4.596
R72663 out.n5079 out.n5078 4.596
R72664 out.n5790 out.n5789 4.596
R72665 out.n2876 out.n2875 4.596
R72666 out.n2765 out.n2764 4.596
R72667 out.n5537 out.n5536 4.596
R72668 out.n1461 out.n1460 4.596
R72669 out.n5333 out.n5332 4.596
R72670 out.n5207 out.n5206 4.596
R72671 out.n1301 out.n1300 4.596
R72672 out.n6691 out.n6690 4.596
R72673 out.n6586 out.n6585 4.596
R72674 out.n6362 out.n6361 4.596
R72675 out.n2000 out.n1999 4.596
R72676 out.n2045 out.n2044 4.596
R72677 out.n6136 out.n6135 4.596
R72678 out.n6016 out.n6015 4.596
R72679 out.n6924 out.n6923 4.596
R72680 out.n1780 out.n1779 4.596
R72681 out.n1669 out.n1668 4.596
R72682 out.n7395 out.n7394 4.596
R72683 out.n2305 out.n2304 4.596
R72684 out.n7174 out.n7173 4.596
R72685 out.n2510 out.n2509 4.596
R72686 out.n2566 out.n2565 4.596
R72687 out.n7745 out.n7744 4.596
R72688 out.n7529 out.n7528 4.596
R72689 out.n2680 out.n2679 4.596
R72690 out.n13163 out.n13162 4.589
R72691 out.n12697 out.n12696 4.589
R72692 out.n12298 out.n12297 4.589
R72693 out.n13531 out.n13530 4.589
R72694 out.n11467 out.n11466 4.589
R72695 out.n11040 out.n11039 4.589
R72696 out.n11878 out.n11877 4.589
R72697 out.n13986 out.n13985 4.589
R72698 out.n10611 out.n10610 4.589
R72699 out.n14318 out.n14317 4.589
R72700 out.n5005 out.n5004 4.589
R72701 out.n13118 out.n13117 4.582
R72702 out.n12742 out.n12741 4.582
R72703 out.n12253 out.n12252 4.582
R72704 out.n13576 out.n13575 4.582
R72705 out.n11422 out.n11421 4.582
R72706 out.n10995 out.n10994 4.582
R72707 out.n11833 out.n11832 4.582
R72708 out.n14031 out.n14030 4.582
R72709 out.n10566 out.n10565 4.582
R72710 out.n14323 out.n14322 4.582
R72711 out.n5010 out.n5009 4.582
R72712 out.n10218 out.n10217 4.574
R72713 out.n10085 out.n10084 4.567
R72714 out.n5288 out.n5287 4.567
R72715 out.n12573 out.n12572 4.56
R72716 out.n13406 out.n13405 4.56
R72717 out.n13861 out.n13860 4.56
R72718 out.n14229 out.n14228 4.56
R72719 out.n10146 out.n10081 4.558
R72720 out.n10167 out.n10077 4.558
R72721 out.n10165 out.n10080 4.558
R72722 out.n10214 out.n10208 4.558
R72723 out.n10214 out.n10213 4.558
R72724 out.n10229 out.n10059 4.558
R72725 out.n12994 out.n12993 4.558
R72726 out.n13079 out.n12877 4.558
R72727 out.n12568 out.n12567 4.558
R72728 out.n12794 out.n12415 4.558
R72729 out.n12129 out.n12128 4.558
R72730 out.n12214 out.n12010 4.558
R72731 out.n13401 out.n13400 4.558
R72732 out.n13628 out.n13260 4.558
R72733 out.n11306 out.n11305 4.558
R72734 out.n11388 out.n11175 4.558
R72735 out.n10876 out.n10875 4.558
R72736 out.n10961 out.n10752 4.558
R72737 out.n11709 out.n11708 4.558
R72738 out.n11794 out.n11592 4.558
R72739 out.n13856 out.n13855 4.558
R72740 out.n14083 out.n13715 4.558
R72741 out.n10442 out.n10441 4.558
R72742 out.n10527 out.n10325 4.558
R72743 out.n14423 out.n14370 4.558
R72744 out.n14219 out.n14218 4.558
R72745 out.n1006 out.n1005 4.558
R72746 out.n5097 out.n5059 4.558
R72747 out.n2744 out.n2743 4.558
R72748 out.n2849 out.n2848 4.558
R72749 out.n1517 out.n1516 4.558
R72750 out.n5407 out.n5402 4.558
R72751 out.n1146 out.n1145 4.558
R72752 out.n5357 out.n5183 4.558
R72753 out.n5359 out.n5180 4.558
R72754 out.n5247 out.n5196 4.558
R72755 out.n1220 out.n1219 4.558
R72756 out.n2156 out.n2155 4.558
R72757 out.n6476 out.n6471 4.558
R72758 out.n1873 out.n1872 4.558
R72759 out.n1973 out.n1972 4.558
R72760 out.n1600 out.n1599 4.558
R72761 out.n6171 out.n5881 4.558
R72762 out.n5894 out.n5889 4.558
R72763 out.n1648 out.n1647 4.558
R72764 out.n1753 out.n1752 4.558
R72765 out.n2364 out.n2363 4.558
R72766 out.n7268 out.n7263 4.558
R72767 out.n7216 out.n7029 4.558
R72768 out.n7046 out.n7041 4.558
R72769 out.n2493 out.n2492 4.558
R72770 out.n2701 out.n2700 4.558
R72771 out.n7549 out.n7544 4.558
R72772 out.n9445 out.n9429 4.531
R72773 out.n12999 out.n12998 4.517
R72774 out.n12134 out.n12133 4.517
R72775 out.n11177 out.n11176 4.517
R72776 out.n10881 out.n10880 4.517
R72777 out.n11714 out.n11713 4.517
R72778 out.n10447 out.n10446 4.517
R72779 out.n1016 out.n1015 4.517
R72780 out.n6094 out.n6093 4.517
R72781 out.n9445 out.n9428 4.5
R72782 out.n9443 out.n9442 4.5
R72783 out.n9445 out.n9430 4.5
R72784 out.n9432 out.n9430 4.5
R72785 out.n9443 out.n9430 4.5
R72786 out.n9443 out.n9426 4.5
R72787 out.n9432 out.n9426 4.5
R72788 out.n9445 out.n9426 4.5
R72789 out.n9445 out.n9444 4.5
R72790 out.n9444 out.n9432 4.5
R72791 out.n9444 out.n9443 4.5
R72792 out.n9432 out.n9428 4.5
R72793 out.n9443 out.n9428 4.5
R72794 out.n10113 out.n10112 4.5
R72795 out.n10088 out.n10087 4.5
R72796 out.n10128 out.n10127 4.5
R72797 out.n10131 out.n10095 4.5
R72798 out.n10139 out.n10138 4.5
R72799 out.n10164 out.n10163 4.5
R72800 out.n10158 out.n10157 4.5
R72801 out.n10153 out.n10152 4.5
R72802 out.n10066 out.n10065 4.5
R72803 out.n10186 out.n10185 4.5
R72804 out.n10204 out.n10203 4.5
R72805 out.n10225 out.n10224 4.5
R72806 out.n10221 out.n10220 4.5
R72807 out.n10270 out.n10269 4.5
R72808 out.n10262 out.n10261 4.5
R72809 out.n10245 out.n10244 4.5
R72810 out.n10238 out.n10237 4.5
R72811 out.n12838 out.n12837 4.5
R72812 out.n12940 out.n12939 4.5
R72813 out.n12952 out.n12951 4.5
R72814 out.n12960 out.n12959 4.5
R72815 out.n12967 out.n12966 4.5
R72816 out.n12888 out.n12887 4.5
R72817 out.n12882 out.n12881 4.5
R72818 out.n12982 out.n12981 4.5
R72819 out.n12990 out.n12989 4.5
R72820 out.n13011 out.n13010 4.5
R72821 out.n13056 out.n13055 4.5
R72822 out.n13067 out.n13066 4.5
R72823 out.n13078 out.n13077 4.5
R72824 out.n12868 out.n12867 4.5
R72825 out.n13090 out.n13089 4.5
R72826 out.n13110 out.n13109 4.5
R72827 out.n13121 out.n13120 4.5
R72828 out.n13166 out.n13165 4.5
R72829 out.n13177 out.n13176 4.5
R72830 out.n13190 out.n13189 4.5
R72831 out.n13202 out.n13201 4.5
R72832 out.n13211 out.n13210 4.5
R72833 out.n13223 out.n13222 4.5
R72834 out.n12815 out.n12814 4.5
R72835 out.n12465 out.n12464 4.5
R72836 out.n12514 out.n12513 4.5
R72837 out.n12525 out.n12524 4.5
R72838 out.n12534 out.n12533 4.5
R72839 out.n12540 out.n12539 4.5
R72840 out.n12451 out.n12450 4.5
R72841 out.n12445 out.n12444 4.5
R72842 out.n12556 out.n12555 4.5
R72843 out.n12565 out.n12564 4.5
R72844 out.n12576 out.n12575 4.5
R72845 out.n12587 out.n12586 4.5
R72846 out.n12634 out.n12633 4.5
R72847 out.n12645 out.n12644 4.5
R72848 out.n12656 out.n12655 4.5
R72849 out.n12434 out.n12433 4.5
R72850 out.n12428 out.n12427 4.5
R72851 out.n12425 out.n12424 4.5
R72852 out.n12689 out.n12688 4.5
R72853 out.n12700 out.n12699 4.5
R72854 out.n12745 out.n12744 4.5
R72855 out.n12756 out.n12755 4.5
R72856 out.n12779 out.n12778 4.5
R72857 out.n12788 out.n12787 4.5
R72858 out.n12797 out.n12796 4.5
R72859 out.n12379 out.n12378 4.5
R72860 out.n12075 out.n12074 4.5
R72861 out.n12087 out.n12086 4.5
R72862 out.n12095 out.n12094 4.5
R72863 out.n12102 out.n12101 4.5
R72864 out.n12021 out.n12020 4.5
R72865 out.n12015 out.n12014 4.5
R72866 out.n12117 out.n12116 4.5
R72867 out.n12125 out.n12124 4.5
R72868 out.n12146 out.n12145 4.5
R72869 out.n12191 out.n12190 4.5
R72870 out.n12202 out.n12201 4.5
R72871 out.n12213 out.n12212 4.5
R72872 out.n12001 out.n12000 4.5
R72873 out.n12225 out.n12224 4.5
R72874 out.n12245 out.n12244 4.5
R72875 out.n12256 out.n12255 4.5
R72876 out.n12301 out.n12300 4.5
R72877 out.n12312 out.n12311 4.5
R72878 out.n12325 out.n12324 4.5
R72879 out.n12337 out.n12336 4.5
R72880 out.n12346 out.n12345 4.5
R72881 out.n12358 out.n12357 4.5
R72882 out.n13654 out.n13653 4.5
R72883 out.n13661 out.n13660 4.5
R72884 out.n13347 out.n13346 4.5
R72885 out.n13358 out.n13357 4.5
R72886 out.n13367 out.n13366 4.5
R72887 out.n13373 out.n13372 4.5
R72888 out.n13295 out.n13294 4.5
R72889 out.n13289 out.n13288 4.5
R72890 out.n13389 out.n13388 4.5
R72891 out.n13398 out.n13397 4.5
R72892 out.n13409 out.n13408 4.5
R72893 out.n13420 out.n13419 4.5
R72894 out.n13467 out.n13466 4.5
R72895 out.n13478 out.n13477 4.5
R72896 out.n13489 out.n13488 4.5
R72897 out.n13278 out.n13277 4.5
R72898 out.n13272 out.n13271 4.5
R72899 out.n13269 out.n13268 4.5
R72900 out.n13523 out.n13522 4.5
R72901 out.n13534 out.n13533 4.5
R72902 out.n13579 out.n13578 4.5
R72903 out.n13590 out.n13589 4.5
R72904 out.n13613 out.n13612 4.5
R72905 out.n13622 out.n13621 4.5
R72906 out.n13631 out.n13630 4.5
R72907 out.n11547 out.n11546 4.5
R72908 out.n11252 out.n11251 4.5
R72909 out.n11264 out.n11263 4.5
R72910 out.n11272 out.n11271 4.5
R72911 out.n11279 out.n11278 4.5
R72912 out.n11189 out.n11188 4.5
R72913 out.n11183 out.n11182 4.5
R72914 out.n11294 out.n11293 4.5
R72915 out.n11302 out.n11301 4.5
R72916 out.n11320 out.n11319 4.5
R72917 out.n11365 out.n11364 4.5
R72918 out.n11376 out.n11375 4.5
R72919 out.n11387 out.n11386 4.5
R72920 out.n11166 out.n11165 4.5
R72921 out.n11399 out.n11398 4.5
R72922 out.n11157 out.n11156 4.5
R72923 out.n11425 out.n11424 4.5
R72924 out.n11470 out.n11469 4.5
R72925 out.n11481 out.n11480 4.5
R72926 out.n11494 out.n11493 4.5
R72927 out.n11506 out.n11505 4.5
R72928 out.n11515 out.n11514 4.5
R72929 out.n11527 out.n11526 4.5
R72930 out.n11123 out.n11122 4.5
R72931 out.n10822 out.n10821 4.5
R72932 out.n10834 out.n10833 4.5
R72933 out.n10842 out.n10841 4.5
R72934 out.n10849 out.n10848 4.5
R72935 out.n10763 out.n10762 4.5
R72936 out.n10757 out.n10756 4.5
R72937 out.n10864 out.n10863 4.5
R72938 out.n10872 out.n10871 4.5
R72939 out.n10893 out.n10892 4.5
R72940 out.n10938 out.n10937 4.5
R72941 out.n10949 out.n10948 4.5
R72942 out.n10960 out.n10959 4.5
R72943 out.n10743 out.n10742 4.5
R72944 out.n10972 out.n10971 4.5
R72945 out.n10734 out.n10733 4.5
R72946 out.n10998 out.n10997 4.5
R72947 out.n11043 out.n11042 4.5
R72948 out.n11054 out.n11053 4.5
R72949 out.n11067 out.n11066 4.5
R72950 out.n11079 out.n11078 4.5
R72951 out.n11088 out.n11087 4.5
R72952 out.n11100 out.n11099 4.5
R72953 out.n11959 out.n11958 4.5
R72954 out.n11655 out.n11654 4.5
R72955 out.n11667 out.n11666 4.5
R72956 out.n11675 out.n11674 4.5
R72957 out.n11682 out.n11681 4.5
R72958 out.n11603 out.n11602 4.5
R72959 out.n11597 out.n11596 4.5
R72960 out.n11697 out.n11696 4.5
R72961 out.n11705 out.n11704 4.5
R72962 out.n11726 out.n11725 4.5
R72963 out.n11771 out.n11770 4.5
R72964 out.n11782 out.n11781 4.5
R72965 out.n11793 out.n11792 4.5
R72966 out.n11583 out.n11582 4.5
R72967 out.n11805 out.n11804 4.5
R72968 out.n11825 out.n11824 4.5
R72969 out.n11836 out.n11835 4.5
R72970 out.n11881 out.n11880 4.5
R72971 out.n11892 out.n11891 4.5
R72972 out.n11905 out.n11904 4.5
R72973 out.n11917 out.n11916 4.5
R72974 out.n11926 out.n11925 4.5
R72975 out.n11938 out.n11937 4.5
R72976 out.n13687 out.n13686 4.5
R72977 out.n13694 out.n13693 4.5
R72978 out.n13802 out.n13801 4.5
R72979 out.n13813 out.n13812 4.5
R72980 out.n13822 out.n13821 4.5
R72981 out.n13828 out.n13827 4.5
R72982 out.n13750 out.n13749 4.5
R72983 out.n13744 out.n13743 4.5
R72984 out.n13844 out.n13843 4.5
R72985 out.n13853 out.n13852 4.5
R72986 out.n13864 out.n13863 4.5
R72987 out.n13875 out.n13874 4.5
R72988 out.n13922 out.n13921 4.5
R72989 out.n13933 out.n13932 4.5
R72990 out.n13944 out.n13943 4.5
R72991 out.n13733 out.n13732 4.5
R72992 out.n13727 out.n13726 4.5
R72993 out.n13724 out.n13723 4.5
R72994 out.n13978 out.n13977 4.5
R72995 out.n13989 out.n13988 4.5
R72996 out.n14034 out.n14033 4.5
R72997 out.n14045 out.n14044 4.5
R72998 out.n14068 out.n14067 4.5
R72999 out.n14077 out.n14076 4.5
R73000 out.n14086 out.n14085 4.5
R73001 out.n10692 out.n10691 4.5
R73002 out.n10388 out.n10387 4.5
R73003 out.n10400 out.n10399 4.5
R73004 out.n10408 out.n10407 4.5
R73005 out.n10415 out.n10414 4.5
R73006 out.n10336 out.n10335 4.5
R73007 out.n10330 out.n10329 4.5
R73008 out.n10430 out.n10429 4.5
R73009 out.n10438 out.n10437 4.5
R73010 out.n10459 out.n10458 4.5
R73011 out.n10504 out.n10503 4.5
R73012 out.n10515 out.n10514 4.5
R73013 out.n10526 out.n10525 4.5
R73014 out.n10316 out.n10315 4.5
R73015 out.n10538 out.n10537 4.5
R73016 out.n10558 out.n10557 4.5
R73017 out.n10569 out.n10568 4.5
R73018 out.n10614 out.n10613 4.5
R73019 out.n10625 out.n10624 4.5
R73020 out.n10638 out.n10637 4.5
R73021 out.n10650 out.n10649 4.5
R73022 out.n10659 out.n10658 4.5
R73023 out.n10671 out.n10670 4.5
R73024 out.n14165 out.n14164 4.5
R73025 out.n14386 out.n14385 4.5
R73026 out.n14379 out.n14378 4.5
R73027 out.n14422 out.n14421 4.5
R73028 out.n14360 out.n14359 4.5
R73029 out.n14349 out.n14348 4.5
R73030 out.n14335 out.n14334 4.5
R73031 out.n14326 out.n14325 4.5
R73032 out.n14321 out.n14320 4.5
R73033 out.n14312 out.n14311 4.5
R73034 out.n14303 out.n14302 4.5
R73035 out.n14292 out.n14291 4.5
R73036 out.n14281 out.n14280 4.5
R73037 out.n14485 out.n14484 4.5
R73038 out.n14266 out.n14265 4.5
R73039 out.n14257 out.n14256 4.5
R73040 out.n14241 out.n14240 4.5
R73041 out.n14232 out.n14231 4.5
R73042 out.n14222 out.n14221 4.5
R73043 out.n14214 out.n14213 4.5
R73044 out.n14203 out.n14202 4.5
R73045 out.n14196 out.n14195 4.5
R73046 out.n14533 out.n14532 4.5
R73047 out.n14542 out.n14541 4.5
R73048 out.n14185 out.n14184 4.5
R73049 out.n14555 out.n14554 4.5
R73050 out.n14560 out.n14559 4.5
R73051 out.n10282 out.n10281 4.5
R73052 out.n13234 out.n13233 4.5
R73053 out.n12408 out.n12407 4.5
R73054 out.n11982 out.n11981 4.5
R73055 out.n13253 out.n13252 4.5
R73056 out.n11142 out.n11141 4.5
R73057 out.n10719 out.n10718 4.5
R73058 out.n11565 out.n11564 4.5
R73059 out.n13708 out.n13707 4.5
R73060 out.n10298 out.n10297 4.5
R73061 out.n942 out.n941 4.5
R73062 out.n970 out.n969 4.5
R73063 out.n976 out.n975 4.5
R73064 out.n1074 out.n1073 4.5
R73065 out.n1066 out.n1065 4.5
R73066 out.n984 out.n983 4.5
R73067 out.n991 out.n990 4.5
R73068 out.n1000 out.n999 4.5
R73069 out.n1009 out.n1008 4.5
R73070 out.n1026 out.n1025 4.5
R73071 out.n5075 out.n5074 4.5
R73072 out.n5068 out.n5067 4.5
R73073 out.n5096 out.n5095 4.5
R73074 out.n5049 out.n5048 4.5
R73075 out.n5038 out.n5037 4.5
R73076 out.n5022 out.n5021 4.5
R73077 out.n5013 out.n5012 4.5
R73078 out.n5008 out.n5007 4.5
R73079 out.n4999 out.n4998 4.5
R73080 out.n4990 out.n4989 4.5
R73081 out.n4978 out.n4977 4.5
R73082 out.n4967 out.n4966 4.5
R73083 out.n5159 out.n5158 4.5
R73084 out.n5167 out.n5166 4.5
R73085 out.n5849 out.n5848 4.5
R73086 out.n5638 out.n5637 4.5
R73087 out.n5822 out.n5821 4.5
R73088 out.n5831 out.n5830 4.5
R73089 out.n5813 out.n5812 4.5
R73090 out.n5751 out.n5750 4.5
R73091 out.n5647 out.n5646 4.5
R73092 out.n5738 out.n5737 4.5
R73093 out.n5726 out.n5725 4.5
R73094 out.n5653 out.n5652 4.5
R73095 out.n5713 out.n5712 4.5
R73096 out.n5691 out.n5690 4.5
R73097 out.n5699 out.n5698 4.5
R73098 out.n5706 out.n5705 4.5
R73099 out.n5683 out.n5682 4.5
R73100 out.n2859 out.n2858 4.5
R73101 out.n2852 out.n2851 4.5
R73102 out.n2845 out.n2844 4.5
R73103 out.n2835 out.n2834 4.5
R73104 out.n2827 out.n2826 4.5
R73105 out.n2821 out.n2820 4.5
R73106 out.n2812 out.n2811 4.5
R73107 out.n2780 out.n2779 4.5
R73108 out.n2789 out.n2788 4.5
R73109 out.n2796 out.n2795 4.5
R73110 out.n2807 out.n2806 4.5
R73111 out.n2940 out.n2939 4.5
R73112 out.n5395 out.n5394 4.5
R73113 out.n5578 out.n5577 4.5
R73114 out.n5587 out.n5586 4.5
R73115 out.n5567 out.n5566 4.5
R73116 out.n5556 out.n5555 4.5
R73117 out.n5507 out.n5506 4.5
R73118 out.n5498 out.n5497 4.5
R73119 out.n5406 out.n5405 4.5
R73120 out.n5485 out.n5484 4.5
R73121 out.n5412 out.n5411 4.5
R73122 out.n5418 out.n5417 4.5
R73123 out.n5469 out.n5468 4.5
R73124 out.n5452 out.n5451 4.5
R73125 out.n5429 out.n5428 4.5
R73126 out.n1419 out.n1418 4.5
R73127 out.n1412 out.n1411 4.5
R73128 out.n1403 out.n1402 4.5
R73129 out.n1374 out.n1373 4.5
R73130 out.n1381 out.n1380 4.5
R73131 out.n1388 out.n1387 4.5
R73132 out.n1498 out.n1497 4.5
R73133 out.n1529 out.n1528 4.5
R73134 out.n5177 out.n5176 4.5
R73135 out.n5362 out.n5361 4.5
R73136 out.n5356 out.n5355 4.5
R73137 out.n5347 out.n5346 4.5
R73138 out.n5291 out.n5290 4.5
R73139 out.n5269 out.n5268 4.5
R73140 out.n5260 out.n5259 4.5
R73141 out.n5189 out.n5188 4.5
R73142 out.n5239 out.n5238 4.5
R73143 out.n5246 out.n5245 4.5
R73144 out.n5230 out.n5229 4.5
R73145 out.n1223 out.n1222 4.5
R73146 out.n1216 out.n1215 4.5
R73147 out.n1206 out.n1205 4.5
R73148 out.n1198 out.n1197 4.5
R73149 out.n1191 out.n1190 4.5
R73150 out.n1186 out.n1185 4.5
R73151 out.n1289 out.n1288 4.5
R73152 out.n1281 out.n1280 4.5
R73153 out.n1274 out.n1273 4.5
R73154 out.n1334 out.n1333 4.5
R73155 out.n6454 out.n6453 4.5
R73156 out.n6732 out.n6731 4.5
R73157 out.n6741 out.n6740 4.5
R73158 out.n6721 out.n6720 4.5
R73159 out.n6710 out.n6709 4.5
R73160 out.n6671 out.n6670 4.5
R73161 out.n6662 out.n6661 4.5
R73162 out.n6475 out.n6474 4.5
R73163 out.n6649 out.n6648 4.5
R73164 out.n6481 out.n6480 4.5
R73165 out.n6487 out.n6486 4.5
R73166 out.n6633 out.n6632 4.5
R73167 out.n6497 out.n6496 4.5
R73168 out.n6615 out.n6614 4.5
R73169 out.n6523 out.n6522 4.5
R73170 out.n6529 out.n6528 4.5
R73171 out.n6538 out.n6537 4.5
R73172 out.n2136 out.n2135 4.5
R73173 out.n2103 out.n2102 4.5
R73174 out.n2110 out.n2109 4.5
R73175 out.n2121 out.n2120 4.5
R73176 out.n2167 out.n2166 4.5
R73177 out.n6421 out.n6420 4.5
R73178 out.n6210 out.n6209 4.5
R73179 out.n6394 out.n6393 4.5
R73180 out.n6403 out.n6402 4.5
R73181 out.n6385 out.n6384 4.5
R73182 out.n6328 out.n6327 4.5
R73183 out.n6224 out.n6223 4.5
R73184 out.n6315 out.n6314 4.5
R73185 out.n6303 out.n6302 4.5
R73186 out.n6230 out.n6229 4.5
R73187 out.n6290 out.n6289 4.5
R73188 out.n6268 out.n6267 4.5
R73189 out.n6276 out.n6275 4.5
R73190 out.n6283 out.n6282 4.5
R73191 out.n6260 out.n6259 4.5
R73192 out.n1983 out.n1982 4.5
R73193 out.n1976 out.n1975 4.5
R73194 out.n1969 out.n1968 4.5
R73195 out.n1959 out.n1958 4.5
R73196 out.n1951 out.n1950 4.5
R73197 out.n1945 out.n1944 4.5
R73198 out.n1936 out.n1935 4.5
R73199 out.n1904 out.n1903 4.5
R73200 out.n1913 out.n1912 4.5
R73201 out.n1920 out.n1919 4.5
R73202 out.n1931 out.n1930 4.5
R73203 out.n2069 out.n2068 4.5
R73204 out.n5877 out.n5876 4.5
R73205 out.n6170 out.n6169 4.5
R73206 out.n6159 out.n6158 4.5
R73207 out.n6148 out.n6147 4.5
R73208 out.n6108 out.n6107 4.5
R73209 out.n5893 out.n5892 4.5
R73210 out.n6085 out.n6084 4.5
R73211 out.n5899 out.n5898 4.5
R73212 out.n6072 out.n6071 4.5
R73213 out.n6057 out.n6056 4.5
R73214 out.n6065 out.n6064 4.5
R73215 out.n6049 out.n6048 4.5
R73216 out.n6037 out.n6036 4.5
R73217 out.n5920 out.n5919 4.5
R73218 out.n5928 out.n5927 4.5
R73219 out.n5983 out.n5982 4.5
R73220 out.n5934 out.n5933 4.5
R73221 out.n5970 out.n5969 4.5
R73222 out.n5962 out.n5961 4.5
R73223 out.n1558 out.n1557 4.5
R73224 out.n1563 out.n1562 4.5
R73225 out.n1568 out.n1567 4.5
R73226 out.n5941 out.n5940 4.5
R73227 out.n5947 out.n5946 4.5
R73228 out.n1610 out.n1609 4.5
R73229 out.n6983 out.n6982 4.5
R73230 out.n6772 out.n6771 4.5
R73231 out.n6956 out.n6955 4.5
R73232 out.n6965 out.n6964 4.5
R73233 out.n6947 out.n6946 4.5
R73234 out.n6885 out.n6884 4.5
R73235 out.n6781 out.n6780 4.5
R73236 out.n6872 out.n6871 4.5
R73237 out.n6860 out.n6859 4.5
R73238 out.n6787 out.n6786 4.5
R73239 out.n6847 out.n6846 4.5
R73240 out.n6825 out.n6824 4.5
R73241 out.n6833 out.n6832 4.5
R73242 out.n6840 out.n6839 4.5
R73243 out.n6817 out.n6816 4.5
R73244 out.n1763 out.n1762 4.5
R73245 out.n1756 out.n1755 4.5
R73246 out.n1749 out.n1748 4.5
R73247 out.n1739 out.n1738 4.5
R73248 out.n1731 out.n1730 4.5
R73249 out.n1725 out.n1724 4.5
R73250 out.n1716 out.n1715 4.5
R73251 out.n1684 out.n1683 4.5
R73252 out.n1693 out.n1692 4.5
R73253 out.n1700 out.n1699 4.5
R73254 out.n1711 out.n1710 4.5
R73255 out.n1844 out.n1843 4.5
R73256 out.n7256 out.n7255 4.5
R73257 out.n7436 out.n7435 4.5
R73258 out.n7445 out.n7444 4.5
R73259 out.n7425 out.n7424 4.5
R73260 out.n7414 out.n7413 4.5
R73261 out.n7365 out.n7364 4.5
R73262 out.n7356 out.n7355 4.5
R73263 out.n7267 out.n7266 4.5
R73264 out.n7343 out.n7342 4.5
R73265 out.n7273 out.n7272 4.5
R73266 out.n7279 out.n7278 4.5
R73267 out.n7327 out.n7326 4.5
R73268 out.n7310 out.n7309 4.5
R73269 out.n7290 out.n7289 4.5
R73270 out.n2263 out.n2262 4.5
R73271 out.n2256 out.n2255 4.5
R73272 out.n2247 out.n2246 4.5
R73273 out.n2218 out.n2217 4.5
R73274 out.n2225 out.n2224 4.5
R73275 out.n2232 out.n2231 4.5
R73276 out.n2345 out.n2344 4.5
R73277 out.n2376 out.n2375 4.5
R73278 out.n7229 out.n7228 4.5
R73279 out.n7022 out.n7021 4.5
R73280 out.n7206 out.n7205 4.5
R73281 out.n7215 out.n7214 4.5
R73282 out.n7197 out.n7196 4.5
R73283 out.n7045 out.n7044 4.5
R73284 out.n7134 out.n7133 4.5
R73285 out.n7122 out.n7121 4.5
R73286 out.n7051 out.n7050 4.5
R73287 out.n7109 out.n7108 4.5
R73288 out.n7087 out.n7086 4.5
R73289 out.n7095 out.n7094 4.5
R73290 out.n7102 out.n7101 4.5
R73291 out.n7079 out.n7078 4.5
R73292 out.n2475 out.n2474 4.5
R73293 out.n2468 out.n2467 4.5
R73294 out.n2459 out.n2458 4.5
R73295 out.n2427 out.n2426 4.5
R73296 out.n2435 out.n2434 4.5
R73297 out.n2441 out.n2440 4.5
R73298 out.n2454 out.n2453 4.5
R73299 out.n2592 out.n2591 4.5
R73300 out.n7483 out.n7482 4.5
R73301 out.n7777 out.n7776 4.5
R73302 out.n7786 out.n7785 4.5
R73303 out.n7768 out.n7767 4.5
R73304 out.n7711 out.n7710 4.5
R73305 out.n7497 out.n7496 4.5
R73306 out.n7506 out.n7505 4.5
R73307 out.n7516 out.n7515 4.5
R73308 out.n7523 out.n7522 4.5
R73309 out.n7693 out.n7692 4.5
R73310 out.n7672 out.n7671 4.5
R73311 out.n7680 out.n7679 4.5
R73312 out.n7687 out.n7686 4.5
R73313 out.n7664 out.n7663 4.5
R73314 out.n7620 out.n7619 4.5
R73315 out.n7548 out.n7547 4.5
R73316 out.n7557 out.n7556 4.5
R73317 out.n7567 out.n7566 4.5
R73318 out.n7574 out.n7573 4.5
R73319 out.n7601 out.n7600 4.5
R73320 out.n7581 out.n7580 4.5
R73321 out.n2644 out.n2643 4.5
R73322 out.n2652 out.n2651 4.5
R73323 out.n2658 out.n2657 4.5
R73324 out.n2661 out.n2660 4.5
R73325 out.n2711 out.n2710 4.5
R73326 out.n5601 out.n5600 4.5
R73327 out.n5600 out.n5599 4.5
R73328 out.n7813 out.n7812 4.5
R73329 out.n7459 out.n7458 4.5
R73330 out.n7458 out.n7457 4.5
R73331 out.n6756 out.n6755 4.5
R73332 out.n6434 out.n6428 4.5
R73333 out.n6433 out.n6432 4.5
R73334 out.n6432 out.n6431 4.5
R73335 out.n6996 out.n6990 4.5
R73336 out.n6995 out.n6994 4.5
R73337 out.n6994 out.n6993 4.5
R73338 out.n7460 out.n7454 4.5
R73339 out.n7242 out.n7236 4.5
R73340 out.n7241 out.n7240 4.5
R73341 out.n7240 out.n7239 4.5
R73342 out.n5857 out.n5856 4.5
R73343 out.n5633 out.n5632 4.5
R73344 out.n5632 out.n5631 4.5
R73345 out.n5602 out.n5596 4.5
R73346 out.n5386 out.n5173 4.5
R73347 out.n5385 out.n5384 4.5
R73348 out.n5384 out.n5383 4.5
R73349 out.n5169 out.n5168 4.5
R73350 out.n1128 out.n1127 4.5
R73351 out.n10178 out.n10177 4.47
R73352 out.n12835 out.n12834 4.384
R73353 out.n12376 out.n12375 4.384
R73354 out.n11196 out.n11195 4.384
R73355 out.n11120 out.n11119 4.384
R73356 out.n11956 out.n11955 4.384
R73357 out.n10689 out.n10688 4.384
R73358 out.n1116 out.n1115 4.384
R73359 out.n939 out.n938 4.384
R73360 out.n5648 out.n5643 4.384
R73361 out.n1445 out.n1444 4.384
R73362 out.n1439 out.n1438 4.384
R73363 out.n6565 out.n6564 4.384
R73364 out.n6510 out.n6509 4.384
R73365 out.n6225 out.n6220 4.384
R73366 out.n5921 out.n5916 4.384
R73367 out.n5929 out.n5924 4.384
R73368 out.n6782 out.n6777 4.384
R73369 out.n2289 out.n2288 4.384
R73370 out.n2283 out.n2282 4.384
R73371 out.n2407 out.n2406 4.384
R73372 out.n7498 out.n7493 4.384
R73373 out.n2434 out.n2433 4.363
R73374 out.n10232 out.n10231 4.328
R73375 out.n5846 out.n5845 4.328
R73376 out.n6418 out.n6417 4.328
R73377 out.n6980 out.n6979 4.328
R73378 out.n7801 out.n7800 4.328
R73379 out.n10117 out.n10116 4.326
R73380 out.n5273 out.n5272 4.326
R73381 out.n12458 out.n12457 4.223
R73382 out.n13651 out.n13650 4.223
R73383 out.n13684 out.n13683 4.223
R73384 out.n2750 out.n2749 4.223
R73385 out.n5499 out.n5494 4.223
R73386 out.n1152 out.n1151 4.223
R73387 out.n6663 out.n6658 4.223
R73388 out.n1879 out.n1878 4.223
R73389 out.n1654 out.n1653 4.223
R73390 out.n7357 out.n7352 4.223
R73391 out.n2498 out.n2497 4.223
R73392 out.n2695 out.n2694 4.223
R73393 out.n5848 out.n5846 4.162
R73394 out.n6420 out.n6418 4.162
R73395 out.n6982 out.n6980 4.162
R73396 out.n10112 out.n10110 4.154
R73397 out.n13089 out.n13087 4.154
R73398 out.n12778 out.n12777 4.154
R73399 out.n12224 out.n12222 4.154
R73400 out.n13612 out.n13611 4.154
R73401 out.n11398 out.n11396 4.154
R73402 out.n10971 out.n10969 4.154
R73403 out.n11804 out.n11802 4.154
R73404 out.n14067 out.n14066 4.154
R73405 out.n10537 out.n10535 4.154
R73406 out.n5037 out.n5035 4.154
R73407 out.n5268 out.n5266 4.154
R73408 out.n2788 out.n2786 4.141
R73409 out.n1387 out.n1385 4.141
R73410 out.n2109 out.n2107 4.141
R73411 out.n1912 out.n1910 4.141
R73412 out.n1692 out.n1690 4.141
R73413 out.n2231 out.n2229 4.141
R73414 out.n2651 out.n2649 4.141
R73415 out.n2788 out.n2787 3.987
R73416 out.n1912 out.n1911 3.987
R73417 out.n1692 out.n1691 3.987
R73418 out.n2651 out.n2650 3.987
R73419 out.n10104 out.n10103 3.951
R73420 out.n5257 out.n5256 3.951
R73421 out.n7226 out.n7225 3.951
R73422 out.n10157 out.n10156 3.95
R73423 out.n12552 out.n12551 3.95
R73424 out.n13385 out.n13384 3.95
R73425 out.n13840 out.n13839 3.95
R73426 out.n14211 out.n14210 3.95
R73427 out.n1151 out.n1150 3.879
R73428 out.n2497 out.n2496 3.879
R73429 out.n5301 out.n5300 3.843
R73430 out.n12584 out.n12583 3.836
R73431 out.n13417 out.n13416 3.836
R73432 out.n13872 out.n13871 3.836
R73433 out.n14238 out.n14237 3.836
R73434 out.n13008 out.n13007 3.829
R73435 out.n12143 out.n12142 3.829
R73436 out.n11317 out.n11316 3.829
R73437 out.n10890 out.n10889 3.829
R73438 out.n11723 out.n11722 3.829
R73439 out.n10456 out.n10455 3.829
R73440 out.n14162 out.n14161 3.829
R73441 out.n1023 out.n1022 3.829
R73442 out.n6105 out.n6104 3.829
R73443 out.n5748 out.n5747 3.821
R73444 out.n6325 out.n6324 3.821
R73445 out.n6882 out.n6881 3.821
R73446 out.n7708 out.n7707 3.821
R73447 out.n1228 out.n1227 3.814
R73448 out.n7144 out.n7143 3.814
R73449 out.n1541 out.n1540 3.77
R73450 out.n13108 out.n13107 3.764
R73451 out.n12574 out.n12573 3.764
R73452 out.n12754 out.n12753 3.764
R73453 out.n12243 out.n12242 3.764
R73454 out.n13407 out.n13406 3.764
R73455 out.n13588 out.n13587 3.764
R73456 out.n11155 out.n11154 3.764
R73457 out.n10732 out.n10731 3.764
R73458 out.n11823 out.n11822 3.764
R73459 out.n13862 out.n13861 3.764
R73460 out.n14043 out.n14042 3.764
R73461 out.n10556 out.n10555 3.764
R73462 out.n14333 out.n14332 3.764
R73463 out.n14230 out.n14229 3.764
R73464 out.n5020 out.n5019 3.764
R73465 out.n2734 out.n2732 3.764
R73466 out.n1429 out.n1427 3.764
R73467 out.n1229 out.n1228 3.764
R73468 out.n6517 out.n6515 3.764
R73469 out.n1863 out.n1861 3.764
R73470 out.n1557 out.n1555 3.764
R73471 out.n1638 out.n1636 3.764
R73472 out.n2273 out.n2271 3.764
R73473 out.n7145 out.n7144 3.764
R73474 out.n2434 out.n2432 3.764
R73475 out.n10211 out.n10209 3.686
R73476 out.n2826 out.n2824 3.624
R73477 out.n5411 out.n5409 3.624
R73478 out.n1418 out.n1416 3.624
R73479 out.n1373 out.n1372 3.624
R73480 out.n6480 out.n6478 3.624
R73481 out.n6522 out.n6520 3.624
R73482 out.n2135 out.n2134 3.624
R73483 out.n1950 out.n1948 3.624
R73484 out.n5933 out.n5931 3.624
R73485 out.n1730 out.n1728 3.624
R73486 out.n7272 out.n7270 3.624
R73487 out.n2262 out.n2260 3.624
R73488 out.n2217 out.n2216 3.624
R73489 out.n2474 out.n2472 3.624
R73490 out.n7573 out.n7571 3.624
R73491 out.n1562 out.n1561 3.611
R73492 out.n10185 out.n10182 3.573
R73493 out.n12979 out.n12978 3.573
R73494 out.n12114 out.n12113 3.573
R73495 out.n11291 out.n11290 3.573
R73496 out.n10861 out.n10860 3.573
R73497 out.n11694 out.n11693 3.573
R73498 out.n10427 out.n10426 3.573
R73499 out.n997 out.n996 3.573
R73500 out.n6082 out.n6081 3.573
R73501 out.n5734 out.n5733 3.572
R73502 out.n6311 out.n6310 3.572
R73503 out.n6868 out.n6867 3.572
R73504 out.n7502 out.n7501 3.572
R73505 out.n1444 out.n1443 3.565
R73506 out.n6564 out.n6563 3.565
R73507 out.n2288 out.n2287 3.565
R73508 out.n12981 out.n12979 3.416
R73509 out.n12116 out.n12114 3.416
R73510 out.n11293 out.n11291 3.416
R73511 out.n10863 out.n10861 3.416
R73512 out.n11696 out.n11694 3.416
R73513 out.n10429 out.n10427 3.416
R73514 out.n999 out.n997 3.416
R73515 out.n1143 out.n1142 3.416
R73516 out.n5259 out.n5257 3.416
R73517 out.n6084 out.n6082 3.416
R73518 out.n7228 out.n7226 3.416
R73519 out.n2490 out.n2489 3.416
R73520 out.n5402 out.n5401 3.388
R73521 out.n6471 out.n6470 3.388
R73522 out.n7263 out.n7262 3.388
R73523 out.n2779 out.n2777 3.388
R73524 out.n1380 out.n1378 3.388
R73525 out.n2102 out.n2100 3.388
R73526 out.n1903 out.n1901 3.388
R73527 out.n1539 out.n1538 3.388
R73528 out.n5946 out.n5945 3.388
R73529 out.n1683 out.n1681 3.388
R73530 out.n2224 out.n2222 3.388
R73531 out.n2392 out.n2390 3.388
R73532 out.n2453 out.n2452 3.388
R73533 out.n2643 out.n2641 3.388
R73534 out.n1115 out.n1114 3.354
R73535 out.n5924 out.n5923 3.354
R73536 out.n2426 out.n2425 3.247
R73537 out.n5723 out.n5722 3.197
R73538 out.n6300 out.n6299 3.197
R73539 out.n6857 out.n6856 3.197
R73540 out.n7513 out.n7512 3.197
R73541 out.n1212 out.n1211 3.195
R73542 out.n7130 out.n7129 3.195
R73543 out.n10095 out.n10094 3.189
R73544 out.n10141 out.n10140 3.105
R73545 out.n10198 out.n10197 3.105
R73546 out.n12912 out.n12911 3.105
R73547 out.n13037 out.n13036 3.105
R73548 out.n13129 out.n13128 3.105
R73549 out.n13152 out.n13151 3.105
R73550 out.n12488 out.n12487 3.105
R73551 out.n12613 out.n12612 3.105
R73552 out.n12710 out.n12709 3.105
R73553 out.n12733 out.n12732 3.105
R73554 out.n12047 out.n12046 3.105
R73555 out.n12172 out.n12171 3.105
R73556 out.n12264 out.n12263 3.105
R73557 out.n12287 out.n12286 3.105
R73558 out.n13321 out.n13320 3.105
R73559 out.n13446 out.n13445 3.105
R73560 out.n13544 out.n13543 3.105
R73561 out.n13567 out.n13566 3.105
R73562 out.n11224 out.n11223 3.105
R73563 out.n11346 out.n11345 3.105
R73564 out.n11433 out.n11432 3.105
R73565 out.n11456 out.n11455 3.105
R73566 out.n10794 out.n10793 3.105
R73567 out.n10919 out.n10918 3.105
R73568 out.n11006 out.n11005 3.105
R73569 out.n11029 out.n11028 3.105
R73570 out.n11627 out.n11626 3.105
R73571 out.n11752 out.n11751 3.105
R73572 out.n11844 out.n11843 3.105
R73573 out.n11867 out.n11866 3.105
R73574 out.n13776 out.n13775 3.105
R73575 out.n13901 out.n13900 3.105
R73576 out.n13999 out.n13998 3.105
R73577 out.n14022 out.n14021 3.105
R73578 out.n10360 out.n10359 3.105
R73579 out.n10485 out.n10484 3.105
R73580 out.n10577 out.n10576 3.105
R73581 out.n10600 out.n10599 3.105
R73582 out.n14406 out.n14405 3.105
R73583 out.n14438 out.n14437 3.105
R73584 out.n14461 out.n14460 3.105
R73585 out.n14500 out.n14499 3.105
R73586 out.n1089 out.n1088 3.105
R73587 out.n1034 out.n1033 3.105
R73588 out.n5112 out.n5111 3.105
R73589 out.n5135 out.n5134 3.105
R73590 out.n5783 out.n5782 3.105
R73591 out.n2871 out.n2870 3.105
R73592 out.n5530 out.n5529 3.105
R73593 out.n1456 out.n1455 3.105
R73594 out.n5324 out.n5323 3.105
R73595 out.n5200 out.n5199 3.105
R73596 out.n1308 out.n1307 3.105
R73597 out.n6462 out.n6461 3.105
R73598 out.n6579 out.n6578 3.105
R73599 out.n6355 out.n6354 3.105
R73600 out.n1995 out.n1994 3.105
R73601 out.n6129 out.n6128 3.105
R73602 out.n5908 out.n5907 3.105
R73603 out.n6917 out.n6916 3.105
R73604 out.n1775 out.n1774 3.105
R73605 out.n7388 out.n7387 3.105
R73606 out.n2300 out.n2299 3.105
R73607 out.n7033 out.n7032 3.105
R73608 out.n2517 out.n2516 3.105
R73609 out.n7738 out.n7737 3.105
R73610 out.n7534 out.n7533 3.105
R73611 out.n1233 out.n1232 3.09
R73612 out.n7155 out.n7154 3.09
R73613 out.n12462 out.n12461 3.083
R73614 out.n13658 out.n13657 3.083
R73615 out.n13691 out.n13690 3.083
R73616 out.n5504 out.n5503 3.083
R73617 out.n6668 out.n6667 3.083
R73618 out.n7362 out.n7361 3.083
R73619 out.n12842 out.n12841 3.076
R73620 out.n12382 out.n12381 3.076
R73621 out.n11200 out.n11199 3.076
R73622 out.n10770 out.n10769 3.076
R73623 out.n11963 out.n11962 3.076
R73624 out.n10696 out.n10695 3.076
R73625 out.n1106 out.n1105 3.076
R73626 out.n5995 out.n5994 3.076
R73627 out.n2856 out.n2855 3.068
R73628 out.n1980 out.n1979 3.068
R73629 out.n1760 out.n1759 3.068
R73630 out.n7617 out.n7616 3.068
R73631 out.n12555 out.n12553 3.033
R73632 out.n13388 out.n13386 3.033
R73633 out.n13843 out.n13841 3.033
R73634 out.n14213 out.n14212 3.033
R73635 out.n5737 out.n5735 3.033
R73636 out.n6314 out.n6312 3.033
R73637 out.n6871 out.n6869 3.033
R73638 out.n7505 out.n7503 3.033
R73639 out.n10134 out.n10133 3.033
R73640 out.n10194 out.n10193 3.033
R73641 out.n10207 out.n10206 3.033
R73642 out.n10251 out.n10250 3.033
R73643 out.n12844 out.n12843 3.033
R73644 out.n13000 out.n12999 3.033
R73645 out.n12862 out.n12861 3.033
R73646 out.n13217 out.n13216 3.033
R73647 out.n12661 out.n12660 3.033
R73648 out.n12767 out.n12766 3.033
R73649 out.n12384 out.n12383 3.033
R73650 out.n12135 out.n12134 3.033
R73651 out.n11995 out.n11994 3.033
R73652 out.n12352 out.n12351 3.033
R73653 out.n13494 out.n13493 3.033
R73654 out.n13601 out.n13600 3.033
R73655 out.n11202 out.n11201 3.033
R73656 out.n11178 out.n11177 3.033
R73657 out.n11160 out.n11159 3.033
R73658 out.n11521 out.n11520 3.033
R73659 out.n10772 out.n10771 3.033
R73660 out.n10882 out.n10881 3.033
R73661 out.n10737 out.n10736 3.033
R73662 out.n11094 out.n11093 3.033
R73663 out.n11965 out.n11964 3.033
R73664 out.n11715 out.n11714 3.033
R73665 out.n11577 out.n11576 3.033
R73666 out.n11932 out.n11931 3.033
R73667 out.n13949 out.n13948 3.033
R73668 out.n14056 out.n14055 3.033
R73669 out.n10698 out.n10697 3.033
R73670 out.n10448 out.n10447 3.033
R73671 out.n10310 out.n10309 3.033
R73672 out.n10665 out.n10664 3.033
R73673 out.n14345 out.n14344 3.033
R73674 out.n14479 out.n14478 3.033
R73675 out.n1017 out.n1016 3.033
R73676 out.n5033 out.n5032 3.033
R73677 out.n5153 out.n5152 3.033
R73678 out.n5837 out.n5836 3.033
R73679 out.n5378 out.n5377 3.033
R73680 out.n5279 out.n5278 3.033
R73681 out.n1230 out.n1229 3.033
R73682 out.n6409 out.n6408 3.033
R73683 out.n6095 out.n6094 3.033
R73684 out.n5997 out.n5996 3.033
R73685 out.n6971 out.n6970 3.033
R73686 out.n7146 out.n7145 3.033
R73687 out.n7792 out.n7791 3.033
R73688 out.n6190 out.n6189 3.033
R73689 out.n2401 out.n2400 3.032
R73690 out.n1351 out.n1350 3.024
R73691 out.n2085 out.n2084 3.024
R73692 out.n2195 out.n2194 3.024
R73693 out.n10086 out.n10085 3.011
R73694 out.n12843 out.n12842 3.011
R73695 out.n13175 out.n13174 3.011
R73696 out.n13232 out.n13231 3.011
R73697 out.n12643 out.n12642 3.011
R73698 out.n12687 out.n12686 3.011
R73699 out.n12383 out.n12382 3.011
R73700 out.n12310 out.n12309 3.011
R73701 out.n11980 out.n11979 3.011
R73702 out.n13476 out.n13475 3.011
R73703 out.n13521 out.n13520 3.011
R73704 out.n11201 out.n11200 3.011
R73705 out.n11479 out.n11478 3.011
R73706 out.n11140 out.n11139 3.011
R73707 out.n10771 out.n10770 3.011
R73708 out.n11052 out.n11051 3.011
R73709 out.n10717 out.n10716 3.011
R73710 out.n11964 out.n11963 3.011
R73711 out.n11890 out.n11889 3.011
R73712 out.n11563 out.n11562 3.011
R73713 out.n13931 out.n13930 3.011
R73714 out.n13976 out.n13975 3.011
R73715 out.n10697 out.n10696 3.011
R73716 out.n10623 out.n10622 3.011
R73717 out.n10296 out.n10295 3.011
R73718 out.n14310 out.n14309 3.011
R73719 out.n14264 out.n14263 3.011
R73720 out.n4997 out.n4996 3.011
R73721 out.n2731 out.n2730 3.011
R73722 out.n5749 out.n5748 3.011
R73723 out.n5682 out.n5681 3.011
R73724 out.n1342 out.n1341 3.011
R73725 out.n5451 out.n5450 3.011
R73726 out.n5428 out.n5427 3.011
R73727 out.n1497 out.n1496 3.011
R73728 out.n5289 out.n5288 3.011
R73729 out.n2078 out.n2077 3.011
R73730 out.n6496 out.n6495 3.011
R73731 out.n6614 out.n6613 3.011
R73732 out.n2120 out.n2119 3.011
R73733 out.n1860 out.n1859 3.011
R73734 out.n6326 out.n6325 3.011
R73735 out.n6259 out.n6258 3.011
R73736 out.n5996 out.n5995 3.011
R73737 out.n1635 out.n1634 3.011
R73738 out.n6883 out.n6882 3.011
R73739 out.n6816 out.n6815 3.011
R73740 out.n2186 out.n2185 3.011
R73741 out.n7309 out.n7308 3.011
R73742 out.n7289 out.n7288 3.011
R73743 out.n2344 out.n2343 3.011
R73744 out.n2426 out.n2424 3.011
R73745 out.n2622 out.n2621 3.011
R73746 out.n7709 out.n7708 3.011
R73747 out.n7663 out.n7662 3.011
R73748 out.n10145 out.n10083 2.953
R73749 out.n10171 out.n10070 2.953
R73750 out.n10170 out.n10073 2.953
R73751 out.n10168 out.n10074 2.953
R73752 out.n10166 out.n10078 2.953
R73753 out.n10214 out.n10211 2.953
R73754 out.n10228 out.n10061 2.953
R73755 out.n10248 out.n10055 2.953
R73756 out.n10230 out.n10056 2.953
R73757 out.n12968 out.n12892 2.953
R73758 out.n13080 out.n12875 2.953
R73759 out.n13081 out.n12874 2.953
R73760 out.n13081 out.n12871 2.953
R73761 out.n13215 out.n12859 2.953
R73762 out.n13215 out.n12857 2.953
R73763 out.n12541 out.n12455 2.953
R73764 out.n12662 out.n12437 2.953
R73765 out.n12662 out.n12440 2.953
R73766 out.n12792 out.n12421 2.953
R73767 out.n12792 out.n12419 2.953
R73768 out.n12793 out.n12416 2.953
R73769 out.n12103 out.n12025 2.953
R73770 out.n12215 out.n12008 2.953
R73771 out.n12216 out.n12007 2.953
R73772 out.n12216 out.n12004 2.953
R73773 out.n12350 out.n11992 2.953
R73774 out.n12350 out.n11989 2.953
R73775 out.n13374 out.n13299 2.953
R73776 out.n13495 out.n13281 2.953
R73777 out.n13495 out.n13284 2.953
R73778 out.n13626 out.n13266 2.953
R73779 out.n13626 out.n13263 2.953
R73780 out.n13627 out.n13261 2.953
R73781 out.n11280 out.n11193 2.953
R73782 out.n11389 out.n11173 2.953
R73783 out.n11390 out.n11172 2.953
R73784 out.n11390 out.n11169 2.953
R73785 out.n11519 out.n11152 2.953
R73786 out.n11519 out.n11149 2.953
R73787 out.n10850 out.n10767 2.953
R73788 out.n10962 out.n10750 2.953
R73789 out.n10963 out.n10749 2.953
R73790 out.n10963 out.n10746 2.953
R73791 out.n11092 out.n10729 2.953
R73792 out.n11092 out.n10726 2.953
R73793 out.n11683 out.n11607 2.953
R73794 out.n11795 out.n11590 2.953
R73795 out.n11796 out.n11589 2.953
R73796 out.n11796 out.n11587 2.953
R73797 out.n11930 out.n11574 2.953
R73798 out.n11930 out.n11572 2.953
R73799 out.n13829 out.n13754 2.953
R73800 out.n13950 out.n13737 2.953
R73801 out.n13950 out.n13739 2.953
R73802 out.n14081 out.n13721 2.953
R73803 out.n14081 out.n13719 2.953
R73804 out.n14082 out.n13716 2.953
R73805 out.n10416 out.n10340 2.953
R73806 out.n10528 out.n10323 2.953
R73807 out.n10529 out.n10322 2.953
R73808 out.n10529 out.n10320 2.953
R73809 out.n10663 out.n10307 2.953
R73810 out.n10663 out.n10305 2.953
R73811 out.n14424 out.n14368 2.953
R73812 out.n14425 out.n14367 2.953
R73813 out.n14425 out.n14365 2.953
R73814 out.n14477 out.n14275 2.953
R73815 out.n14477 out.n14273 2.953
R73816 out.n14530 out.n14190 2.953
R73817 out.n1063 out.n979 2.953
R73818 out.n5098 out.n5057 2.953
R73819 out.n5099 out.n5056 2.953
R73820 out.n5099 out.n5054 2.953
R73821 out.n5151 out.n4961 2.953
R73822 out.n5151 out.n4958 2.953
R73823 out.n5838 out.n5641 2.953
R73824 out.n5588 out.n5399 2.953
R73825 out.n5371 out.n5370 2.953
R73826 out.n5371 out.n5367 2.953
R73827 out.n5358 out.n5181 2.953
R73828 out.n5248 out.n5194 2.953
R73829 out.n5249 out.n5192 2.953
R73830 out.n6742 out.n6458 2.953
R73831 out.n6410 out.n6213 2.953
R73832 out.n6178 out.n6177 2.953
R73833 out.n6178 out.n6174 2.953
R73834 out.n6172 out.n5879 2.953
R73835 out.n6066 out.n5904 2.953
R73836 out.n6972 out.n6775 2.953
R73837 out.n7446 out.n7260 2.953
R73838 out.n7217 out.n7027 2.953
R73839 out.n7218 out.n7025 2.953
R73840 out.n7793 out.n7486 2.953
R73841 out.n2779 out.n2778 2.871
R73842 out.n1903 out.n1902 2.871
R73843 out.n1683 out.n1682 2.871
R73844 out.n2643 out.n2642 2.871
R73845 out.n10093 out.n10092 2.826
R73846 out.n1203 out.n1202 2.82
R73847 out.n7119 out.n7118 2.82
R73848 out.n10224 out.n10223 2.819
R73849 out.n5482 out.n5481 2.819
R73850 out.n6646 out.n6645 2.819
R73851 out.n7340 out.n7339 2.819
R73852 out.n5761 out.n5760 2.722
R73853 out.n6338 out.n6337 2.722
R73854 out.n6895 out.n6894 2.722
R73855 out.n7721 out.n7720 2.722
R73856 out.n2741 out.n2740 2.67
R73857 out.n5725 out.n5723 2.67
R73858 out.n5484 out.n5482 2.67
R73859 out.n1436 out.n1435 2.67
R73860 out.n6648 out.n6646 2.67
R73861 out.n6507 out.n6506 2.67
R73862 out.n1870 out.n1869 2.67
R73863 out.n6302 out.n6300 2.67
R73864 out.n1645 out.n1644 2.67
R73865 out.n6859 out.n6857 2.67
R73866 out.n7342 out.n7340 2.67
R73867 out.n2280 out.n2279 2.67
R73868 out.n7515 out.n7513 2.67
R73869 out.n2858 out.n2856 2.641
R73870 out.n1982 out.n1980 2.641
R73871 out.n1762 out.n1760 2.641
R73872 out.n7619 out.n7617 2.641
R73873 out.n1145 out.n1144 2.639
R73874 out.n2492 out.n2491 2.639
R73875 out.n10155 out.n10154 2.635
R73876 out.n10268 out.n10267 2.635
R73877 out.n12939 out.n12938 2.635
R73878 out.n12951 out.n12950 2.635
R73879 out.n12074 out.n12073 2.635
R73880 out.n12086 out.n12085 2.635
R73881 out.n11251 out.n11250 2.635
R73882 out.n11263 out.n11262 2.635
R73883 out.n10821 out.n10820 2.635
R73884 out.n10833 out.n10832 2.635
R73885 out.n11654 out.n11653 2.635
R73886 out.n11666 out.n11665 2.635
R73887 out.n10387 out.n10386 2.635
R73888 out.n10399 out.n10398 2.635
R73889 out.n969 out.n968 2.635
R73890 out.n975 out.n974 2.635
R73891 out.n2834 out.n2833 2.635
R73892 out.n2826 out.n2825 2.635
R73893 out.n5411 out.n5410 2.635
R73894 out.n1418 out.n1417 2.635
R73895 out.n1373 out.n1371 2.635
R73896 out.n1362 out.n1361 2.635
R73897 out.n5229 out.n5228 2.635
R73898 out.n1288 out.n1287 2.635
R73899 out.n6480 out.n6479 2.635
R73900 out.n6522 out.n6521 2.635
R73901 out.n2135 out.n2133 2.635
R73902 out.n2096 out.n2095 2.635
R73903 out.n1958 out.n1957 2.635
R73904 out.n1950 out.n1949 2.635
R73905 out.n6048 out.n6047 2.635
R73906 out.n6036 out.n6035 2.635
R73907 out.n5933 out.n5932 2.635
R73908 out.n1567 out.n1566 2.635
R73909 out.n1738 out.n1737 2.635
R73910 out.n1730 out.n1729 2.635
R73911 out.n7272 out.n7271 2.635
R73912 out.n2262 out.n2261 2.635
R73913 out.n2217 out.n2215 2.635
R73914 out.n2206 out.n2205 2.635
R73915 out.n2389 out.n2388 2.635
R73916 out.n7196 out.n7195 2.635
R73917 out.n7086 out.n7085 2.635
R73918 out.n2474 out.n2473 2.635
R73919 out.n7566 out.n7565 2.635
R73920 out.n7573 out.n7572 2.635
R73921 out.n1438 out.n1437 2.605
R73922 out.n6509 out.n6508 2.605
R73923 out.n2282 out.n2281 2.605
R73924 out.n1557 out.n1556 2.495
R73925 out.n10127 out.n10124 2.442
R73926 out.n5980 out.n5979 2.442
R73927 out.n2841 out.n2840 2.44
R73928 out.n1965 out.n1964 2.44
R73929 out.n1745 out.n1744 2.44
R73930 out.n7553 out.n7552 2.44
R73931 out.n10174 out.n10173 2.28
R73932 out.n9434 out.n9429 2.268
R73933 out.n10127 out.n10126 2.258
R73934 out.n10064 out.n10063 2.258
R73935 out.n10219 out.n10218 2.258
R73936 out.n10281 out.n10280 2.258
R73937 out.n13009 out.n13008 2.258
R73938 out.n13065 out.n13064 2.258
R73939 out.n12463 out.n12462 2.258
R73940 out.n12524 out.n12523 2.258
R73941 out.n12523 out.n12522 2.258
R73942 out.n12633 out.n12632 2.258
R73943 out.n12406 out.n12405 2.258
R73944 out.n12144 out.n12143 2.258
R73945 out.n12200 out.n12199 2.258
R73946 out.n13659 out.n13658 2.258
R73947 out.n13357 out.n13356 2.258
R73948 out.n13356 out.n13355 2.258
R73949 out.n13466 out.n13465 2.258
R73950 out.n13251 out.n13250 2.258
R73951 out.n11318 out.n11317 2.258
R73952 out.n11374 out.n11373 2.258
R73953 out.n10891 out.n10890 2.258
R73954 out.n10947 out.n10946 2.258
R73955 out.n11724 out.n11723 2.258
R73956 out.n11780 out.n11779 2.258
R73957 out.n13692 out.n13691 2.258
R73958 out.n13812 out.n13811 2.258
R73959 out.n13811 out.n13810 2.258
R73960 out.n13921 out.n13920 2.258
R73961 out.n13706 out.n13705 2.258
R73962 out.n10457 out.n10456 2.258
R73963 out.n10513 out.n10512 2.258
R73964 out.n14163 out.n14162 2.258
R73965 out.n14377 out.n14376 2.258
R73966 out.n14256 out.n14255 2.258
R73967 out.n14183 out.n14182 2.258
R73968 out.n14184 out.n14183 2.258
R73969 out.n1024 out.n1023 2.258
R73970 out.n5066 out.n5065 2.258
R73971 out.n5812 out.n5811 2.258
R73972 out.n5690 out.n5689 2.258
R73973 out.n5566 out.n5565 2.258
R73974 out.n5565 out.n5564 2.258
R73975 out.n5505 out.n5504 2.258
R73976 out.n1402 out.n1401 2.258
R73977 out.n1205 out.n1204 2.258
R73978 out.n6720 out.n6719 2.258
R73979 out.n6719 out.n6718 2.258
R73980 out.n6669 out.n6668 2.258
R73981 out.n6537 out.n6536 2.258
R73982 out.n6384 out.n6383 2.258
R73983 out.n6267 out.n6266 2.258
R73984 out.n6157 out.n6156 2.258
R73985 out.n6106 out.n6105 2.258
R73986 out.n5982 out.n5981 2.258
R73987 out.n1549 out.n1548 2.258
R73988 out.n6946 out.n6945 2.258
R73989 out.n6824 out.n6823 2.258
R73990 out.n7424 out.n7423 2.258
R73991 out.n7423 out.n7422 2.258
R73992 out.n7363 out.n7362 2.258
R73993 out.n2246 out.n2245 2.258
R73994 out.n7121 out.n7120 2.258
R73995 out.n2418 out.n2417 2.258
R73996 out.n7767 out.n7766 2.258
R73997 out.n7671 out.n7670 2.258
R73998 out.n6192 out.n6191 2.25
R73999 out.n9442 out.n9427 2.249
R74000 out.n13642 out.n13641 2.249
R74001 out.n11539 out.n11538 2.249
R74002 out.n11112 out.n11111 2.249
R74003 out.n14097 out.n14096 2.249
R74004 out.n14563 out.n14562 2.249
R74005 out.n13244 out.n13243 2.249
R74006 out.n12823 out.n12822 2.248
R74007 out.n13670 out.n13669 2.248
R74008 out.n13703 out.n13702 2.248
R74009 out.n9440 out.n9439 2.247
R74010 out.n13245 out.n12853 2.247
R74011 out.n12393 out.n12392 2.247
R74012 out.n11555 out.n11554 2.247
R74013 out.n11132 out.n11131 2.247
R74014 out.n7815 out.n7814 2.247
R74015 out.n6758 out.n6757 2.247
R74016 out.n13245 out.n13238 2.245
R74017 out.n9440 out.n9438 2.245
R74018 out.n10131 out.n10093 2.102
R74019 out.n2832 out.n2831 2.066
R74020 out.n1956 out.n1955 2.066
R74021 out.n1736 out.n1735 2.066
R74022 out.n7564 out.n7563 2.066
R74023 out.n1141 out.n1140 2.064
R74024 out.n2484 out.n2483 2.064
R74025 out.n12821 out.n12820 2.025
R74026 out.n13668 out.n13667 2.025
R74027 out.n13701 out.n13700 2.025
R74028 out.n12852 out.n12851 2.014
R74029 out.n12391 out.n12390 2.014
R74030 out.n11553 out.n11552 2.014
R74031 out.n11130 out.n11129 2.014
R74032 out.n11973 out.n11972 2.014
R74033 out.n10706 out.n10705 2.014
R74034 out.n1205 out.n1203 1.925
R74035 out.n5982 out.n5980 1.925
R74036 out.n7121 out.n7119 1.925
R74037 out.n1215 out.n1213 1.91
R74038 out.n7133 out.n7131 1.91
R74039 out.n2743 out.n2742 1.89
R74040 out.n1872 out.n1871 1.89
R74041 out.n1647 out.n1646 1.89
R74042 out.n2700 out.n2699 1.89
R74043 out.n10152 out.n10151 1.882
R74044 out.n10184 out.n10183 1.882
R74045 out.n10224 out.n10222 1.882
R74046 out.n12959 out.n12958 1.882
R74047 out.n12881 out.n12880 1.882
R74048 out.n13066 out.n13065 1.882
R74049 out.n13165 out.n13164 1.882
R74050 out.n12444 out.n12443 1.882
R74051 out.n12699 out.n12698 1.882
R74052 out.n12407 out.n12406 1.882
R74053 out.n12094 out.n12093 1.882
R74054 out.n12014 out.n12013 1.882
R74055 out.n12201 out.n12200 1.882
R74056 out.n12300 out.n12299 1.882
R74057 out.n13288 out.n13287 1.882
R74058 out.n13533 out.n13532 1.882
R74059 out.n13252 out.n13251 1.882
R74060 out.n11271 out.n11270 1.882
R74061 out.n11182 out.n11181 1.882
R74062 out.n11375 out.n11374 1.882
R74063 out.n11469 out.n11468 1.882
R74064 out.n10841 out.n10840 1.882
R74065 out.n10756 out.n10755 1.882
R74066 out.n10948 out.n10947 1.882
R74067 out.n11042 out.n11041 1.882
R74068 out.n11674 out.n11673 1.882
R74069 out.n11596 out.n11595 1.882
R74070 out.n11781 out.n11780 1.882
R74071 out.n11880 out.n11879 1.882
R74072 out.n13743 out.n13742 1.882
R74073 out.n13988 out.n13987 1.882
R74074 out.n13707 out.n13706 1.882
R74075 out.n10407 out.n10406 1.882
R74076 out.n10329 out.n10328 1.882
R74077 out.n10514 out.n10513 1.882
R74078 out.n10613 out.n10612 1.882
R74079 out.n14378 out.n14377 1.882
R74080 out.n14320 out.n14319 1.882
R74081 out.n14202 out.n14200 1.882
R74082 out.n1073 out.n1072 1.882
R74083 out.n990 out.n989 1.882
R74084 out.n5067 out.n5066 1.882
R74085 out.n5007 out.n5006 1.882
R74086 out.n5725 out.n5724 1.882
R74087 out.n5652 out.n5651 1.882
R74088 out.n2842 out.n2841 1.882
R74089 out.n2844 out.n2843 1.882
R74090 out.n2820 out.n2819 1.882
R74091 out.n2761 out.n2760 1.882
R74092 out.n5484 out.n5483 1.882
R74093 out.n5417 out.n5416 1.882
R74094 out.n1452 out.n1451 1.882
R74095 out.n1411 out.n1410 1.882
R74096 out.n5346 out.n5345 1.882
R74097 out.n5238 out.n5237 1.882
R74098 out.n1197 out.n1196 1.882
R74099 out.n1280 out.n1279 1.882
R74100 out.n6648 out.n6647 1.882
R74101 out.n6486 out.n6485 1.882
R74102 out.n6500 out.n6499 1.882
R74103 out.n6528 out.n6527 1.882
R74104 out.n6302 out.n6301 1.882
R74105 out.n6229 out.n6228 1.882
R74106 out.n1966 out.n1965 1.882
R74107 out.n1968 out.n1967 1.882
R74108 out.n1944 out.n1943 1.882
R74109 out.n1890 out.n1889 1.882
R74110 out.n6158 out.n6157 1.882
R74111 out.n5898 out.n5897 1.882
R74112 out.n6056 out.n6055 1.882
R74113 out.n5969 out.n5968 1.882
R74114 out.n6859 out.n6858 1.882
R74115 out.n6786 out.n6785 1.882
R74116 out.n1746 out.n1745 1.882
R74117 out.n1748 out.n1747 1.882
R74118 out.n1724 out.n1723 1.882
R74119 out.n1665 out.n1664 1.882
R74120 out.n7342 out.n7341 1.882
R74121 out.n7278 out.n7277 1.882
R74122 out.n2296 out.n2295 1.882
R74123 out.n2255 out.n2254 1.882
R74124 out.n7205 out.n7204 1.882
R74125 out.n7050 out.n7049 1.882
R74126 out.n7094 out.n7093 1.882
R74127 out.n2467 out.n2466 1.882
R74128 out.n2458 out.n2457 1.882
R74129 out.n7515 out.n7514 1.882
R74130 out.n7522 out.n7521 1.882
R74131 out.n7554 out.n7553 1.882
R74132 out.n7556 out.n7555 1.882
R74133 out.n7600 out.n7599 1.882
R74134 out.n2636 out.n2635 1.882
R74135 out.n10273 out.n10272 1.844
R74136 out.n10274 out.n10273 1.823
R74137 out.n10213 out.n10212 1.799
R74138 out.n14180 out.n14179 1.691
R74139 out.n2478 out.n2477 1.69
R74140 out.n12905 out.n12904 1.614
R74141 out.n12481 out.n12480 1.614
R74142 out.n12040 out.n12039 1.614
R74143 out.n13314 out.n13313 1.614
R74144 out.n11217 out.n11216 1.614
R74145 out.n10787 out.n10786 1.614
R74146 out.n11620 out.n11619 1.614
R74147 out.n13769 out.n13768 1.614
R74148 out.n10353 out.n10352 1.614
R74149 out.n1096 out.n1095 1.614
R74150 out.n5776 out.n5775 1.614
R74151 out.n5523 out.n5522 1.614
R74152 out.n1242 out.n1241 1.614
R74153 out.n6467 out.n6466 1.614
R74154 out.n6217 out.n6216 1.614
R74155 out.n5913 out.n5912 1.614
R74156 out.n6910 out.n6909 1.614
R74157 out.n7381 out.n7380 1.614
R74158 out.n7038 out.n7037 1.614
R74159 out.n7490 out.n7489 1.614
R74160 out.n10151 out.n10150 1.505
R74161 out.n10065 out.n10064 1.505
R74162 out.n10185 out.n10184 1.505
R74163 out.n10280 out.n10279 1.505
R74164 out.n10261 out.n10260 1.505
R74165 out.n12950 out.n12949 1.505
R74166 out.n12981 out.n12980 1.505
R74167 out.n13119 out.n13118 1.505
R74168 out.n13120 out.n13119 1.505
R74169 out.n13233 out.n13232 1.505
R74170 out.n12533 out.n12532 1.505
R74171 out.n12585 out.n12584 1.505
R74172 out.n12644 out.n12643 1.505
R74173 out.n12744 out.n12743 1.505
R74174 out.n12743 out.n12742 1.505
R74175 out.n12085 out.n12084 1.505
R74176 out.n12116 out.n12115 1.505
R74177 out.n12254 out.n12253 1.505
R74178 out.n12255 out.n12254 1.505
R74179 out.n11981 out.n11980 1.505
R74180 out.n13366 out.n13365 1.505
R74181 out.n13418 out.n13417 1.505
R74182 out.n13477 out.n13476 1.505
R74183 out.n13578 out.n13577 1.505
R74184 out.n13577 out.n13576 1.505
R74185 out.n11262 out.n11261 1.505
R74186 out.n11293 out.n11292 1.505
R74187 out.n11423 out.n11422 1.505
R74188 out.n11424 out.n11423 1.505
R74189 out.n11141 out.n11140 1.505
R74190 out.n10832 out.n10831 1.505
R74191 out.n10863 out.n10862 1.505
R74192 out.n10996 out.n10995 1.505
R74193 out.n10997 out.n10996 1.505
R74194 out.n10718 out.n10717 1.505
R74195 out.n11665 out.n11664 1.505
R74196 out.n11696 out.n11695 1.505
R74197 out.n11834 out.n11833 1.505
R74198 out.n11835 out.n11834 1.505
R74199 out.n11564 out.n11563 1.505
R74200 out.n13821 out.n13820 1.505
R74201 out.n13873 out.n13872 1.505
R74202 out.n13932 out.n13931 1.505
R74203 out.n14033 out.n14032 1.505
R74204 out.n14032 out.n14031 1.505
R74205 out.n10398 out.n10397 1.505
R74206 out.n10429 out.n10428 1.505
R74207 out.n10567 out.n10566 1.505
R74208 out.n10568 out.n10567 1.505
R74209 out.n10297 out.n10296 1.505
R74210 out.n14324 out.n14323 1.505
R74211 out.n14325 out.n14324 1.505
R74212 out.n14265 out.n14264 1.505
R74213 out.n14239 out.n14238 1.505
R74214 out.n14541 out.n14540 1.505
R74215 out.n974 out.n973 1.505
R74216 out.n999 out.n998 1.505
R74217 out.n5011 out.n5010 1.505
R74218 out.n5012 out.n5011 1.505
R74219 out.n5821 out.n5820 1.505
R74220 out.n5811 out.n5810 1.505
R74221 out.n5698 out.n5697 1.505
R74222 out.n2811 out.n2810 1.505
R74223 out.n5577 out.n5576 1.505
R74224 out.n5450 out.n5449 1.505
R74225 out.n5345 out.n5344 1.505
R74226 out.n5259 out.n5258 1.505
R74227 out.n1213 out.n1212 1.505
R74228 out.n1215 out.n1214 1.505
R74229 out.n1162 out.n1161 1.505
R74230 out.n6731 out.n6730 1.505
R74231 out.n6495 out.n6494 1.505
R74232 out.n6393 out.n6392 1.505
R74233 out.n6383 out.n6382 1.505
R74234 out.n6275 out.n6274 1.505
R74235 out.n1935 out.n1934 1.505
R74236 out.n6084 out.n6083 1.505
R74237 out.n6047 out.n6046 1.505
R74238 out.n5927 out.n5926 1.505
R74239 out.n1566 out.n1565 1.505
R74240 out.n6955 out.n6954 1.505
R74241 out.n6945 out.n6944 1.505
R74242 out.n6832 out.n6831 1.505
R74243 out.n1715 out.n1714 1.505
R74244 out.n7435 out.n7434 1.505
R74245 out.n7308 out.n7307 1.505
R74246 out.n2392 out.n2391 1.505
R74247 out.n7228 out.n7227 1.505
R74248 out.n7131 out.n7130 1.505
R74249 out.n7133 out.n7132 1.505
R74250 out.n2507 out.n2506 1.505
R74251 out.n7776 out.n7775 1.505
R74252 out.n7766 out.n7765 1.505
R74253 out.n7679 out.n7678 1.505
R74254 out.n7580 out.n7579 1.505
R74255 out.n10286 out.n10283 1.498
R74256 out.n11975 out.n11974 1.498
R74257 out.n10708 out.n10707 1.498
R74258 out.n9440 out.n9431 1.49
R74259 out.n9441 out.n9440 1.489
R74260 out.n9440 out.n9435 1.488
R74261 out.n5461 out.n5460 1.428
R74262 out.n6626 out.n6625 1.428
R74263 out.n7319 out.n7318 1.428
R74264 out.n5461 out.n5458 1.426
R74265 out.n6626 out.n6623 1.426
R74266 out.n7319 out.n7316 1.426
R74267 out.n5955 out.n5952 1.411
R74268 out.n2804 out.n2800 1.397
R74269 out.n1928 out.n1924 1.397
R74270 out.n1708 out.n1704 1.397
R74271 out.n7591 out.n7587 1.397
R74272 out.n2449 out.n2445 1.385
R74273 out.n5873 out.n5872 1.362
R74274 out.n7808 out.n7807 1.351
R74275 out.n6751 out.n6750 1.332
R74276 out.n1354 out.n1353 1.186
R74277 out.n2088 out.n2087 1.186
R74278 out.n2198 out.n2197 1.186
R74279 out.n2834 out.n2832 1.179
R74280 out.n1958 out.n1956 1.179
R74281 out.n1738 out.n1736 1.179
R74282 out.n7566 out.n7564 1.179
R74283 out.n10126 out.n10125 1.129
R74284 out.n10163 out.n10162 1.129
R74285 out.n10157 out.n10155 1.129
R74286 out.n10220 out.n10219 1.129
R74287 out.n10244 out.n10243 1.129
R74288 out.n10237 out.n10236 1.129
R74289 out.n12966 out.n12965 1.129
R74290 out.n12887 out.n12886 1.129
R74291 out.n13077 out.n13076 1.129
R74292 out.n12867 out.n12866 1.129
R74293 out.n13176 out.n13175 1.129
R74294 out.n13210 out.n13208 1.129
R74295 out.n12450 out.n12449 1.129
R74296 out.n12555 out.n12554 1.129
R74297 out.n12553 out.n12552 1.129
R74298 out.n12586 out.n12585 1.129
R74299 out.n12433 out.n12432 1.129
R74300 out.n12688 out.n12687 1.129
R74301 out.n12787 out.n12785 1.129
R74302 out.n12796 out.n12795 1.129
R74303 out.n12101 out.n12100 1.129
R74304 out.n12020 out.n12019 1.129
R74305 out.n12212 out.n12211 1.129
R74306 out.n12000 out.n11999 1.129
R74307 out.n12311 out.n12310 1.129
R74308 out.n12345 out.n12343 1.129
R74309 out.n13294 out.n13293 1.129
R74310 out.n13388 out.n13387 1.129
R74311 out.n13386 out.n13385 1.129
R74312 out.n13419 out.n13418 1.129
R74313 out.n13277 out.n13276 1.129
R74314 out.n13522 out.n13521 1.129
R74315 out.n13621 out.n13619 1.129
R74316 out.n13630 out.n13629 1.129
R74317 out.n11278 out.n11277 1.129
R74318 out.n11188 out.n11187 1.129
R74319 out.n11386 out.n11385 1.129
R74320 out.n11165 out.n11164 1.129
R74321 out.n11480 out.n11479 1.129
R74322 out.n11514 out.n11512 1.129
R74323 out.n10848 out.n10847 1.129
R74324 out.n10762 out.n10761 1.129
R74325 out.n10959 out.n10958 1.129
R74326 out.n10742 out.n10741 1.129
R74327 out.n11053 out.n11052 1.129
R74328 out.n11087 out.n11085 1.129
R74329 out.n11681 out.n11680 1.129
R74330 out.n11602 out.n11601 1.129
R74331 out.n11792 out.n11791 1.129
R74332 out.n11582 out.n11581 1.129
R74333 out.n11891 out.n11890 1.129
R74334 out.n11925 out.n11923 1.129
R74335 out.n13749 out.n13748 1.129
R74336 out.n13843 out.n13842 1.129
R74337 out.n13841 out.n13840 1.129
R74338 out.n13874 out.n13873 1.129
R74339 out.n13732 out.n13731 1.129
R74340 out.n13977 out.n13976 1.129
R74341 out.n14076 out.n14074 1.129
R74342 out.n14085 out.n14084 1.129
R74343 out.n10414 out.n10413 1.129
R74344 out.n10335 out.n10334 1.129
R74345 out.n10525 out.n10524 1.129
R74346 out.n10315 out.n10314 1.129
R74347 out.n10624 out.n10623 1.129
R74348 out.n10658 out.n10656 1.129
R74349 out.n14421 out.n14420 1.129
R74350 out.n14359 out.n14358 1.129
R74351 out.n14311 out.n14310 1.129
R74352 out.n14280 out.n14278 1.129
R74353 out.n14240 out.n14239 1.129
R74354 out.n14212 out.n14211 1.129
R74355 out.n14213 out.n14209 1.129
R74356 out.n14195 out.n14193 1.129
R74357 out.n1065 out.n1064 1.129
R74358 out.n983 out.n982 1.129
R74359 out.n5095 out.n5094 1.129
R74360 out.n5048 out.n5047 1.129
R74361 out.n4998 out.n4997 1.129
R74362 out.n4966 out.n4964 1.129
R74363 out.n2734 out.n2733 1.129
R74364 out.n5848 out.n5847 1.129
R74365 out.n5637 out.n5636 1.129
R74366 out.n5735 out.n5734 1.129
R74367 out.n5737 out.n5736 1.129
R74368 out.n5712 out.n5711 1.129
R74369 out.n2868 out.n2867 1.129
R74370 out.n2851 out.n2850 1.129
R74371 out.n5599 out.n5598 1.129
R74372 out.n5394 out.n5393 1.129
R74373 out.n5405 out.n5404 1.129
R74374 out.n5468 out.n5467 1.129
R74375 out.n5355 out.n5354 1.129
R74376 out.n5188 out.n5187 1.129
R74377 out.n5245 out.n5244 1.129
R74378 out.n1190 out.n1189 1.129
R74379 out.n1273 out.n1272 1.129
R74380 out.n6755 out.n6754 1.129
R74381 out.n6453 out.n6452 1.129
R74382 out.n6474 out.n6473 1.129
R74383 out.n6632 out.n6631 1.129
R74384 out.n1863 out.n1862 1.129
R74385 out.n6420 out.n6419 1.129
R74386 out.n6209 out.n6208 1.129
R74387 out.n6312 out.n6311 1.129
R74388 out.n6314 out.n6313 1.129
R74389 out.n6289 out.n6288 1.129
R74390 out.n1992 out.n1991 1.129
R74391 out.n1975 out.n1974 1.129
R74392 out.n5876 out.n5875 1.129
R74393 out.n6169 out.n6168 1.129
R74394 out.n6071 out.n6070 1.129
R74395 out.n6064 out.n6063 1.129
R74396 out.n5961 out.n5960 1.129
R74397 out.n1638 out.n1637 1.129
R74398 out.n6982 out.n6981 1.129
R74399 out.n6771 out.n6770 1.129
R74400 out.n6869 out.n6868 1.129
R74401 out.n6871 out.n6870 1.129
R74402 out.n6846 out.n6845 1.129
R74403 out.n1772 out.n1771 1.129
R74404 out.n1755 out.n1754 1.129
R74405 out.n7457 out.n7456 1.129
R74406 out.n7255 out.n7254 1.129
R74407 out.n7266 out.n7265 1.129
R74408 out.n7326 out.n7325 1.129
R74409 out.n7021 out.n7020 1.129
R74410 out.n7214 out.n7213 1.129
R74411 out.n7108 out.n7107 1.129
R74412 out.n7101 out.n7100 1.129
R74413 out.n2624 out.n2623 1.129
R74414 out.n7482 out.n7481 1.129
R74415 out.n7503 out.n7502 1.129
R74416 out.n7505 out.n7504 1.129
R74417 out.n7692 out.n7691 1.129
R74418 out.n7538 out.n7537 1.129
R74419 out.n7547 out.n7546 1.129
R74420 out.n9461 out.n9460 1.11
R74421 out.n2749 out.n2748 1.066
R74422 out.n1878 out.n1877 1.066
R74423 out.n1653 out.n1652 1.066
R74424 out.n2694 out.n2693 1.066
R74425 out.n1126 out.n1125 1.066
R74426 out.n10178 out.n10174 1.002
R74427 out.n10177 out.n10175 0.944
R74428 out.n12457 out.n12456 0.886
R74429 out.n13650 out.n13649 0.886
R74430 out.n13683 out.n13682 0.886
R74431 out.n5494 out.n5493 0.886
R74432 out.n6658 out.n6657 0.886
R74433 out.n7352 out.n7351 0.886
R74434 out.n1151 out.n1149 0.874
R74435 out.n2497 out.n2495 0.874
R74436 out.n2590 out.n2589 0.841
R74437 out.n2938 out.n2937 0.84
R74438 out.n2067 out.n2066 0.84
R74439 out.n1842 out.n1841 0.84
R74440 out.n1331 out.n1330 0.835
R74441 out.n12851 out.n12850 0.831
R74442 out.n12390 out.n12389 0.831
R74443 out.n11552 out.n11551 0.831
R74444 out.n11129 out.n11128 0.831
R74445 out.n11972 out.n11971 0.831
R74446 out.n10705 out.n10704 0.831
R74447 out.n12820 out.n12819 0.825
R74448 out.n13667 out.n13666 0.825
R74449 out.n13700 out.n13699 0.825
R74450 out.n14178 out.n14177 0.818
R74451 out.n1527 out.n1526 0.804
R74452 out.n2374 out.n2373 0.804
R74453 out.n2844 out.n2842 0.788
R74454 out.n1968 out.n1966 0.788
R74455 out.n1748 out.n1746 0.788
R74456 out.n7556 out.n7554 0.788
R74457 out.n10100 out.n10099 0.76
R74458 out.n2406 out.n2405 0.755
R74459 out.n10112 out.n10111 0.752
R74460 out.n10087 out.n10086 0.752
R74461 out.n10138 out.n10137 0.752
R74462 out.n10203 out.n10202 0.752
R74463 out.n10269 out.n10268 0.752
R74464 out.n12837 out.n12836 0.752
R74465 out.n12938 out.n12937 0.752
R74466 out.n12989 out.n12988 0.752
R74467 out.n13010 out.n13009 0.752
R74468 out.n13089 out.n13088 0.752
R74469 out.n13109 out.n13108 0.752
R74470 out.n13164 out.n13163 0.752
R74471 out.n13222 out.n13221 0.752
R74472 out.n12539 out.n12538 0.752
R74473 out.n12809 out.n12808 0.752
R74474 out.n12632 out.n12631 0.752
R74475 out.n12655 out.n12654 0.752
R74476 out.n12698 out.n12697 0.752
R74477 out.n12755 out.n12754 0.752
R74478 out.n12778 out.n12776 0.752
R74479 out.n12378 out.n12377 0.752
R74480 out.n12073 out.n12072 0.752
R74481 out.n12124 out.n12123 0.752
R74482 out.n12145 out.n12144 0.752
R74483 out.n12224 out.n12223 0.752
R74484 out.n12244 out.n12243 0.752
R74485 out.n12299 out.n12298 0.752
R74486 out.n12357 out.n12356 0.752
R74487 out.n13372 out.n13371 0.752
R74488 out.n13645 out.n13644 0.752
R74489 out.n13465 out.n13464 0.752
R74490 out.n13488 out.n13487 0.752
R74491 out.n13532 out.n13531 0.752
R74492 out.n13589 out.n13588 0.752
R74493 out.n13612 out.n13610 0.752
R74494 out.n11546 out.n11545 0.752
R74495 out.n11250 out.n11249 0.752
R74496 out.n11301 out.n11300 0.752
R74497 out.n11319 out.n11318 0.752
R74498 out.n11398 out.n11397 0.752
R74499 out.n11156 out.n11155 0.752
R74500 out.n11468 out.n11467 0.752
R74501 out.n11526 out.n11525 0.752
R74502 out.n11122 out.n11121 0.752
R74503 out.n10820 out.n10819 0.752
R74504 out.n10871 out.n10870 0.752
R74505 out.n10892 out.n10891 0.752
R74506 out.n10971 out.n10970 0.752
R74507 out.n10733 out.n10732 0.752
R74508 out.n11041 out.n11040 0.752
R74509 out.n11099 out.n11098 0.752
R74510 out.n11958 out.n11957 0.752
R74511 out.n11653 out.n11652 0.752
R74512 out.n11704 out.n11703 0.752
R74513 out.n11725 out.n11724 0.752
R74514 out.n11804 out.n11803 0.752
R74515 out.n11824 out.n11823 0.752
R74516 out.n11879 out.n11878 0.752
R74517 out.n11937 out.n11936 0.752
R74518 out.n13827 out.n13826 0.752
R74519 out.n13678 out.n13677 0.752
R74520 out.n13920 out.n13919 0.752
R74521 out.n13943 out.n13942 0.752
R74522 out.n13987 out.n13986 0.752
R74523 out.n14044 out.n14043 0.752
R74524 out.n14067 out.n14065 0.752
R74525 out.n10691 out.n10690 0.752
R74526 out.n10386 out.n10385 0.752
R74527 out.n10437 out.n10436 0.752
R74528 out.n10458 out.n10457 0.752
R74529 out.n10537 out.n10536 0.752
R74530 out.n10557 out.n10556 0.752
R74531 out.n10612 out.n10611 0.752
R74532 out.n10670 out.n10669 0.752
R74533 out.n14164 out.n14163 0.752
R74534 out.n14348 out.n14347 0.752
R74535 out.n14334 out.n14333 0.752
R74536 out.n14319 out.n14318 0.752
R74537 out.n14484 out.n14483 0.752
R74538 out.n14255 out.n14254 0.752
R74539 out.n14532 out.n14531 0.752
R74540 out.n14559 out.n14558 0.752
R74541 out.n941 out.n940 0.752
R74542 out.n968 out.n967 0.752
R74543 out.n1008 out.n1007 0.752
R74544 out.n1025 out.n1024 0.752
R74545 out.n5037 out.n5036 0.752
R74546 out.n5021 out.n5020 0.752
R74547 out.n5006 out.n5005 0.752
R74548 out.n5158 out.n5157 0.752
R74549 out.n5830 out.n5829 0.752
R74550 out.n5705 out.n5704 0.752
R74551 out.n5681 out.n5680 0.752
R74552 out.n5586 out.n5585 0.752
R74553 out.n5427 out.n5426 0.752
R74554 out.n5383 out.n5382 0.752
R74555 out.n5176 out.n5175 0.752
R74556 out.n5290 out.n5289 0.752
R74557 out.n5268 out.n5267 0.752
R74558 out.n5228 out.n5227 0.752
R74559 out.n1222 out.n1221 0.752
R74560 out.n6740 out.n6739 0.752
R74561 out.n6613 out.n6612 0.752
R74562 out.n6402 out.n6401 0.752
R74563 out.n6282 out.n6281 0.752
R74564 out.n6258 out.n6257 0.752
R74565 out.n6107 out.n6106 0.752
R74566 out.n5892 out.n5891 0.752
R74567 out.n6035 out.n6034 0.752
R74568 out.n5919 out.n5918 0.752
R74569 out.n5945 out.n5944 0.752
R74570 out.n6964 out.n6963 0.752
R74571 out.n6839 out.n6838 0.752
R74572 out.n6815 out.n6814 0.752
R74573 out.n7444 out.n7443 0.752
R74574 out.n7288 out.n7287 0.752
R74575 out.n7239 out.n7238 0.752
R74576 out.n7195 out.n7194 0.752
R74577 out.n7044 out.n7043 0.752
R74578 out.n2452 out.n2451 0.752
R74579 out.n7785 out.n7784 0.752
R74580 out.n7686 out.n7685 0.752
R74581 out.n7662 out.n7661 0.752
R74582 out.n5595 out.n5594 0.671
R74583 out.n6752 out.n6751 0.671
R74584 out.n7453 out.n7452 0.671
R74585 out.n7235 out.n7234 0.662
R74586 out.n5855 out.n5854 0.652
R74587 out.n6427 out.n6426 0.652
R74588 out.n6989 out.n6988 0.652
R74589 out.n7809 out.n7808 0.652
R74590 out.n6191 out.n5873 0.646
R74591 out.n5173 out.n5171 0.613
R74592 out.n9652 out.t9 0.612
R74593 out.n9661 out.t15 0.612
R74594 out.n5643 out.n5642 0.586
R74595 out.n6220 out.n6219 0.586
R74596 out.n6777 out.n6776 0.586
R74597 out.n7493 out.n7492 0.586
R74598 out.n1398 out.n1397 0.579
R74599 out.n2117 out.n2116 0.579
R74600 out.n2242 out.n2241 0.579
R74601 out.n12834 out.n12833 0.575
R74602 out.n12375 out.n12374 0.575
R74603 out.n11195 out.n11194 0.575
R74604 out.n11119 out.n11118 0.575
R74605 out.n11955 out.n11954 0.575
R74606 out.n10688 out.n10687 0.575
R74607 out.n938 out.n937 0.575
R74608 out.n5916 out.n5915 0.575
R74609 out.n1444 out.n1442 0.575
R74610 out.n6564 out.n6562 0.575
R74611 out.n2288 out.n2286 0.575
R74612 out.n2449 out.n2448 0.572
R74613 out.n2804 out.n2803 0.568
R74614 out.n1928 out.n1927 0.568
R74615 out.n1708 out.n1707 0.568
R74616 out.n7591 out.n7590 0.568
R74617 out.n1398 out.n1395 0.566
R74618 out.n2117 out.n2114 0.566
R74619 out.n5955 out.n5954 0.566
R74620 out.n2242 out.n2239 0.566
R74621 out.n10273 out.t40 0.553
R74622 out.n10273 out.t52 0.553
R74623 out.n12851 out.t50 0.553
R74624 out.n12851 out.t42 0.553
R74625 out.n12820 out.t54 0.553
R74626 out.n12820 out.t28 0.553
R74627 out.n12390 out.t46 0.553
R74628 out.n12390 out.t39 0.553
R74629 out.n13667 out.t30 0.553
R74630 out.n13667 out.t49 0.553
R74631 out.n11552 out.t60 0.553
R74632 out.n11552 out.t34 0.553
R74633 out.n11129 out.t27 0.553
R74634 out.n11129 out.t45 0.553
R74635 out.n11972 out.t37 0.553
R74636 out.n11972 out.t56 0.553
R74637 out.n13700 out.t22 0.553
R74638 out.n13700 out.t64 0.553
R74639 out.n10705 out.t33 0.553
R74640 out.n10705 out.t25 0.553
R74641 out.n14178 out.t62 0.553
R74642 out.n14178 out.t58 0.553
R74643 out.n1124 out.t61 0.553
R74644 out.n1124 out.t57 0.553
R74645 out.n2937 out.t35 0.553
R74646 out.n2937 out.t55 0.553
R74647 out.n1526 out.t65 0.553
R74648 out.n1526 out.t63 0.553
R74649 out.n1330 out.t31 0.553
R74650 out.n1330 out.t23 0.553
R74651 out.n6750 out.t38 0.553
R74652 out.n6750 out.t51 0.553
R74653 out.n2066 out.t48 0.553
R74654 out.n2066 out.t41 0.553
R74655 out.n5872 out.t53 0.553
R74656 out.n5872 out.t26 0.553
R74657 out.n1841 out.t44 0.553
R74658 out.n1841 out.t36 0.553
R74659 out.n2373 out.t29 0.553
R74660 out.n2373 out.t47 0.553
R74661 out.n2589 out.t59 0.553
R74662 out.n2589 out.t32 0.553
R74663 out.n7807 out.t24 0.553
R74664 out.n7807 out.t43 0.553
R74665 out.n6184 out.n6183 0.552
R74666 out.n1438 out.n1436 0.533
R74667 out.n6509 out.n6507 0.533
R74668 out.n5924 out.n5922 0.533
R74669 out.n2282 out.n2280 0.533
R74670 out.n1528 out.n1527 0.516
R74671 out.n2166 out.n2165 0.516
R74672 out.n2375 out.n2374 0.516
R74673 out.n1609 out.n1608 0.509
R74674 out.n14179 out.n14178 0.504
R74675 out.n9660 out.n9659 0.501
R74676 out.n9659 out.n9658 0.501
R74677 out.n9658 out.n9657 0.501
R74678 out.n9657 out.n9656 0.501
R74679 out.n9656 out.n9655 0.501
R74680 out.n9655 out.n9654 0.501
R74681 out.n9654 out.n9653 0.501
R74682 out.n9653 out.n9652 0.501
R74683 out.n9669 out.n9668 0.501
R74684 out.n9668 out.n9667 0.501
R74685 out.n9667 out.n9666 0.501
R74686 out.n9666 out.n9665 0.501
R74687 out.n9665 out.n9664 0.501
R74688 out.n9664 out.n9663 0.501
R74689 out.n9663 out.n9662 0.501
R74690 out.n9662 out.n9661 0.501
R74691 out.n10011 out.t82 0.49
R74692 out.n2591 out.n2590 0.477
R74693 out.n2939 out.n2938 0.475
R74694 out.n2068 out.n2067 0.475
R74695 out.n1843 out.n1842 0.475
R74696 out.n2710 out.n2709 0.475
R74697 out.n1332 out.n1331 0.471
R74698 out.n14177 out.n14176 0.47
R74699 out.n10275 out.n10274 0.468
R74700 out.n12819 out.n12818 0.465
R74701 out.n13666 out.n13665 0.465
R74702 out.n13699 out.n13698 0.465
R74703 out.n11128 out.n11127 0.461
R74704 out.n11551 out.n11550 0.461
R74705 out.n12850 out.n12849 0.461
R74706 out.n11971 out.n11970 0.461
R74707 out.n10704 out.n10703 0.461
R74708 out.n12389 out.n12388 0.461
R74709 out.n2700 out.n2698 0.432
R74710 out.n1516 out.n1515 0.418
R74711 out.n2155 out.n2154 0.418
R74712 out.n2363 out.n2362 0.418
R74713 out.n10083 out.n10082 0.379
R74714 out.n13189 out.n13188 0.376
R74715 out.n13201 out.n13200 0.376
R74716 out.n12814 out.n12813 0.376
R74717 out.n12464 out.n12463 0.376
R74718 out.n12564 out.n12563 0.376
R74719 out.n12575 out.n12574 0.376
R74720 out.n12427 out.n12426 0.376
R74721 out.n12424 out.n12423 0.376
R74722 out.n12324 out.n12323 0.376
R74723 out.n12336 out.n12335 0.376
R74724 out.n13653 out.n13652 0.376
R74725 out.n13660 out.n13659 0.376
R74726 out.n13397 out.n13396 0.376
R74727 out.n13408 out.n13407 0.376
R74728 out.n13271 out.n13270 0.376
R74729 out.n13268 out.n13267 0.376
R74730 out.n11493 out.n11492 0.376
R74731 out.n11505 out.n11504 0.376
R74732 out.n11066 out.n11065 0.376
R74733 out.n11078 out.n11077 0.376
R74734 out.n11904 out.n11903 0.376
R74735 out.n11916 out.n11915 0.376
R74736 out.n13686 out.n13685 0.376
R74737 out.n13693 out.n13692 0.376
R74738 out.n13852 out.n13851 0.376
R74739 out.n13863 out.n13862 0.376
R74740 out.n13726 out.n13725 0.376
R74741 out.n13723 out.n13722 0.376
R74742 out.n10637 out.n10636 0.376
R74743 out.n10649 out.n10648 0.376
R74744 out.n14154 out.n14153 0.376
R74745 out.n14302 out.n14301 0.376
R74746 out.n14291 out.n14290 0.376
R74747 out.n14231 out.n14230 0.376
R74748 out.n14221 out.n14220 0.376
R74749 out.n4989 out.n4988 0.376
R74750 out.n4977 out.n4976 0.376
R74751 out.n5631 out.n5630 0.376
R74752 out.n5750 out.n5749 0.376
R74753 out.n5646 out.n5645 0.376
R74754 out.n2858 out.n2857 0.376
R74755 out.n5506 out.n5505 0.376
R74756 out.n5497 out.n5496 0.376
R74757 out.n1429 out.n1428 0.376
R74758 out.n5361 out.n5360 0.376
R74759 out.n6670 out.n6669 0.376
R74760 out.n6661 out.n6660 0.376
R74761 out.n6517 out.n6516 0.376
R74762 out.n6431 out.n6430 0.376
R74763 out.n6327 out.n6326 0.376
R74764 out.n6223 out.n6222 0.376
R74765 out.n1982 out.n1981 0.376
R74766 out.n6993 out.n6992 0.376
R74767 out.n6884 out.n6883 0.376
R74768 out.n6780 out.n6779 0.376
R74769 out.n1762 out.n1761 0.376
R74770 out.n7364 out.n7363 0.376
R74771 out.n7355 out.n7354 0.376
R74772 out.n2273 out.n2272 0.376
R74773 out.n7812 out.n7811 0.376
R74774 out.n7710 out.n7709 0.376
R74775 out.n7496 out.n7495 0.376
R74776 out.n7619 out.n7618 0.376
R74777 out.n5196 out.n5195 0.373
R74778 out.n7029 out.n7028 0.373
R74779 out.n12877 out.n12876 0.362
R74780 out.n12415 out.n12414 0.362
R74781 out.n12010 out.n12009 0.362
R74782 out.n13260 out.n13259 0.362
R74783 out.n11175 out.n11174 0.362
R74784 out.n10752 out.n10751 0.362
R74785 out.n11592 out.n11591 0.362
R74786 out.n13715 out.n13714 0.362
R74787 out.n10325 out.n10324 0.362
R74788 out.n5059 out.n5058 0.362
R74789 out.n5881 out.n5880 0.362
R74790 out.n14370 out.n14369 0.362
R74791 out.n10080 out.n10079 0.351
R74792 out.n5183 out.n5182 0.351
R74793 out.n10013 out.n10012 0.338
R74794 out.n10012 out.n10011 0.338
R74795 out.n9670 out.n9669 0.338
R74796 out.n9671 out.n9660 0.336
R74797 out.n5168 out.n4956 0.306
R74798 out.n10133 out.n10132 0.298
R74799 out.n12567 out.n12566 0.261
R74800 out.n13400 out.n13399 0.261
R74801 out.n13855 out.n13854 0.261
R74802 out.n14218 out.n14217 0.261
R74803 out.n2848 out.n2847 0.261
R74804 out.n1972 out.n1971 0.261
R74805 out.n1752 out.n1751 0.261
R74806 out.n7544 out.n7543 0.261
R74807 out.n11974 out.n11973 0.255
R74808 out.n10707 out.n10706 0.255
R74809 out.n12853 out.n12852 0.252
R74810 out.n12392 out.n12391 0.252
R74811 out.n11554 out.n11553 0.252
R74812 out.n11131 out.n11130 0.252
R74813 out.n1219 out.n1218 0.25
R74814 out.n7041 out.n7040 0.25
R74815 out.n10211 out.n10210 0.247
R74816 out.n12822 out.n12821 0.245
R74817 out.n13669 out.n13668 0.245
R74818 out.n13702 out.n13701 0.245
R74819 out.n1599 out.n1598 0.238
R74820 out.t85 out.t66 0.225
R74821 out.t71 out.t85 0.225
R74822 out.t83 out.t71 0.225
R74823 out.t82 out.t83 0.225
R74824 out.t84 out.t72 0.225
R74825 out.t70 out.t84 0.225
R74826 out.t80 out.t70 0.225
R74827 out.t79 out.t80 0.225
R74828 out.t78 out.t81 0.225
R74829 out.t68 out.t78 0.225
R74830 out.t76 out.t68 0.225
R74831 out.t75 out.t76 0.225
R74832 out.t77 out.t69 0.225
R74833 out.t67 out.t77 0.225
R74834 out.t74 out.t67 0.225
R74835 out.t73 out.t74 0.225
R74836 out.n1125 out.n1124 0.216
R74837 out.n9484 out.n9483 0.205
R74838 out.n9497 out.n9496 0.205
R74839 out.n9503 out.n9502 0.205
R74840 out.n9469 out.n9424 0.202
R74841 out.n9464 out.n9463 0.198
R74842 out.n10253 out.n10252 0.189
R74843 out.n12832 out.n12831 0.189
R74844 out.n12810 out.n12809 0.189
R74845 out.n12373 out.n12372 0.189
R74846 out.n13646 out.n13645 0.189
R74847 out.n11544 out.n11543 0.189
R74848 out.n11117 out.n11116 0.189
R74849 out.n11953 out.n11952 0.189
R74850 out.n13679 out.n13678 0.189
R74851 out.n10686 out.n10685 0.189
R74852 out.n14538 out.n14537 0.189
R74853 out.n5580 out.n5579 0.189
R74854 out.n6734 out.n6733 0.189
R74855 out.n7438 out.n7437 0.189
R74856 out.n7788 out.n7787 0.189
R74857 out.n7806 out.n7805 0.189
R74858 out.n10072 out.n10071 0.188
R74859 out.n10054 out.n10053 0.188
R74860 out.n5833 out.n5832 0.188
R74861 out.n2936 out.n2935 0.188
R74862 out.n6405 out.n6404 0.188
R74863 out.n2065 out.n2064 0.188
R74864 out.n6967 out.n6966 0.188
R74865 out.n1840 out.n1839 0.188
R74866 out.n2588 out.n2587 0.188
R74867 out.n9454 out.t0 0.186
R74868 out.n17312 out 0.185
R74869 out.n10077 out.n10075 0.185
R74870 out.n10059 out.n10058 0.185
R74871 out.n12993 out.n12991 0.185
R74872 out.n12128 out.n12126 0.185
R74873 out.n11305 out.n11303 0.185
R74874 out.n10875 out.n10873 0.185
R74875 out.n11708 out.n11706 0.185
R74876 out.n10441 out.n10439 0.185
R74877 out.n1005 out.n1003 0.185
R74878 out.n2743 out.n2741 0.185
R74879 out.n5402 out.n5400 0.185
R74880 out.n1145 out.n1143 0.185
R74881 out.n5180 out.n5178 0.185
R74882 out.n6471 out.n6469 0.185
R74883 out.n1872 out.n1870 0.185
R74884 out.n5889 out.n5887 0.185
R74885 out.n1647 out.n1645 0.185
R74886 out.n7263 out.n7261 0.185
R74887 out.n2492 out.n2490 0.185
R74888 out.n9466 out.n9465 0.18
R74889 out.n10258 out.n10257 0.178
R74890 out.n13219 out.n13218 0.178
R74891 out.n12658 out.n12657 0.178
R74892 out.n12354 out.n12353 0.178
R74893 out.n13491 out.n13490 0.178
R74894 out.n11523 out.n11522 0.178
R74895 out.n11096 out.n11095 0.178
R74896 out.n11934 out.n11933 0.178
R74897 out.n13946 out.n13945 0.178
R74898 out.n10667 out.n10666 0.178
R74899 out.n14481 out.n14480 0.178
R74900 out.n7779 out.n7778 0.178
R74901 out.n9673 out.n9672 0.177
R74902 out.n10241 out.n10240 0.177
R74903 out.n5155 out.n5154 0.177
R74904 out.n5824 out.n5823 0.177
R74905 out.n1328 out.n1327 0.177
R74906 out.n6396 out.n6395 0.177
R74907 out.n6958 out.n6957 0.177
R74908 out.n7208 out.n7207 0.177
R74909 out.n9469 out.n9466 0.169
R74910 out.n5380 out.n5379 0.166
R74911 out.n12812 out.n12811 0.155
R74912 out.n13648 out.n13647 0.155
R74913 out.n13681 out.n13680 0.155
R74914 out.n14547 out.n14546 0.155
R74915 out.n5571 out.n5570 0.155
R74916 out.n6725 out.n6724 0.155
R74917 out.n7429 out.n7428 0.155
R74918 out.n15388 out.n15387 0.154
R74919 out.n12649 out.n12648 0.144
R74920 out.n13482 out.n13481 0.144
R74921 out.n13937 out.n13936 0.144
R74922 out.n13228 out.n13227 0.144
R74923 out.n12363 out.n12362 0.144
R74924 out.n11532 out.n11531 0.144
R74925 out.n11105 out.n11104 0.144
R74926 out.n11943 out.n11942 0.144
R74927 out.n10676 out.n10675 0.144
R74928 out.n14490 out.n14489 0.144
R74929 out.n5164 out.n5163 0.144
R74930 out.n9671 out.n9670 0.139
R74931 out.n10012 out.t75 0.138
R74932 out.n10011 out.t79 0.137
R74933 out.n10013 out.t73 0.137
R74934 out.n12762 out.n12761 0.133
R74935 out.n13596 out.n13595 0.133
R74936 out.n14051 out.n14050 0.133
R74937 out.n10193 out.n10192 0.133
R74938 out.n13100 out.n13099 0.132
R74939 out.n12235 out.n12234 0.132
R74940 out.n11409 out.n11408 0.132
R74941 out.n10982 out.n10981 0.132
R74942 out.n11815 out.n11814 0.132
R74943 out.n10548 out.n10547 0.132
R74944 out.n14155 out.n14154 0.132
R74945 out.n1118 out.n1117 0.132
R74946 out.n13097 out.n13095 0.127
R74947 out.n12232 out.n12230 0.127
R74948 out.n11406 out.n11404 0.127
R74949 out.n10979 out.n10977 0.127
R74950 out.n11812 out.n11810 0.127
R74951 out.n10545 out.n10543 0.127
R74952 out.n14430 out.n14354 0.127
R74953 out.n5104 out.n5043 0.127
R74954 out.n12675 out.n12673 0.124
R74955 out.n13508 out.n13506 0.124
R74956 out.n13963 out.n13961 0.124
R74957 out.n13071 out.n13070 0.122
R74958 out.n12206 out.n12205 0.122
R74959 out.n11380 out.n11379 0.122
R74960 out.n10953 out.n10952 0.122
R74961 out.n11786 out.n11785 0.122
R74962 out.n10519 out.n10518 0.122
R74963 out.n14157 out.n14156 0.122
R74964 out.n1120 out.n1119 0.122
R74965 out.n12802 out.n12801 0.121
R74966 out.n13636 out.n13635 0.121
R74967 out.n14091 out.n14090 0.121
R74968 out.n6163 out.n6162 0.121
R74969 out.n5276 out.n5274 0.12
R74970 out.n9652 out.t7 0.111
R74971 out.n9653 out.t18 0.111
R74972 out.n9654 out.t4 0.111
R74973 out.n9655 out.t2 0.111
R74974 out.n9656 out.t13 0.111
R74975 out.n9657 out.t11 0.111
R74976 out.n9658 out.t10 0.111
R74977 out.n9659 out.t16 0.111
R74978 out.n9660 out.t14 0.111
R74979 out.n9661 out.t19 0.111
R74980 out.n9662 out.t21 0.111
R74981 out.n9663 out.t20 0.111
R74982 out.n9664 out.t5 0.111
R74983 out.n9665 out.t6 0.111
R74984 out.n9666 out.t12 0.111
R74985 out.n9667 out.t17 0.111
R74986 out.n9668 out.t3 0.111
R74987 out.n9669 out.t8 0.111
R74988 out.n13183 out.n13182 0.11
R74989 out.n12318 out.n12317 0.11
R74990 out.n11487 out.n11486 0.11
R74991 out.n11060 out.n11059 0.11
R74992 out.n11898 out.n11897 0.11
R74993 out.n10631 out.n10630 0.11
R74994 out.n4983 out.n4982 0.11
R74995 out.n12679 out.n12678 0.11
R74996 out.n13513 out.n13512 0.11
R74997 out.n13968 out.n13967 0.11
R74998 out.n10137 out.n10136 0.109
R74999 out.n5853 out.n5851 0.105
R75000 out.n5264 out.n5262 0.105
R75001 out.n6425 out.n6423 0.105
R75002 out.n6987 out.n6985 0.105
R75003 out.n7233 out.n7231 0.105
R75004 out.n7804 out.n7802 0.105
R75005 out.n14472 out.n14294 0.103
R75006 out.n5146 out.n4980 0.103
R75007 out.n13103 out.n13097 0.099
R75008 out.n11818 out.n11812 0.099
R75009 out.n10551 out.n10545 0.099
R75010 out.n11412 out.n11411 0.098
R75011 out.n10985 out.n10984 0.098
R75012 out.n12986 out.n12984 0.098
R75013 out.n12561 out.n12559 0.098
R75014 out.n12121 out.n12119 0.098
R75015 out.n13394 out.n13392 0.098
R75016 out.n11298 out.n11296 0.098
R75017 out.n10868 out.n10866 0.098
R75018 out.n11701 out.n11699 0.098
R75019 out.n13849 out.n13847 0.098
R75020 out.n10434 out.n10432 0.098
R75021 out.n5730 out.n5728 0.098
R75022 out.n6307 out.n6305 0.098
R75023 out.n6089 out.n6087 0.098
R75024 out.n6864 out.n6862 0.098
R75025 out.n7126 out.n7124 0.098
R75026 out.n7701 out.n7518 0.098
R75027 out.n12238 out.n12237 0.098
R75028 out.n13103 out.n13102 0.098
R75029 out.n11818 out.n11817 0.098
R75030 out.n10551 out.n10550 0.098
R75031 out.n14343 out.n14342 0.098
R75032 out.n5030 out.n5029 0.098
R75033 out.n1493 out.n1407 0.097
R75034 out.n5454 out.n5453 0.097
R75035 out.n2340 out.n2251 0.097
R75036 out.n7312 out.n7311 0.097
R75037 out.n12238 out.n12232 0.097
R75038 out.n13603 out.n13593 0.097
R75039 out.n14058 out.n14048 0.097
R75040 out.n13192 out.n13180 0.095
R75041 out.n11907 out.n11895 0.095
R75042 out.n10640 out.n10628 0.095
R75043 out.n14529 out.n14191 0.094
R75044 out.n1270 out.n1193 0.094
R75045 out.n10985 out.n10979 0.094
R75046 out.n12327 out.n12315 0.093
R75047 out.n13516 out.n13508 0.093
R75048 out.n13971 out.n13963 0.093
R75049 out.n1062 out.n986 0.093
R75050 out.n14476 out.n14276 0.093
R75051 out.n5150 out.n4962 0.093
R75052 out.n10188 out.n10179 0.092
R75053 out.n12769 out.n12759 0.092
R75054 out.n11412 out.n11406 0.092
R75055 out.n10130 out.n10121 0.091
R75056 out.n11069 out.n11057 0.091
R75057 out.n10107 out.n10105 0.091
R75058 out.n5743 out.n5741 0.091
R75059 out.n5489 out.n5487 0.091
R75060 out.n6653 out.n6651 0.091
R75061 out.n6320 out.n6318 0.091
R75062 out.n5987 out.n5985 0.091
R75063 out.n6877 out.n6875 0.091
R75064 out.n7347 out.n7345 0.091
R75065 out.n7139 out.n7137 0.091
R75066 out.n7703 out.n7509 0.091
R75067 out.n7609 out.n7569 0.091
R75068 out.n5444 out.n5420 0.091
R75069 out.n7302 out.n7281 0.091
R75070 out.n2929 out.n2745 0.09
R75071 out.n2895 out.n2853 0.09
R75072 out.n2058 out.n1874 0.09
R75073 out.n2019 out.n1977 0.09
R75074 out.n1833 out.n1649 0.09
R75075 out.n1799 out.n1757 0.09
R75076 out.n2907 out.n2906 0.09
R75077 out.n1491 out.n1414 0.09
R75078 out.n1811 out.n1810 0.09
R75079 out.n2338 out.n2258 0.09
R75080 out.n12682 out.n12675 0.09
R75081 out.n11496 out.n11484 0.09
R75082 out.n14523 out.n14216 0.09
R75083 out.n5284 out.n5276 0.089
R75084 out.n6074 out.n6067 0.089
R75085 out.n6540 out.n6533 0.089
R75086 out.n6635 out.n6628 0.089
R75087 out.n2124 out.n2123 0.089
R75088 out.n5964 out.n5957 0.089
R75089 out.n7594 out.n7593 0.089
R75090 out.n6619 out.n6618 0.089
R75091 out.n14527 out.n14198 0.088
R75092 out.n1060 out.n993 0.088
R75093 out.n2031 out.n2030 0.088
R75094 out.n10107 out.n10101 0.088
R75095 out.n13083 out.n13082 0.088
R75096 out.n12970 out.n12969 0.088
R75097 out.n11798 out.n11797 0.088
R75098 out.n11685 out.n11684 0.088
R75099 out.n10531 out.n10530 0.088
R75100 out.n10418 out.n10417 0.088
R75101 out.n13214 out.n13206 0.088
R75102 out.n11929 out.n11921 0.088
R75103 out.n10662 out.n10654 0.088
R75104 out.n7695 out.n7688 0.088
R75105 out.n2663 out.n2662 0.088
R75106 out.n1056 out.n1011 0.087
R75107 out.n7804 out.n7799 0.087
R75108 out.n2929 out.n2746 0.087
R75109 out.n1833 out.n1650 0.087
R75110 out.n1322 out.n1147 0.087
R75111 out.n1259 out.n1224 0.087
R75112 out.n2581 out.n2404 0.087
R75113 out.n2534 out.n2494 0.087
R75114 out.n1054 out.n1018 0.087
R75115 out.n1489 out.n1421 0.087
R75116 out.n5442 out.n5430 0.087
R75117 out.n2336 out.n2265 0.087
R75118 out.n7300 out.n7291 0.087
R75119 out.n2552 out.n2551 0.086
R75120 out.n1322 out.n1148 0.086
R75121 out.n2545 out.n2544 0.086
R75122 out.n10188 out.n10187 0.086
R75123 out.n1483 out.n1441 0.086
R75124 out.n2330 out.n2285 0.086
R75125 out.n14415 out.n14371 0.086
R75126 out.n5089 out.n5060 0.086
R75127 out.n14521 out.n14224 0.086
R75128 out.n14470 out.n14304 0.086
R75129 out.n5144 out.n4991 0.086
R75130 out.n7704 out.n7703 0.085
R75131 out.n12218 out.n12217 0.085
R75132 out.n12105 out.n12104 0.085
R75133 out.n13625 out.n13617 0.085
R75134 out.n13376 out.n13375 0.085
R75135 out.n14080 out.n14072 0.085
R75136 out.n13831 out.n13830 0.085
R75137 out.n12682 out.n12681 0.085
R75138 out.n12349 out.n12341 0.085
R75139 out.n13497 out.n13496 0.085
R75140 out.n13952 out.n13951 0.085
R75141 out.n7220 out.n7219 0.085
R75142 out.n2547 out.n2546 0.085
R75143 out.n13516 out.n13515 0.085
R75144 out.n13971 out.n13970 0.085
R75145 out.n2058 out.n1875 0.084
R75146 out.n1483 out.n1440 0.084
R75147 out.n6557 out.n6518 0.084
R75148 out.n2330 out.n2284 0.084
R75149 out.n7611 out.n7560 0.084
R75150 out.n2129 out.n2128 0.084
R75151 out.n1570 out.n1569 0.084
R75152 out.n6543 out.n6542 0.084
R75153 out.n6617 out.n6606 0.084
R75154 out.n5972 out.n5965 0.084
R75155 out.n10965 out.n10964 0.084
R75156 out.n10852 out.n10851 0.084
R75157 out.n6412 out.n6411 0.084
R75158 out.n11091 out.n11083 0.083
R75159 out.n5251 out.n5250 0.083
R75160 out.n2033 out.n2032 0.083
R75161 out.n7666 out.n7655 0.083
R75162 out.n1487 out.n1426 0.083
R75163 out.n2334 out.n2270 0.083
R75164 out.n10188 out.n10186 0.083
R75165 out.n10130 out.n10128 0.083
R75166 out.n14523 out.n14223 0.083
R75167 out.n7697 out.n7696 0.083
R75168 out.n2555 out.n2554 0.083
R75169 out.n7612 out.n7611 0.083
R75170 out.n12973 out.n12972 0.082
R75171 out.n12954 out.n12943 0.082
R75172 out.n11688 out.n11687 0.082
R75173 out.n11669 out.n11658 0.082
R75174 out.n10421 out.n10420 0.082
R75175 out.n10402 out.n10391 0.082
R75176 out.n6723 out.n6713 0.082
R75177 out.n6637 out.n6636 0.082
R75178 out.n6076 out.n6075 0.082
R75179 out.n6051 out.n6040 0.082
R75180 out.n2666 out.n2665 0.082
R75181 out.n7603 out.n7596 0.082
R75182 out.n12791 out.n12783 0.082
R75183 out.n12543 out.n12542 0.082
R75184 out.n11392 out.n11391 0.082
R75185 out.n11282 out.n11281 0.082
R75186 out.n5840 out.n5839 0.082
R75187 out.n6974 out.n6973 0.082
R75188 out.n12664 out.n12663 0.082
R75189 out.n11518 out.n11510 0.082
R75190 out.n2909 out.n2908 0.082
R75191 out.n1813 out.n1812 0.082
R75192 out.n14413 out.n14380 0.082
R75193 out.n5087 out.n5069 0.082
R75194 out.n13402 out.n13394 0.082
R75195 out.n13857 out.n13849 0.082
R75196 out.n13114 out.n13105 0.081
R75197 out.n13004 out.n12997 0.081
R75198 out.n11829 out.n11820 0.081
R75199 out.n11719 out.n11712 0.081
R75200 out.n10562 out.n10553 0.081
R75201 out.n10452 out.n10445 0.081
R75202 out.n6101 out.n6092 0.081
R75203 out.n14176 out.n14166 0.081
R75204 out.n1052 out.n1027 0.081
R75205 out.n2581 out.n2579 0.081
R75206 out.n12995 out.n12986 0.081
R75207 out.n11710 out.n11701 0.081
R75208 out.n10443 out.n10434 0.081
R75209 out.n6090 out.n6089 0.081
R75210 out.n13238 out.n13230 0.08
R75211 out.n12089 out.n12078 0.08
R75212 out.n13360 out.n13350 0.08
R75213 out.n13815 out.n13805 0.08
R75214 out.n7081 out.n7072 0.08
R75215 out.n14468 out.n14313 0.08
R75216 out.n5142 out.n5000 0.08
R75217 out.n6546 out.n6545 0.08
R75218 out.n6605 out.n6597 0.08
R75219 out.n7654 out.n7646 0.08
R75220 out.n7605 out.n7604 0.08
R75221 out.n2138 out.n2131 0.08
R75222 out.n1573 out.n1572 0.08
R75223 out.n1056 out.n1010 0.08
R75224 out.n14519 out.n14233 0.08
R75225 out.n12108 out.n12107 0.08
R75226 out.n13379 out.n13378 0.08
R75227 out.n13834 out.n13833 0.08
R75228 out.n7113 out.n7112 0.08
R75229 out.n6654 out.n6653 0.08
R75230 out.n13069 out.n13059 0.08
R75231 out.n11784 out.n11774 0.08
R75232 out.n10517 out.n10507 0.08
R75233 out.n6161 out.n6151 0.08
R75234 out.n7140 out.n7139 0.08
R75235 out.n7770 out.n7760 0.08
R75236 out.n14411 out.n14387 0.08
R75237 out.n5085 out.n5076 0.08
R75238 out.n2048 out.n2043 0.08
R75239 out.n12130 out.n12121 0.08
R75240 out.n6558 out.n6557 0.08
R75241 out.n5533 out.n5532 0.08
R75242 out.n7391 out.n7390 0.08
R75243 out.n1317 out.n1157 0.079
R75244 out.n6262 out.n6251 0.079
R75245 out.n12249 out.n12240 0.079
R75246 out.n12139 out.n12132 0.079
R75247 out.n13592 out.n13582 0.079
R75248 out.n13480 out.n13470 0.079
R75249 out.n14047 out.n14037 0.079
R75250 out.n13935 out.n13925 0.079
R75251 out.n2562 out.n2557 0.079
R75252 out.n1085 out.n1084 0.079
R75253 out.n13179 out.n13169 0.079
R75254 out.n11894 out.n11884 0.079
R75255 out.n10627 out.n10617 0.079
R75256 out.n7795 out.n7794 0.079
R75257 out.n6321 out.n6320 0.079
R75258 out.n1606 out.n1544 0.079
R75259 out.n10836 out.n10825 0.079
R75260 out.n5974 out.n5973 0.079
R75261 out.n1259 out.n1257 0.079
R75262 out.n12942 out.n12932 0.079
R75263 out.n11657 out.n11647 0.079
R75264 out.n10390 out.n10380 0.079
R75265 out.n6712 out.n6704 0.079
R75266 out.n6640 out.n6639 0.079
R75267 out.n6039 out.n6029 0.079
R75268 out.n2669 out.n2668 0.079
R75269 out.n1304 out.n1299 0.079
R75270 out.n10877 out.n10868 0.079
R75271 out.n6744 out.n6743 0.078
R75272 out.n6180 out.n6179 0.078
R75273 out.n10855 out.n10854 0.078
R75274 out.n1268 out.n1266 0.078
R75275 out.n6294 out.n6293 0.078
R75276 out.n5779 out.n5778 0.078
R75277 out.n5526 out.n5525 0.078
R75278 out.n6913 out.n6912 0.078
R75279 out.n7384 out.n7383 0.078
R75280 out.n2569 out.n2564 0.078
R75281 out.n12204 out.n12194 0.078
R75282 out.n12664 out.n12435 0.078
R75283 out.n7715 out.n7706 0.078
R75284 out.n1092 out.n1087 0.078
R75285 out.n1311 out.n1306 0.078
R75286 out.n12314 out.n12304 0.078
R75287 out.n13527 out.n13518 0.078
R75288 out.n13413 out.n13404 0.078
R75289 out.n13982 out.n13973 0.078
R75290 out.n13868 out.n13859 0.078
R75291 out.n5251 out.n5190 0.078
R75292 out.n14503 out.n14498 0.078
R75293 out.n5203 out.n5202 0.078
R75294 out.n13497 out.n13279 0.078
R75295 out.n13952 out.n13734 0.078
R75296 out.n7220 out.n7023 0.078
R75297 out.n1606 out.n1604 0.078
R75298 out.n14441 out.n14436 0.078
R75299 out.n14409 out.n14403 0.078
R75300 out.n5115 out.n5110 0.078
R75301 out.n12527 out.n12517 0.078
R75302 out.n5569 out.n5559 0.078
R75303 out.n7427 out.n7417 0.078
R75304 out.n7695 out.n7694 0.078
R75305 out.n2663 out.n2659 0.078
R75306 out.n10991 out.n10987 0.078
R75307 out.n10886 out.n10879 0.078
R75308 out.n14466 out.n14458 0.078
R75309 out.n5140 out.n5132 0.078
R75310 out.n12543 out.n12452 0.078
R75311 out.n11392 out.n11167 0.078
R75312 out.n11282 out.n11190 0.078
R75313 out.n5840 out.n5639 0.078
R75314 out.n6974 out.n6773 0.078
R75315 out.n14174 out.n14172 0.078
R75316 out.n1050 out.n1048 0.078
R75317 out.n1104 out.n1102 0.078
R75318 out.n7759 out.n7751 0.078
R75319 out.n6540 out.n6539 0.078
R75320 out.n6635 out.n6634 0.078
R75321 out.n2124 out.n2111 0.078
R75322 out.n5964 out.n5963 0.078
R75323 out.n7594 out.n7582 0.078
R75324 out.n6596 out.n6590 0.078
R75325 out.n1580 out.n1575 0.078
R75326 out.n7645 out.n7637 0.078
R75327 out.n10965 out.n10744 0.078
R75328 out.n10852 out.n10764 0.078
R75329 out.n6412 out.n6211 0.078
R75330 out.n12218 out.n12002 0.077
R75331 out.n12105 out.n12022 0.077
R75332 out.n13376 out.n13296 0.077
R75333 out.n13831 out.n13751 0.077
R75334 out.n12569 out.n12561 0.077
R75335 out.n7111 out.n7110 0.077
R75336 out.n14517 out.n14510 0.077
R75337 out.n5988 out.n5987 0.077
R75338 out.n11266 out.n11255 0.077
R75339 out.n5685 out.n5674 0.077
R75340 out.n6819 out.n6808 0.077
R75341 out.n13083 out.n12869 0.077
R75342 out.n12970 out.n12889 0.077
R75343 out.n11798 out.n11584 0.077
R75344 out.n11685 out.n11604 0.077
R75345 out.n10531 out.n10317 0.077
R75346 out.n10418 out.n10337 0.077
R75347 out.n7071 out.n7063 0.077
R75348 out.n6292 out.n6291 0.077
R75349 out.n1922 out.n1921 0.077
R75350 out.n11307 out.n11298 0.077
R75351 out.n2534 out.n2532 0.077
R75352 out.n6074 out.n6073 0.077
R75353 out.n5715 out.n5714 0.077
R75354 out.n2798 out.n2797 0.077
R75355 out.n5471 out.n5470 0.077
R75356 out.n1390 out.n1389 0.077
R75357 out.n6849 out.n6848 0.077
R75358 out.n1702 out.n1701 0.077
R75359 out.n7329 out.n7328 0.077
R75360 out.n2234 out.n2233 0.077
R75361 out.n14506 out.n14505 0.077
R75362 out.n14447 out.n14443 0.077
R75363 out.n14457 out.n14451 0.077
R75364 out.n5121 out.n5117 0.077
R75365 out.n5131 out.n5125 0.077
R75366 out.n1099 out.n1094 0.077
R75367 out.n1245 out.n1240 0.077
R75368 out.n6351 out.n6350 0.077
R75369 out.n2443 out.n2442 0.077
R75370 out.n5744 out.n5743 0.077
R75371 out.n6878 out.n6877 0.077
R75372 out.n2923 out.n2762 0.077
R75373 out.n1511 out.n1363 0.077
R75374 out.n2150 out.n2097 0.077
R75375 out.n2052 out.n1891 0.077
R75376 out.n1827 out.n1666 0.077
R75377 out.n2358 out.n2207 0.077
R75378 out.n2573 out.n2419 0.077
R75379 out.n2688 out.n2637 0.077
R75380 out.n2520 out.n2515 0.077
R75381 out.n12077 out.n12067 0.077
R75382 out.n13349 out.n13341 0.077
R75383 out.n13804 out.n13796 0.077
R75384 out.n7199 out.n7189 0.077
R75385 out.n12546 out.n12545 0.077
R75386 out.n11285 out.n11284 0.077
R75387 out.n5717 out.n5716 0.077
R75388 out.n5473 out.n5472 0.077
R75389 out.n6851 out.n6850 0.077
R75390 out.n7331 out.n7330 0.077
R75391 out.n10951 out.n10941 0.077
R75392 out.n12758 out.n12748 0.077
R75393 out.n12647 out.n12637 0.077
R75394 out.n11418 out.n11414 0.077
R75395 out.n11313 out.n11309 0.077
R75396 out.n2019 out.n2017 0.077
R75397 out.n14362 out.n14361 0.077
R75398 out.n5051 out.n5050 0.077
R75399 out.n11056 out.n11046 0.077
R75400 out.n6553 out.n6548 0.077
R75401 out.n13058 out.n13050 0.076
R75402 out.n12931 out.n12923 0.076
R75403 out.n11773 out.n11765 0.076
R75404 out.n11646 out.n11638 0.076
R75405 out.n10506 out.n10498 0.076
R75406 out.n10379 out.n10371 0.076
R75407 out.n6703 out.n6695 0.076
R75408 out.n6150 out.n6142 0.076
R75409 out.n6028 out.n6020 0.076
R75410 out.n2676 out.n2671 0.076
R75411 out.n2543 out.n2541 0.076
R75412 out.n1113 out.n1111 0.076
R75413 out.n7149 out.n7142 0.076
R75414 out.n2145 out.n2140 0.076
R75415 out.n14402 out.n14396 0.076
R75416 out.n1044 out.n1039 0.076
R75417 out.n1481 out.n1447 0.076
R75418 out.n2328 out.n2291 0.076
R75419 out.n2931 out.n2738 0.076
R75420 out.n2898 out.n2846 0.076
R75421 out.n2060 out.n1867 0.076
R75422 out.n2022 out.n1970 0.076
R75423 out.n1835 out.n1642 0.076
R75424 out.n1802 out.n1750 0.076
R75425 out.n2707 out.n2628 0.076
R75426 out.n5232 out.n5222 0.076
R75427 out.n7170 out.n7169 0.076
R75428 out.n13125 out.n13116 0.076
R75429 out.n13015 out.n13006 0.076
R75430 out.n11840 out.n11831 0.076
R75431 out.n11730 out.n11721 0.076
R75432 out.n10573 out.n10564 0.076
R75433 out.n10463 out.n10454 0.076
R75434 out.n6112 out.n6103 0.076
R75435 out.n6000 out.n5993 0.076
R75436 out.n6589 out.n6583 0.076
R75437 out.n7750 out.n7742 0.076
R75438 out.n10824 out.n10814 0.075
R75439 out.n6387 out.n6377 0.075
R75440 out.n6250 out.n6242 0.075
R75441 out.n11378 out.n11368 0.075
R75442 out.n2895 out.n2893 0.075
R75443 out.n1799 out.n1797 0.075
R75444 out.n1587 out.n1582 0.075
R75445 out.n1320 out.n1318 0.075
R75446 out.n13168 out.n13158 0.075
R75447 out.n11883 out.n11873 0.075
R75448 out.n10616 out.n10606 0.075
R75449 out.n12066 out.n12058 0.075
R75450 out.n13340 out.n13332 0.075
R75451 out.n13795 out.n13787 0.075
R75452 out.n7062 out.n7054 0.075
R75453 out.n2028 out.n2026 0.075
R75454 out.n7168 out.n7167 0.075
R75455 out.n12693 out.n12684 0.075
R75456 out.n12580 out.n12571 0.075
R75457 out.n11483 out.n11473 0.075
R75458 out.n5295 out.n5286 0.075
R75459 out.n1256 out.n1254 0.075
R75460 out.n7724 out.n7717 0.075
R75461 out.n7628 out.n7624 0.075
R75462 out.n12193 out.n12185 0.075
R75463 out.n13469 out.n13459 0.075
R75464 out.n13924 out.n13914 0.075
R75465 out.n7188 out.n7180 0.075
R75466 out.n6675 out.n6666 0.075
R75467 out.n11254 out.n11244 0.074
R75468 out.n7636 out.n7635 0.074
R75469 out.n5490 out.n5489 0.074
R75470 out.n7348 out.n7347 0.074
R75471 out.n5284 out.n5283 0.074
R75472 out.n13049 out.n13041 0.074
R75473 out.n12922 out.n12916 0.074
R75474 out.n11764 out.n11756 0.074
R75475 out.n11637 out.n11631 0.074
R75476 out.n10497 out.n10489 0.074
R75477 out.n10370 out.n10364 0.074
R75478 out.n6694 out.n6688 0.074
R75479 out.n6141 out.n6133 0.074
R75480 out.n6019 out.n6013 0.074
R75481 out.n6582 out.n6576 0.074
R75482 out.n6687 out.n6686 0.074
R75483 out.n6012 out.n6011 0.074
R75484 out.n7741 out.n7735 0.074
R75485 out.n5349 out.n5339 0.074
R75486 out.n12516 out.n12508 0.074
R75487 out.n5815 out.n5805 0.074
R75488 out.n5673 out.n5665 0.074
R75489 out.n5558 out.n5550 0.074
R75490 out.n6949 out.n6939 0.074
R75491 out.n6807 out.n6799 0.074
R75492 out.n7416 out.n7408 0.074
R75493 out.n12260 out.n12251 0.074
R75494 out.n12150 out.n12141 0.074
R75495 out.n13581 out.n13571 0.074
R75496 out.n14036 out.n14026 0.074
R75497 out.n2151 out.n2150 0.074
R75498 out.n2683 out.n2678 0.074
R75499 out.n12303 out.n12293 0.074
R75500 out.n13538 out.n13529 0.074
R75501 out.n13993 out.n13984 0.074
R75502 out.n6332 out.n6323 0.074
R75503 out.n6241 out.n6233 0.074
R75504 out.n13424 out.n13415 0.074
R75505 out.n13879 out.n13870 0.074
R75506 out.n2904 out.n2902 0.073
R75507 out.n5476 out.n5475 0.073
R75508 out.n1808 out.n1806 0.073
R75509 out.n7334 out.n7333 0.073
R75510 out.n6685 out.n6684 0.073
R75511 out.n6010 out.n6009 0.073
R75512 out.n6125 out.n6124 0.073
R75513 out.n6376 out.n6368 0.073
R75514 out.n10940 out.n10932 0.073
R75515 out.n10813 out.n10805 0.073
R75516 out.n5221 out.n5213 0.073
R75517 out.n7179 out.n7171 0.073
R75518 out.n7730 out.n7726 0.073
R75519 out.n13132 out.n13127 0.073
R75520 out.n13040 out.n13034 0.073
R75521 out.n12915 out.n12909 0.073
R75522 out.n11847 out.n11842 0.073
R75523 out.n11755 out.n11749 0.073
R75524 out.n11630 out.n11624 0.073
R75525 out.n10580 out.n10575 0.073
R75526 out.n10488 out.n10482 0.073
R75527 out.n10363 out.n10357 0.073
R75528 out.n6132 out.n6126 0.073
R75529 out.n12184 out.n12176 0.073
R75530 out.n13331 out.n13325 0.073
R75531 out.n13786 out.n13780 0.073
R75532 out.n5264 out.n5184 0.073
R75533 out.n2583 out.n2396 0.073
R75534 out.n2537 out.n2488 0.073
R75535 out.n11002 out.n10993 0.073
R75536 out.n10897 out.n10888 0.073
R75537 out.n10775 out.n10768 0.073
R75538 out.n13157 out.n13149 0.073
R75539 out.n11872 out.n11864 0.073
R75540 out.n10605 out.n10597 0.073
R75541 out.n7634 out.n7633 0.073
R75542 out.n5590 out.n5589 0.073
R75543 out.n7448 out.n7447 0.073
R75544 out.n2688 out.n2686 0.073
R75545 out.n13023 out.n13017 0.073
R75546 out.n12899 out.n12895 0.073
R75547 out.n11738 out.n11732 0.073
R75548 out.n11614 out.n11610 0.073
R75549 out.n10471 out.n10465 0.073
R75550 out.n10347 out.n10343 0.073
R75551 out.n6120 out.n6114 0.073
R75552 out.n6006 out.n6002 0.073
R75553 out.n13458 out.n13450 0.073
R75554 out.n13913 out.n13905 0.073
R75555 out.n12057 out.n12051 0.073
R75556 out.n5755 out.n5746 0.073
R75557 out.n6889 out.n6880 0.073
R75558 out.n7158 out.n7151 0.072
R75559 out.n2528 out.n2526 0.072
R75560 out.n7622 out.n7614 0.072
R75561 out.n2055 out.n2054 0.072
R75562 out.n6681 out.n6677 0.072
R75563 out.n5804 out.n5796 0.072
R75564 out.n6938 out.n6930 0.072
R75565 out.n11045 out.n11035 0.072
R75566 out.n6664 out.n6656 0.072
R75567 out.n6566 out.n6560 0.072
R75568 out.n2926 out.n2925 0.072
R75569 out.n1830 out.n1829 0.072
R75570 out.n13138 out.n13134 0.072
R75571 out.n13148 out.n13142 0.072
R75572 out.n13033 out.n13027 0.072
R75573 out.n12908 out.n12902 0.072
R75574 out.n11853 out.n11849 0.072
R75575 out.n11863 out.n11857 0.072
R75576 out.n11748 out.n11742 0.072
R75577 out.n11623 out.n11617 0.072
R75578 out.n10586 out.n10582 0.072
R75579 out.n10596 out.n10590 0.072
R75580 out.n10481 out.n10475 0.072
R75581 out.n10356 out.n10350 0.072
R75582 out.n7734 out.n7733 0.072
R75583 out.n1262 out.n1217 0.072
R75584 out.n9438 out.n9437 0.072
R75585 out.n12849 out.n12847 0.072
R75586 out.n11970 out.n11968 0.072
R75587 out.n10703 out.n10701 0.072
R75588 out.n5212 out.n5204 0.072
R75589 out.n5991 out.n5990 0.072
R75590 out.n12636 out.n12626 0.072
R75591 out.n12507 out.n12499 0.072
R75592 out.n11367 out.n11359 0.072
R75593 out.n11243 out.n11235 0.072
R75594 out.n5664 out.n5656 0.072
R75595 out.n5549 out.n5541 0.072
R75596 out.n6798 out.n6790 0.072
R75597 out.n7407 out.n7399 0.072
R75598 out.n12175 out.n12169 0.072
R75599 out.n12050 out.n12044 0.072
R75600 out.n13449 out.n13443 0.072
R75601 out.n13904 out.n13898 0.072
R75602 out.n12267 out.n12262 0.071
R75603 out.n13570 out.n13564 0.071
R75604 out.n14025 out.n14019 0.071
R75605 out.n5304 out.n5297 0.071
R75606 out.n1253 out.n1251 0.071
R75607 out.n10931 out.n10923 0.071
R75608 out.n10804 out.n10798 0.071
R75609 out.n5338 out.n5330 0.071
R75610 out.n6367 out.n6359 0.071
R75611 out.n12292 out.n12284 0.071
R75612 out.n13547 out.n13540 0.071
R75613 out.n14002 out.n13995 0.071
R75614 out.n13665 out.n13663 0.071
R75615 out.n13698 out.n13696 0.071
R75616 out.n12747 out.n12737 0.071
R75617 out.n11429 out.n11420 0.071
R75618 out.n11324 out.n11315 0.071
R75619 out.n11205 out.n11198 0.071
R75620 out.n12158 out.n12152 0.071
R75621 out.n12034 out.n12030 0.071
R75622 out.n13432 out.n13426 0.071
R75623 out.n13308 out.n13304 0.071
R75624 out.n13887 out.n13881 0.071
R75625 out.n13763 out.n13759 0.071
R75626 out.n12704 out.n12695 0.071
R75627 out.n11472 out.n11462 0.071
R75628 out.n12591 out.n12582 0.071
R75629 out.n12469 out.n12460 0.071
R75630 out.n5511 out.n5502 0.071
R75631 out.n7369 out.n7360 0.071
R75632 out.n13324 out.n13318 0.071
R75633 out.n13779 out.n13773 0.071
R75634 out.n12273 out.n12269 0.071
R75635 out.n12283 out.n12277 0.071
R75636 out.n13553 out.n13549 0.071
R75637 out.n13563 out.n13557 0.071
R75638 out.n13317 out.n13311 0.071
R75639 out.n14008 out.n14004 0.071
R75640 out.n14018 out.n14012 0.071
R75641 out.n13772 out.n13766 0.071
R75642 out.n1512 out.n1511 0.071
R75643 out.n2359 out.n2358 0.071
R75644 out.n7164 out.n7160 0.07
R75645 out.n10922 out.n10916 0.07
R75646 out.n10797 out.n10791 0.07
R75647 out.n6341 out.n6334 0.07
R75648 out.n2013 out.n2011 0.07
R75649 out.n12498 out.n12492 0.07
R75650 out.n5540 out.n5534 0.07
R75651 out.n7398 out.n7392 0.07
R75652 out.n11009 out.n11004 0.07
R75653 out.n5329 out.n5321 0.07
R75654 out.n6358 out.n6352 0.07
R75655 out.n12625 out.n12617 0.07
R75656 out.n11034 out.n11026 0.07
R75657 out.n11358 out.n11350 0.07
R75658 out.n11234 out.n11228 0.07
R75659 out.n5795 out.n5787 0.07
R75660 out.n6929 out.n6921 0.07
R75661 out.n12388 out.n12386 0.07
R75662 out.n10130 out.n10129 0.07
R75663 out.n10107 out.n10106 0.07
R75664 out.n10905 out.n10899 0.07
R75665 out.n10781 out.n10777 0.07
R75666 out.n11127 out.n11125 0.07
R75667 out.n12168 out.n12162 0.07
R75668 out.n12043 out.n12037 0.07
R75669 out.n13442 out.n13436 0.07
R75670 out.n13897 out.n13891 0.07
R75671 out.n11025 out.n11019 0.069
R75672 out.n5764 out.n5757 0.069
R75673 out.n2889 out.n2887 0.069
R75674 out.n6898 out.n6891 0.069
R75675 out.n1793 out.n1791 0.069
R75676 out.n11015 out.n11011 0.069
R75677 out.n5320 out.n5315 0.069
R75678 out.n5311 out.n5306 0.069
R75679 out.n1250 out.n1248 0.069
R75680 out.n12736 out.n12730 0.069
R75681 out.n11436 out.n11431 0.069
R75682 out.n11349 out.n11343 0.069
R75683 out.n6347 out.n6343 0.069
R75684 out.n10120 out.n10118 0.069
R75685 out.n13085 out.n12863 0.069
R75686 out.n13148 out.n13146 0.069
R75687 out.n13205 out.n13203 0.069
R75688 out.n13214 out.n13212 0.069
R75689 out.n13033 out.n13031 0.069
R75690 out.n13040 out.n13038 0.069
R75691 out.n12849 out.n12839 0.069
R75692 out.n12908 out.n12906 0.069
R75693 out.n12915 out.n12913 0.069
R75694 out.n12922 out.n12920 0.069
R75695 out.n12666 out.n12429 0.069
R75696 out.n12729 out.n12727 0.069
R75697 out.n12736 out.n12734 0.069
R75698 out.n12782 out.n12780 0.069
R75699 out.n12791 out.n12789 0.069
R75700 out.n12609 out.n12607 0.069
R75701 out.n12616 out.n12614 0.069
R75702 out.n12818 out.n12816 0.069
R75703 out.n12484 out.n12482 0.069
R75704 out.n12491 out.n12489 0.069
R75705 out.n12498 out.n12496 0.069
R75706 out.n12220 out.n11996 0.069
R75707 out.n12283 out.n12281 0.069
R75708 out.n12340 out.n12338 0.069
R75709 out.n12349 out.n12347 0.069
R75710 out.n12168 out.n12166 0.069
R75711 out.n12175 out.n12173 0.069
R75712 out.n12388 out.n12380 0.069
R75713 out.n12043 out.n12041 0.069
R75714 out.n12050 out.n12048 0.069
R75715 out.n12057 out.n12055 0.069
R75716 out.n13499 out.n13273 0.069
R75717 out.n13563 out.n13561 0.069
R75718 out.n13570 out.n13568 0.069
R75719 out.n13616 out.n13614 0.069
R75720 out.n13625 out.n13623 0.069
R75721 out.n13442 out.n13440 0.069
R75722 out.n13449 out.n13447 0.069
R75723 out.n13665 out.n13655 0.069
R75724 out.n13317 out.n13315 0.069
R75725 out.n13324 out.n13322 0.069
R75726 out.n13331 out.n13329 0.069
R75727 out.n11394 out.n11161 0.069
R75728 out.n11452 out.n11450 0.069
R75729 out.n11509 out.n11507 0.069
R75730 out.n11518 out.n11516 0.069
R75731 out.n11342 out.n11340 0.069
R75732 out.n11349 out.n11347 0.069
R75733 out.n11550 out.n11548 0.069
R75734 out.n11220 out.n11218 0.069
R75735 out.n11227 out.n11225 0.069
R75736 out.n11234 out.n11232 0.069
R75737 out.n10967 out.n10738 0.069
R75738 out.n11025 out.n11023 0.069
R75739 out.n11082 out.n11080 0.069
R75740 out.n11091 out.n11089 0.069
R75741 out.n10915 out.n10913 0.069
R75742 out.n10922 out.n10920 0.069
R75743 out.n11127 out.n11124 0.069
R75744 out.n10790 out.n10788 0.069
R75745 out.n10797 out.n10795 0.069
R75746 out.n10804 out.n10802 0.069
R75747 out.n11800 out.n11578 0.069
R75748 out.n11863 out.n11861 0.069
R75749 out.n11920 out.n11918 0.069
R75750 out.n11929 out.n11927 0.069
R75751 out.n11748 out.n11746 0.069
R75752 out.n11755 out.n11753 0.069
R75753 out.n11970 out.n11960 0.069
R75754 out.n11623 out.n11621 0.069
R75755 out.n11630 out.n11628 0.069
R75756 out.n11637 out.n11635 0.069
R75757 out.n13954 out.n13728 0.069
R75758 out.n14018 out.n14016 0.069
R75759 out.n14025 out.n14023 0.069
R75760 out.n14071 out.n14069 0.069
R75761 out.n14080 out.n14078 0.069
R75762 out.n13897 out.n13895 0.069
R75763 out.n13904 out.n13902 0.069
R75764 out.n13698 out.n13688 0.069
R75765 out.n13772 out.n13770 0.069
R75766 out.n13779 out.n13777 0.069
R75767 out.n13786 out.n13784 0.069
R75768 out.n10533 out.n10311 0.069
R75769 out.n10596 out.n10594 0.069
R75770 out.n10653 out.n10651 0.069
R75771 out.n10662 out.n10660 0.069
R75772 out.n10481 out.n10479 0.069
R75773 out.n10488 out.n10486 0.069
R75774 out.n10703 out.n10693 0.069
R75775 out.n10356 out.n10354 0.069
R75776 out.n10363 out.n10361 0.069
R75777 out.n10370 out.n10368 0.069
R75778 out.n14525 out.n14215 0.069
R75779 out.n14527 out.n14204 0.069
R75780 out.n14529 out.n14197 0.069
R75781 out.n14428 out.n14355 0.069
R75782 out.n14457 out.n14455 0.069
R75783 out.n14474 out.n14293 0.069
R75784 out.n14476 out.n14282 0.069
R75785 out.n14402 out.n14400 0.069
R75786 out.n14409 out.n14407 0.069
R75787 out.n5102 out.n5044 0.069
R75788 out.n5131 out.n5129 0.069
R75789 out.n5148 out.n4979 0.069
R75790 out.n5150 out.n4968 0.069
R75791 out.n1062 out.n985 0.069
R75792 out.n1060 out.n992 0.069
R75793 out.n1058 out.n1001 0.069
R75794 out.n1113 out.n943 0.069
R75795 out.n1104 out.n946 0.069
R75796 out.n5786 out.n5784 0.069
R75797 out.n5779 out.n5777 0.069
R75798 out.n2886 out.n2869 0.069
R75799 out.n2889 out.n2863 0.069
R75800 out.n2892 out.n2860 0.069
R75801 out.n2901 out.n2836 0.069
R75802 out.n2904 out.n2828 0.069
R75803 out.n2907 out.n2822 0.069
R75804 out.n2925 out.n2755 0.069
R75805 out.n1491 out.n1413 0.069
R75806 out.n1489 out.n1420 0.069
R75807 out.n1487 out.n1425 0.069
R75808 out.n1485 out.n1433 0.069
R75809 out.n1481 out.n1446 0.069
R75810 out.n1474 out.n1453 0.069
R75811 out.n5440 out.n5439 0.069
R75812 out.n5540 out.n5538 0.069
R75813 out.n5533 out.n5531 0.069
R75814 out.n5526 out.n5524 0.069
R75815 out.n1320 out.n1153 0.069
R75816 out.n5320 out.n5318 0.069
R75817 out.n5203 out.n5201 0.069
R75818 out.n1250 out.n1239 0.069
R75819 out.n1265 out.n1207 0.069
R75820 out.n1268 out.n1199 0.069
R75821 out.n1270 out.n1192 0.069
R75822 out.n5364 out.n5363 0.069
R75823 out.n1317 out.n1156 0.069
R75824 out.n1315 out.n1163 0.069
R75825 out.n6575 out.n6504 0.069
R75826 out.n6582 out.n6580 0.069
R75827 out.n6589 out.n6587 0.069
R75828 out.n6596 out.n6594 0.069
R75829 out.n6694 out.n6692 0.069
R75830 out.n6687 out.n6463 0.069
R75831 out.n6685 out.n6468 0.069
R75832 out.n6358 out.n6356 0.069
R75833 out.n6351 out.n6218 0.069
R75834 out.n2010 out.n1993 0.069
R75835 out.n2013 out.n1987 0.069
R75836 out.n2016 out.n1984 0.069
R75837 out.n2025 out.n1960 0.069
R75838 out.n2028 out.n1952 0.069
R75839 out.n2031 out.n1946 0.069
R75840 out.n2054 out.n1884 0.069
R75841 out.n6132 out.n6130 0.069
R75842 out.n6125 out.n5886 0.069
R75843 out.n6019 out.n6017 0.069
R75844 out.n6012 out.n5909 0.069
R75845 out.n6010 out.n5914 0.069
R75846 out.n1592 out.n1550 0.069
R75847 out.n6920 out.n6918 0.069
R75848 out.n6913 out.n6911 0.069
R75849 out.n1790 out.n1773 0.069
R75850 out.n1793 out.n1767 0.069
R75851 out.n1796 out.n1764 0.069
R75852 out.n1805 out.n1740 0.069
R75853 out.n1808 out.n1732 0.069
R75854 out.n1811 out.n1726 0.069
R75855 out.n1829 out.n1659 0.069
R75856 out.n2338 out.n2257 0.069
R75857 out.n2336 out.n2264 0.069
R75858 out.n2334 out.n2269 0.069
R75859 out.n2332 out.n2277 0.069
R75860 out.n2328 out.n2290 0.069
R75861 out.n2321 out.n2297 0.069
R75862 out.n7398 out.n7396 0.069
R75863 out.n7391 out.n7389 0.069
R75864 out.n7384 out.n7382 0.069
R75865 out.n7170 out.n7034 0.069
R75866 out.n7168 out.n7039 0.069
R75867 out.n2525 out.n2508 0.069
R75868 out.n2528 out.n2502 0.069
R75869 out.n2531 out.n2499 0.069
R75870 out.n2543 out.n2476 0.069
R75871 out.n2545 out.n2469 0.069
R75872 out.n2575 out.n2412 0.069
R75873 out.n7741 out.n7739 0.069
R75874 out.n7734 out.n7491 0.069
R75875 out.n7636 out.n7530 0.069
R75876 out.n7634 out.n7535 0.069
R75877 out.n7632 out.n7542 0.069
R75878 out.n2691 out.n2633 0.069
R75879 out.n2531 out.n2529 0.069
R75880 out.n11332 out.n11326 0.069
R75881 out.n11211 out.n11207 0.069
R75882 out.n5786 out.n5780 0.069
R75883 out.n6920 out.n6914 0.069
R75884 out.n12713 out.n12706 0.069
R75885 out.n12616 out.n12610 0.069
R75886 out.n11461 out.n11453 0.069
R75887 out.n10915 out.n10909 0.068
R75888 out.n10790 out.n10784 0.068
R75889 out.n12599 out.n12593 0.068
R75890 out.n12475 out.n12471 0.068
R75891 out.n5517 out.n5513 0.068
R75892 out.n7375 out.n7371 0.068
R75893 out.n12491 out.n12485 0.068
R75894 out.n11227 out.n11221 0.068
R75895 out.n5500 out.n5492 0.068
R75896 out.n7358 out.n7350 0.068
R75897 out.n1525 out.n1346 0.068
R75898 out.n2164 out.n2082 0.068
R75899 out.n2372 out.n2190 0.068
R75900 out.n2540 out.n2482 0.068
R75901 out.n12719 out.n12715 0.068
R75902 out.n12729 out.n12723 0.068
R75903 out.n11442 out.n11438 0.068
R75904 out.n11452 out.n11446 0.068
R75905 out.n5957 out.n5938 0.068
R75906 out.n5770 out.n5766 0.068
R75907 out.n6904 out.n6900 0.068
R75908 out.n2016 out.n2014 0.067
R75909 out.n7804 out.n7803 0.067
R75910 out.n12609 out.n12603 0.067
R75911 out.n12484 out.n12478 0.067
R75912 out.n11342 out.n11336 0.067
R75913 out.n11220 out.n11214 0.067
R75914 out.n2895 out.n2894 0.067
R75915 out.n1799 out.n1798 0.067
R75916 out.n7593 out.n7585 0.067
R75917 out.n2892 out.n2890 0.066
R75918 out.n1796 out.n1794 0.066
R75919 out.n6628 out.n6620 0.066
R75920 out.n13157 out.n13155 0.066
R75921 out.n12292 out.n12290 0.066
R75922 out.n11461 out.n11459 0.066
R75923 out.n11034 out.n11032 0.066
R75924 out.n11872 out.n11870 0.066
R75925 out.n10605 out.n10603 0.066
R75926 out.n14517 out.n14515 0.066
R75927 out.n14466 out.n14464 0.066
R75928 out.n5140 out.n5138 0.066
R75929 out.n5338 out.n5336 0.066
R75930 out.n2019 out.n2018 0.066
R75931 out.n5956 out.n5949 0.066
R75932 out.n11309 out.n11308 0.065
R75933 out.n11496 out.n11495 0.065
R75934 out.n11406 out.n11405 0.065
R75935 out.n15160 out.n10042 0.065
R75936 out.n10879 out.n10878 0.064
R75937 out.n5373 out.n5365 0.064
R75938 out.n1259 out.n1258 0.064
R75939 out.n12769 out.n12768 0.064
R75940 out.n12675 out.n12674 0.064
R75941 out.n11069 out.n11068 0.064
R75942 out.n10979 out.n10978 0.064
R75943 out.n14430 out.n14346 0.064
R75944 out.n5104 out.n5034 0.064
R75945 out.n5276 out.n5275 0.064
R75946 out.n12571 out.n12570 0.064
R75947 out.n5746 out.n5745 0.064
R75948 out.n6880 out.n6879 0.064
R75949 out.n2549 out.n2548 0.064
R75950 out.n5463 out.n5455 0.063
R75951 out.n7321 out.n7313 0.063
R75952 out.n6323 out.n6322 0.063
R75953 out.n2534 out.n2533 0.063
R75954 out.n2035 out.n2034 0.063
R75955 out.n2911 out.n2910 0.063
R75956 out.n1815 out.n1814 0.063
R75957 out.n5502 out.n5501 0.063
R75958 out.n7360 out.n7359 0.063
R75959 out.n7142 out.n7141 0.062
R75960 out.n13192 out.n13190 0.062
R75961 out.n12675 out.n12425 0.062
R75962 out.n12625 out.n12623 0.062
R75963 out.n12327 out.n12325 0.062
R75964 out.n12327 out.n12326 0.062
R75965 out.n12232 out.n12231 0.062
R75966 out.n13508 out.n13269 0.062
R75967 out.n13458 out.n13456 0.062
R75968 out.n11496 out.n11494 0.062
R75969 out.n11069 out.n11067 0.062
R75970 out.n11907 out.n11905 0.062
R75971 out.n13963 out.n13724 0.062
R75972 out.n13913 out.n13911 0.062
R75973 out.n10640 out.n10638 0.062
R75974 out.n14472 out.n14303 0.062
R75975 out.n14174 out.n14171 0.062
R75976 out.n5146 out.n4990 0.062
R75977 out.n1050 out.n1032 0.062
R75978 out.n5804 out.n5802 0.062
R75979 out.n6376 out.n6374 0.062
R75980 out.n6938 out.n6936 0.062
R75981 out.n7759 out.n7757 0.062
R75982 out.n2704 out.n2703 0.062
R75983 out.n12546 out.n12446 0.062
R75984 out.n11285 out.n11184 0.062
R75985 out.n5717 out.n5654 0.062
R75986 out.n5473 out.n5419 0.062
R75987 out.n6851 out.n6788 0.062
R75988 out.n7331 out.n7280 0.062
R75989 out.n7603 out.n7602 0.062
R75990 out.n10855 out.n10758 0.061
R75991 out.n6294 out.n6231 0.061
R75992 out.n6543 out.n6530 0.061
R75993 out.n5972 out.n5971 0.061
R75994 out.n12132 out.n12131 0.061
R75995 out.n12108 out.n12016 0.061
R75996 out.n13379 out.n13290 0.061
R75997 out.n13834 out.n13745 0.061
R75998 out.n7113 out.n7052 0.061
R75999 out.n2552 out.n2436 0.061
R76000 out.n12973 out.n12883 0.061
R76001 out.n11688 out.n11598 0.061
R76002 out.n10421 out.n10331 0.061
R76003 out.n6637 out.n6488 0.061
R76004 out.n6076 out.n5900 0.061
R76005 out.n2666 out.n2653 0.061
R76006 out.n2129 out.n2104 0.061
R76007 out.n1570 out.n1563 0.061
R76008 out.n7697 out.n7524 0.061
R76009 out.n6092 out.n6091 0.061
R76010 out.n965 out.n964 0.061
R76011 out.n1183 out.n1182 0.061
R76012 out.n1915 out.n1914 0.061
R76013 out.n12997 out.n12996 0.06
R76014 out.n11712 out.n11711 0.06
R76015 out.n10445 out.n10444 0.06
R76016 out.n2791 out.n2790 0.06
R76017 out.n1383 out.n1382 0.06
R76018 out.n1695 out.n1694 0.06
R76019 out.n2227 out.n2226 0.06
R76020 out.n5993 out.n5992 0.06
R76021 out.n13404 out.n13403 0.06
R76022 out.n13859 out.n13858 0.06
R76023 out.n13192 out.n13191 0.06
R76024 out.n13097 out.n13096 0.06
R76025 out.n13603 out.n13602 0.06
R76026 out.n13508 out.n13507 0.06
R76027 out.n11907 out.n11906 0.06
R76028 out.n11812 out.n11811 0.06
R76029 out.n14058 out.n14057 0.06
R76030 out.n13963 out.n13962 0.06
R76031 out.n10640 out.n10639 0.06
R76032 out.n10545 out.n10544 0.06
R76033 out.n11418 out.n11417 0.059
R76034 out.n11313 out.n11312 0.059
R76035 out.n10991 out.n10990 0.059
R76036 out.n10886 out.n10885 0.059
R76037 out.n12249 out.n12248 0.059
R76038 out.n12139 out.n12138 0.059
R76039 out.n13097 out.n13086 0.059
R76040 out.n12758 out.n12757 0.059
R76041 out.n12747 out.n12746 0.059
R76042 out.n12736 out.n12735 0.059
R76043 out.n12729 out.n12728 0.059
R76044 out.n12647 out.n12646 0.059
R76045 out.n12636 out.n12635 0.059
R76046 out.n12625 out.n12624 0.059
R76047 out.n12616 out.n12615 0.059
R76048 out.n12527 out.n12526 0.059
R76049 out.n12516 out.n12515 0.059
R76050 out.n12507 out.n12506 0.059
R76051 out.n12498 out.n12497 0.059
R76052 out.n11483 out.n11482 0.059
R76053 out.n11472 out.n11471 0.059
R76054 out.n11461 out.n11460 0.059
R76055 out.n11452 out.n11451 0.059
R76056 out.n11378 out.n11377 0.059
R76057 out.n11367 out.n11366 0.059
R76058 out.n11358 out.n11357 0.059
R76059 out.n11349 out.n11348 0.059
R76060 out.n11266 out.n11265 0.059
R76061 out.n11254 out.n11253 0.059
R76062 out.n11243 out.n11242 0.059
R76063 out.n11234 out.n11233 0.059
R76064 out.n11220 out.n11219 0.059
R76065 out.n11812 out.n11801 0.059
R76066 out.n10545 out.n10534 0.059
R76067 out.n5685 out.n5684 0.059
R76068 out.n5673 out.n5672 0.059
R76069 out.n5664 out.n5663 0.059
R76070 out.n2889 out.n2888 0.059
R76071 out.n5815 out.n5814 0.059
R76072 out.n5804 out.n5803 0.059
R76073 out.n5795 out.n5794 0.059
R76074 out.n5786 out.n5785 0.059
R76075 out.n5569 out.n5568 0.059
R76076 out.n5558 out.n5557 0.059
R76077 out.n5549 out.n5548 0.059
R76078 out.n5540 out.n5539 0.059
R76079 out.n6819 out.n6818 0.059
R76080 out.n6807 out.n6806 0.059
R76081 out.n6798 out.n6797 0.059
R76082 out.n1793 out.n1792 0.059
R76083 out.n6949 out.n6948 0.059
R76084 out.n6938 out.n6937 0.059
R76085 out.n6929 out.n6928 0.059
R76086 out.n6920 out.n6919 0.059
R76087 out.n7427 out.n7426 0.059
R76088 out.n7416 out.n7415 0.059
R76089 out.n7407 out.n7406 0.059
R76090 out.n7398 out.n7397 0.059
R76091 out.n6666 out.n6665 0.059
R76092 out.n2581 out.n2580 0.059
R76093 out.n13114 out.n13113 0.059
R76094 out.n13004 out.n13003 0.059
R76095 out.n11829 out.n11828 0.059
R76096 out.n11719 out.n11718 0.059
R76097 out.n10562 out.n10561 0.059
R76098 out.n10452 out.n10451 0.059
R76099 out.n6101 out.n6100 0.059
R76100 out.n12818 out.n12817 0.058
R76101 out.n11550 out.n11549 0.058
R76102 out.n2892 out.n2891 0.058
R76103 out.n1796 out.n1795 0.058
R76104 out.n14270 out.n14269 0.058
R76105 out.n14339 out.n14338 0.058
R76106 out.n5026 out.n5025 0.058
R76107 out.n1322 out.n1321 0.058
R76108 out.n13097 out.n12862 0.058
R76109 out.n13193 out.n13192 0.058
R76110 out.n13049 out.n13047 0.058
R76111 out.n12769 out.n12767 0.058
R76112 out.n12767 out.n12764 0.058
R76113 out.n12791 out.n12790 0.058
R76114 out.n12609 out.n12608 0.058
R76115 out.n12491 out.n12490 0.058
R76116 out.n12484 out.n12483 0.058
R76117 out.n12232 out.n11995 0.058
R76118 out.n12232 out.n12221 0.058
R76119 out.n12184 out.n12182 0.058
R76120 out.n13603 out.n13601 0.058
R76121 out.n13601 out.n13598 0.058
R76122 out.n13604 out.n13603 0.058
R76123 out.n11406 out.n11160 0.058
R76124 out.n11518 out.n11517 0.058
R76125 out.n11358 out.n11356 0.058
R76126 out.n11342 out.n11341 0.058
R76127 out.n11227 out.n11226 0.058
R76128 out.n10979 out.n10737 0.058
R76129 out.n10931 out.n10929 0.058
R76130 out.n11812 out.n11577 0.058
R76131 out.n11908 out.n11907 0.058
R76132 out.n11764 out.n11762 0.058
R76133 out.n14058 out.n14056 0.058
R76134 out.n14056 out.n14053 0.058
R76135 out.n14059 out.n14058 0.058
R76136 out.n10545 out.n10310 0.058
R76137 out.n10641 out.n10640 0.058
R76138 out.n10497 out.n10495 0.058
R76139 out.n14430 out.n14345 0.058
R76140 out.n14411 out.n14393 0.058
R76141 out.n5104 out.n5033 0.058
R76142 out.n5085 out.n5082 0.058
R76143 out.n2904 out.n2903 0.058
R76144 out.n2909 out.n2816 0.058
R76145 out.n5329 out.n5327 0.058
R76146 out.n5221 out.n5219 0.058
R76147 out.n6141 out.n6139 0.058
R76148 out.n1808 out.n1807 0.058
R76149 out.n1813 out.n1720 0.058
R76150 out.n7188 out.n7186 0.058
R76151 out.n2162 out.n2161 0.058
R76152 out.n2058 out.n2057 0.058
R76153 out.n2929 out.n2928 0.057
R76154 out.n1833 out.n1832 0.057
R76155 out.n2688 out.n2687 0.057
R76156 out.n11056 out.n11055 0.057
R76157 out.n11045 out.n11044 0.057
R76158 out.n11034 out.n11033 0.057
R76159 out.n11025 out.n11024 0.057
R76160 out.n10951 out.n10950 0.057
R76161 out.n10940 out.n10939 0.057
R76162 out.n10931 out.n10930 0.057
R76163 out.n10922 out.n10921 0.057
R76164 out.n10836 out.n10835 0.057
R76165 out.n10824 out.n10823 0.057
R76166 out.n10813 out.n10812 0.057
R76167 out.n10804 out.n10803 0.057
R76168 out.n10797 out.n10796 0.057
R76169 out.n10790 out.n10789 0.057
R76170 out.n5772 out.n5771 0.057
R76171 out.n5232 out.n5231 0.057
R76172 out.n5221 out.n5220 0.057
R76173 out.n5212 out.n5211 0.057
R76174 out.n1250 out.n1249 0.057
R76175 out.n1253 out.n1252 0.057
R76176 out.n1256 out.n1255 0.057
R76177 out.n1268 out.n1267 0.057
R76178 out.n5349 out.n5348 0.057
R76179 out.n5338 out.n5337 0.057
R76180 out.n5329 out.n5328 0.057
R76181 out.n5320 out.n5319 0.057
R76182 out.n6262 out.n6261 0.057
R76183 out.n6250 out.n6249 0.057
R76184 out.n6241 out.n6240 0.057
R76185 out.n2013 out.n2012 0.057
R76186 out.n2028 out.n2027 0.057
R76187 out.n6387 out.n6386 0.057
R76188 out.n6376 out.n6375 0.057
R76189 out.n6367 out.n6366 0.057
R76190 out.n6358 out.n6357 0.057
R76191 out.n6906 out.n6905 0.057
R76192 out.n2016 out.n2015 0.057
R76193 out.n7706 out.n7705 0.057
R76194 out.n7624 out.n7623 0.056
R76195 out.n11127 out.n11126 0.056
R76196 out.n1606 out.n1605 0.056
R76197 out.n12328 out.n12327 0.056
R76198 out.n12314 out.n12313 0.056
R76199 out.n12303 out.n12302 0.056
R76200 out.n12292 out.n12291 0.056
R76201 out.n12283 out.n12282 0.056
R76202 out.n12204 out.n12203 0.056
R76203 out.n12193 out.n12192 0.056
R76204 out.n12184 out.n12183 0.056
R76205 out.n12175 out.n12174 0.056
R76206 out.n12089 out.n12088 0.056
R76207 out.n12077 out.n12076 0.056
R76208 out.n12066 out.n12065 0.056
R76209 out.n12057 out.n12056 0.056
R76210 out.n12043 out.n12042 0.056
R76211 out.n13508 out.n13500 0.056
R76212 out.n13592 out.n13591 0.056
R76213 out.n13581 out.n13580 0.056
R76214 out.n13570 out.n13569 0.056
R76215 out.n13563 out.n13562 0.056
R76216 out.n13480 out.n13479 0.056
R76217 out.n13469 out.n13468 0.056
R76218 out.n13458 out.n13457 0.056
R76219 out.n13449 out.n13448 0.056
R76220 out.n13360 out.n13359 0.056
R76221 out.n13349 out.n13348 0.056
R76222 out.n13340 out.n13339 0.056
R76223 out.n13331 out.n13330 0.056
R76224 out.n13317 out.n13316 0.056
R76225 out.n10979 out.n10968 0.056
R76226 out.n11091 out.n11090 0.056
R76227 out.n10915 out.n10914 0.056
R76228 out.n13963 out.n13955 0.056
R76229 out.n14047 out.n14046 0.056
R76230 out.n14036 out.n14035 0.056
R76231 out.n14025 out.n14024 0.056
R76232 out.n14018 out.n14017 0.056
R76233 out.n13935 out.n13934 0.056
R76234 out.n13924 out.n13923 0.056
R76235 out.n13913 out.n13912 0.056
R76236 out.n13904 out.n13903 0.056
R76237 out.n13815 out.n13814 0.056
R76238 out.n13804 out.n13803 0.056
R76239 out.n13795 out.n13794 0.056
R76240 out.n13786 out.n13785 0.056
R76241 out.n13772 out.n13771 0.056
R76242 out.n14472 out.n14471 0.056
R76243 out.n14430 out.n14429 0.056
R76244 out.n15905 out.n15375 0.056
R76245 out.n5146 out.n5145 0.056
R76246 out.n5104 out.n5103 0.056
R76247 out.n1265 out.n1264 0.056
R76248 out.n5276 out.n5265 0.056
R76249 out.n6445 out.n6438 0.056
R76250 out.n2033 out.n1940 0.056
R76251 out.n6349 out.n6348 0.056
R76252 out.n7008 out.n7003 0.056
R76253 out.n7081 out.n7080 0.056
R76254 out.n7071 out.n7070 0.056
R76255 out.n7062 out.n7061 0.056
R76256 out.n2528 out.n2527 0.056
R76257 out.n7199 out.n7198 0.056
R76258 out.n7188 out.n7187 0.056
R76259 out.n7179 out.n7178 0.056
R76260 out.n7248 out.n7243 0.056
R76261 out.n9439 out.n9433 0.056
R76262 out.n9458 out.n9457 0.056
R76263 out.n6573 out.n6572 0.056
R76264 out.n1483 out.n1482 0.055
R76265 out.n2330 out.n2329 0.055
R76266 out.n14522 out.n14521 0.055
R76267 out.n1056 out.n1055 0.055
R76268 out.n14523 out.n14522 0.055
R76269 out.n1055 out.n1054 0.055
R76270 out.n12388 out.n12387 0.055
R76271 out.n5492 out.n5491 0.055
R76272 out.n7350 out.n7349 0.055
R76273 out.n13665 out.n13664 0.055
R76274 out.n13698 out.n13697 0.055
R76275 out.n12770 out.n12769 0.055
R76276 out.n12721 out.n12720 0.055
R76277 out.n12715 out.n12714 0.055
R76278 out.n12666 out.n12665 0.055
R76279 out.n12561 out.n12560 0.055
R76280 out.n12548 out.n12547 0.055
R76281 out.n12545 out.n12544 0.055
R76282 out.n12507 out.n12505 0.055
R76283 out.n12349 out.n12348 0.055
R76284 out.n12168 out.n12167 0.055
R76285 out.n12050 out.n12049 0.055
R76286 out.n13625 out.n13624 0.055
R76287 out.n13442 out.n13441 0.055
R76288 out.n13340 out.n13338 0.055
R76289 out.n13324 out.n13323 0.055
R76290 out.n11406 out.n11395 0.055
R76291 out.n11444 out.n11443 0.055
R76292 out.n11438 out.n11437 0.055
R76293 out.n11394 out.n11393 0.055
R76294 out.n11298 out.n11297 0.055
R76295 out.n11287 out.n11286 0.055
R76296 out.n11284 out.n11283 0.055
R76297 out.n11070 out.n11069 0.055
R76298 out.n14080 out.n14079 0.055
R76299 out.n13897 out.n13896 0.055
R76300 out.n13795 out.n13793 0.055
R76301 out.n13779 out.n13778 0.055
R76302 out.n14473 out.n14472 0.055
R76303 out.n14431 out.n14430 0.055
R76304 out.n5147 out.n5146 0.055
R76305 out.n5105 out.n5104 0.055
R76306 out.n5795 out.n5793 0.055
R76307 out.n5673 out.n5671 0.055
R76308 out.n2886 out.n2885 0.055
R76309 out.n2901 out.n2900 0.055
R76310 out.n5743 out.n5742 0.055
R76311 out.n5730 out.n5729 0.055
R76312 out.n5719 out.n5718 0.055
R76313 out.n5853 out.n5852 0.055
R76314 out.n5842 out.n5841 0.055
R76315 out.n2923 out.n2763 0.055
R76316 out.n2925 out.n2756 0.055
R76317 out.n1474 out.n1454 0.055
R76318 out.n5549 out.n5547 0.055
R76319 out.n5489 out.n5488 0.055
R76320 out.n5478 out.n5477 0.055
R76321 out.n5475 out.n5474 0.055
R76322 out.n1511 out.n1364 0.055
R76323 out.n1253 out.n1236 0.055
R76324 out.n6703 out.n6701 0.055
R76325 out.n6367 out.n6365 0.055
R76326 out.n6250 out.n6248 0.055
R76327 out.n6929 out.n6927 0.055
R76328 out.n6807 out.n6805 0.055
R76329 out.n1790 out.n1789 0.055
R76330 out.n1805 out.n1804 0.055
R76331 out.n6877 out.n6876 0.055
R76332 out.n6864 out.n6863 0.055
R76333 out.n6853 out.n6852 0.055
R76334 out.n6987 out.n6986 0.055
R76335 out.n6976 out.n6975 0.055
R76336 out.n1827 out.n1667 0.055
R76337 out.n1829 out.n1660 0.055
R76338 out.n2321 out.n2298 0.055
R76339 out.n7407 out.n7405 0.055
R76340 out.n7347 out.n7346 0.055
R76341 out.n7336 out.n7335 0.055
R76342 out.n7333 out.n7332 0.055
R76343 out.n2358 out.n2208 0.055
R76344 out.n2543 out.n2542 0.055
R76345 out.n2547 out.n2463 0.055
R76346 out.n7750 out.n7748 0.055
R76347 out.n7654 out.n7652 0.055
R76348 out.n1514 out.n1513 0.055
R76349 out.n2361 out.n2360 0.055
R76350 out.n2531 out.n2530 0.055
R76351 out.n5590 out.n5396 0.054
R76352 out.n7448 out.n7257 0.054
R76353 out.n6744 out.n6455 0.054
R76354 out.n6180 out.n5878 0.054
R76355 out.n7795 out.n7484 0.054
R76356 out.n13214 out.n13213 0.054
R76357 out.n13179 out.n13178 0.054
R76358 out.n13168 out.n13167 0.054
R76359 out.n13157 out.n13156 0.054
R76360 out.n13148 out.n13147 0.054
R76361 out.n13069 out.n13068 0.054
R76362 out.n13058 out.n13057 0.054
R76363 out.n13049 out.n13048 0.054
R76364 out.n13040 out.n13039 0.054
R76365 out.n13033 out.n13032 0.054
R76366 out.n12954 out.n12953 0.054
R76367 out.n12942 out.n12941 0.054
R76368 out.n12931 out.n12930 0.054
R76369 out.n12922 out.n12921 0.054
R76370 out.n12915 out.n12914 0.054
R76371 out.n12908 out.n12907 0.054
R76372 out.n12846 out.n12845 0.054
R76373 out.n12675 out.n12667 0.054
R76374 out.n11497 out.n11496 0.054
R76375 out.n11017 out.n11016 0.054
R76376 out.n10967 out.n10966 0.054
R76377 out.n10868 out.n10867 0.054
R76378 out.n10857 out.n10856 0.054
R76379 out.n10854 out.n10853 0.054
R76380 out.n11929 out.n11928 0.054
R76381 out.n11894 out.n11893 0.054
R76382 out.n11883 out.n11882 0.054
R76383 out.n11872 out.n11871 0.054
R76384 out.n11863 out.n11862 0.054
R76385 out.n11784 out.n11783 0.054
R76386 out.n11773 out.n11772 0.054
R76387 out.n11764 out.n11763 0.054
R76388 out.n11755 out.n11754 0.054
R76389 out.n11748 out.n11747 0.054
R76390 out.n11669 out.n11668 0.054
R76391 out.n11657 out.n11656 0.054
R76392 out.n11646 out.n11645 0.054
R76393 out.n11637 out.n11636 0.054
R76394 out.n11630 out.n11629 0.054
R76395 out.n11623 out.n11622 0.054
R76396 out.n11967 out.n11966 0.054
R76397 out.n10662 out.n10661 0.054
R76398 out.n10627 out.n10626 0.054
R76399 out.n10616 out.n10615 0.054
R76400 out.n10605 out.n10604 0.054
R76401 out.n10596 out.n10595 0.054
R76402 out.n10517 out.n10516 0.054
R76403 out.n10506 out.n10505 0.054
R76404 out.n10497 out.n10496 0.054
R76405 out.n10488 out.n10487 0.054
R76406 out.n10481 out.n10480 0.054
R76407 out.n10402 out.n10401 0.054
R76408 out.n10390 out.n10389 0.054
R76409 out.n10379 out.n10378 0.054
R76410 out.n10370 out.n10369 0.054
R76411 out.n10363 out.n10362 0.054
R76412 out.n10356 out.n10355 0.054
R76413 out.n10700 out.n10699 0.054
R76414 out.n5264 out.n5263 0.054
R76415 out.n5253 out.n5252 0.054
R76416 out.n1315 out.n1164 0.054
R76417 out.n6723 out.n6722 0.054
R76418 out.n6712 out.n6711 0.054
R76419 out.n6703 out.n6702 0.054
R76420 out.n6694 out.n6693 0.054
R76421 out.n2010 out.n2009 0.054
R76422 out.n2025 out.n2024 0.054
R76423 out.n6320 out.n6319 0.054
R76424 out.n6307 out.n6306 0.054
R76425 out.n6296 out.n6295 0.054
R76426 out.n6425 out.n6424 0.054
R76427 out.n6414 out.n6413 0.054
R76428 out.n2052 out.n1892 0.054
R76429 out.n2054 out.n1885 0.054
R76430 out.n6051 out.n6050 0.054
R76431 out.n6039 out.n6038 0.054
R76432 out.n6028 out.n6027 0.054
R76433 out.n6019 out.n6018 0.054
R76434 out.n6161 out.n6160 0.054
R76435 out.n6150 out.n6149 0.054
R76436 out.n6141 out.n6140 0.054
R76437 out.n6132 out.n6131 0.054
R76438 out.n2540 out.n2539 0.054
R76439 out.n7636 out.n7526 0.054
R76440 out.n7634 out.n7531 0.054
R76441 out.n7734 out.n7487 0.054
R76442 out.n12849 out.n12848 0.054
R76443 out.n11970 out.n11969 0.054
R76444 out.n10703 out.n10702 0.054
R76445 out.n1523 out.n1522 0.054
R76446 out.n2370 out.n2369 0.054
R76447 out.n12693 out.n12692 0.053
R76448 out.n12580 out.n12579 0.053
R76449 out.n9442 out.n9441 0.053
R76450 out.n12782 out.n12781 0.053
R76451 out.n12706 out.n12705 0.053
R76452 out.n12601 out.n12600 0.053
R76453 out.n12477 out.n12476 0.053
R76454 out.n12220 out.n12219 0.053
R76455 out.n12121 out.n12120 0.053
R76456 out.n12110 out.n12109 0.053
R76457 out.n12107 out.n12106 0.053
R76458 out.n13499 out.n13498 0.053
R76459 out.n13394 out.n13393 0.053
R76460 out.n13381 out.n13380 0.053
R76461 out.n13378 out.n13377 0.053
R76462 out.n11011 out.n11010 0.053
R76463 out.n13954 out.n13953 0.053
R76464 out.n13849 out.n13848 0.053
R76465 out.n13836 out.n13835 0.053
R76466 out.n13833 out.n13832 0.053
R76467 out.n5519 out.n5518 0.053
R76468 out.n5313 out.n5312 0.053
R76469 out.n6619 out.n6490 0.053
R76470 out.n6617 out.n6616 0.053
R76471 out.n6605 out.n6604 0.053
R76472 out.n6596 out.n6595 0.053
R76473 out.n6589 out.n6588 0.053
R76474 out.n6582 out.n6581 0.053
R76475 out.n6687 out.n6459 0.053
R76476 out.n6685 out.n6464 0.053
R76477 out.n6012 out.n5905 0.053
R76478 out.n6010 out.n5910 0.053
R76479 out.n6125 out.n5882 0.053
R76480 out.n5949 out.n5948 0.053
R76481 out.n7377 out.n7376 0.053
R76482 out.n2525 out.n2524 0.053
R76483 out.n7139 out.n7138 0.053
R76484 out.n7126 out.n7125 0.053
R76485 out.n7115 out.n7114 0.053
R76486 out.n7233 out.n7232 0.053
R76487 out.n7222 out.n7221 0.053
R76488 out.n2573 out.n2420 0.053
R76489 out.n2575 out.n2413 0.053
R76490 out.n7632 out.n7536 0.053
R76491 out.n7666 out.n7665 0.053
R76492 out.n7654 out.n7653 0.053
R76493 out.n7645 out.n7644 0.053
R76494 out.n7770 out.n7769 0.053
R76495 out.n7759 out.n7758 0.053
R76496 out.n7750 out.n7749 0.053
R76497 out.n7741 out.n7740 0.053
R76498 out.n13527 out.n13526 0.053
R76499 out.n13413 out.n13412 0.053
R76500 out.n13982 out.n13981 0.053
R76501 out.n13868 out.n13867 0.053
R76502 out.n10108 out.n10107 0.052
R76503 out.n12684 out.n12683 0.052
R76504 out.n12593 out.n12592 0.052
R76505 out.n12471 out.n12470 0.052
R76506 out.n12275 out.n12274 0.052
R76507 out.n12269 out.n12268 0.052
R76508 out.n13555 out.n13554 0.052
R76509 out.n13549 out.n13548 0.052
R76510 out.n11509 out.n11508 0.052
R76511 out.n11420 out.n11419 0.052
R76512 out.n11414 out.n11413 0.052
R76513 out.n11334 out.n11333 0.052
R76514 out.n11315 out.n11314 0.052
R76515 out.n11213 out.n11212 0.052
R76516 out.n14010 out.n14009 0.052
R76517 out.n14004 out.n14003 0.052
R76518 out.n15906 out.n15374 0.052
R76519 out.n15159 out.n10044 0.052
R76520 out.n1058 out.n1002 0.052
R76521 out.n2898 out.n2897 0.052
R76522 out.n5766 out.n5765 0.052
R76523 out.n5757 out.n5756 0.052
R76524 out.n2931 out.n2739 0.052
R76525 out.n1485 out.n1434 0.052
R76526 out.n5513 out.n5512 0.052
R76527 out.n6443 out.n6440 0.052
R76528 out.n7007 out.n7006 0.052
R76529 out.n1802 out.n1801 0.052
R76530 out.n6900 out.n6899 0.052
R76531 out.n6891 out.n6890 0.052
R76532 out.n1835 out.n1643 0.052
R76533 out.n2332 out.n2278 0.052
R76534 out.n7371 out.n7370 0.052
R76535 out.n2545 out.n2470 0.052
R76536 out.n7168 out.n7035 0.052
R76537 out.n7104 out.n7103 0.052
R76538 out.n7166 out.n7165 0.052
R76539 out.n2550 out.n2549 0.052
R76540 out.n7247 out.n7246 0.052
R76541 out.n2123 out.n2122 0.052
R76542 out.n2159 out.n2158 0.052
R76543 out.n9436 out.t1 0.051
R76544 out.n5990 out.n5989 0.051
R76545 out.n6656 out.n6655 0.051
R76546 out.n1603 out.n1602 0.051
R76547 out.n13187 out.n13186 0.051
R76548 out.n13140 out.n13139 0.051
R76549 out.n13134 out.n13133 0.051
R76550 out.n13085 out.n13084 0.051
R76551 out.n12986 out.n12985 0.051
R76552 out.n12975 out.n12974 0.051
R76553 out.n12972 out.n12971 0.051
R76554 out.n12931 out.n12929 0.051
R76555 out.n12695 out.n12694 0.051
R76556 out.n12582 out.n12581 0.051
R76557 out.n12322 out.n12321 0.051
R76558 out.n12066 out.n12064 0.051
R76559 out.n13511 out.n13509 0.051
R76560 out.n13616 out.n13615 0.051
R76561 out.n13540 out.n13539 0.051
R76562 out.n11491 out.n11490 0.051
R76563 out.n11431 out.n11430 0.051
R76564 out.n11326 out.n11325 0.051
R76565 out.n11243 out.n11241 0.051
R76566 out.n11207 out.n11206 0.051
R76567 out.n11064 out.n11063 0.051
R76568 out.n11082 out.n11081 0.051
R76569 out.n11004 out.n11003 0.051
R76570 out.n10987 out.n10986 0.051
R76571 out.n10899 out.n10898 0.051
R76572 out.n10813 out.n10811 0.051
R76573 out.n10777 out.n10776 0.051
R76574 out.n11902 out.n11901 0.051
R76575 out.n11855 out.n11854 0.051
R76576 out.n11849 out.n11848 0.051
R76577 out.n11800 out.n11799 0.051
R76578 out.n11701 out.n11700 0.051
R76579 out.n11690 out.n11689 0.051
R76580 out.n11687 out.n11686 0.051
R76581 out.n11646 out.n11644 0.051
R76582 out.n13966 out.n13964 0.051
R76583 out.n14071 out.n14070 0.051
R76584 out.n13995 out.n13994 0.051
R76585 out.n10635 out.n10634 0.051
R76586 out.n10588 out.n10587 0.051
R76587 out.n10582 out.n10581 0.051
R76588 out.n10533 out.n10532 0.051
R76589 out.n10434 out.n10433 0.051
R76590 out.n10423 out.n10422 0.051
R76591 out.n10420 out.n10419 0.051
R76592 out.n10379 out.n10377 0.051
R76593 out.n14521 out.n14520 0.051
R76594 out.n14519 out.n14518 0.051
R76595 out.n14517 out.n14516 0.051
R76596 out.n14497 out.n14496 0.051
R76597 out.n14495 out.n14494 0.051
R76598 out.n14493 out.n14492 0.051
R76599 out.n14300 out.n14299 0.051
R76600 out.n14474 out.n14283 0.051
R76601 out.n14470 out.n14469 0.051
R76602 out.n14468 out.n14467 0.051
R76603 out.n14466 out.n14465 0.051
R76604 out.n14457 out.n14456 0.051
R76605 out.n14435 out.n14434 0.051
R76606 out.n14433 out.n14432 0.051
R76607 out.n14415 out.n14414 0.051
R76608 out.n14413 out.n14412 0.051
R76609 out.n14411 out.n14410 0.051
R76610 out.n14409 out.n14408 0.051
R76611 out.n14174 out.n14173 0.051
R76612 out.n14176 out.n14175 0.051
R76613 out.n4987 out.n4986 0.051
R76614 out.n5148 out.n4969 0.051
R76615 out.n5144 out.n5143 0.051
R76616 out.n5142 out.n5141 0.051
R76617 out.n5140 out.n5139 0.051
R76618 out.n5131 out.n5130 0.051
R76619 out.n5109 out.n5108 0.051
R76620 out.n5107 out.n5106 0.051
R76621 out.n5089 out.n5088 0.051
R76622 out.n5087 out.n5086 0.051
R76623 out.n5085 out.n5084 0.051
R76624 out.n1050 out.n1049 0.051
R76625 out.n1052 out.n1051 0.051
R76626 out.n1054 out.n1053 0.051
R76627 out.n1079 out.n1078 0.051
R76628 out.n1081 out.n1080 0.051
R76629 out.n1083 out.n1082 0.051
R76630 out.n1104 out.n1103 0.051
R76631 out.n1525 out.n1347 0.051
R76632 out.n5280 out.n5279 0.051
R76633 out.n5212 out.n5210 0.051
R76634 out.n1262 out.n1261 0.051
R76635 out.n5306 out.n5305 0.051
R76636 out.n1294 out.n1293 0.051
R76637 out.n1296 out.n1295 0.051
R76638 out.n1298 out.n1297 0.051
R76639 out.n1317 out.n1316 0.051
R76640 out.n6557 out.n6511 0.051
R76641 out.n6653 out.n6652 0.051
R76642 out.n6642 out.n6641 0.051
R76643 out.n6639 out.n6638 0.051
R76644 out.n2150 out.n2098 0.051
R76645 out.n6351 out.n6214 0.051
R76646 out.n2036 out.n2035 0.051
R76647 out.n2038 out.n2037 0.051
R76648 out.n2040 out.n2039 0.051
R76649 out.n6028 out.n6026 0.051
R76650 out.n5987 out.n5986 0.051
R76651 out.n5976 out.n5975 0.051
R76652 out.n6089 out.n6088 0.051
R76653 out.n6078 out.n6077 0.051
R76654 out.n1592 out.n1551 0.051
R76655 out.n2372 out.n2191 0.051
R76656 out.n7179 out.n7177 0.051
R76657 out.n7071 out.n7069 0.051
R76658 out.n7170 out.n7030 0.051
R76659 out.n7611 out.n7550 0.051
R76660 out.n7609 out.n7561 0.051
R76661 out.n7604 out.n7576 0.051
R76662 out.n7632 out.n7631 0.051
R76663 out.n7703 out.n7499 0.051
R76664 out.n7701 out.n7510 0.051
R76665 out.n7696 out.n7525 0.051
R76666 out.n7732 out.n7731 0.051
R76667 out.n2668 out.n2667 0.051
R76668 out.n2671 out.n2670 0.051
R76669 out.n2678 out.n2677 0.051
R76670 out.n2691 out.n2690 0.051
R76671 out.n2153 out.n2152 0.051
R76672 out.n1113 out.n1112 0.051
R76673 out.n9431 out.n9426 0.051
R76674 out.n5476 out.n5413 0.05
R76675 out.n7334 out.n7274 0.05
R76676 out.n2138 out.n2137 0.05
R76677 out.n1573 out.n1558 0.05
R76678 out.n12986 out.n12976 0.05
R76679 out.n13434 out.n13433 0.05
R76680 out.n13426 out.n13425 0.05
R76681 out.n13310 out.n13309 0.05
R76682 out.n13304 out.n13303 0.05
R76683 out.n10993 out.n10992 0.05
R76684 out.n10907 out.n10906 0.05
R76685 out.n10888 out.n10887 0.05
R76686 out.n10783 out.n10782 0.05
R76687 out.n11701 out.n11691 0.05
R76688 out.n13889 out.n13888 0.05
R76689 out.n13881 out.n13880 0.05
R76690 out.n13765 out.n13764 0.05
R76691 out.n13759 out.n13758 0.05
R76692 out.n10434 out.n10424 0.05
R76693 out.n14525 out.n14205 0.05
R76694 out.n14529 out.n14528 0.05
R76695 out.n14527 out.n14526 0.05
R76696 out.n14476 out.n14475 0.05
R76697 out.n14427 out.n14426 0.05
R76698 out.n14402 out.n14401 0.05
R76699 out.n5150 out.n5149 0.05
R76700 out.n5101 out.n5100 0.05
R76701 out.n1060 out.n1059 0.05
R76702 out.n1062 out.n1061 0.05
R76703 out.n2912 out.n2911 0.05
R76704 out.n2914 out.n2913 0.05
R76705 out.n2916 out.n2915 0.05
R76706 out.n5454 out.n5445 0.05
R76707 out.n5444 out.n5443 0.05
R76708 out.n5442 out.n5441 0.05
R76709 out.n1493 out.n1492 0.05
R76710 out.n1501 out.n1500 0.05
R76711 out.n1503 out.n1502 0.05
R76712 out.n5203 out.n5197 0.05
R76713 out.n1270 out.n1269 0.05
R76714 out.n5297 out.n5296 0.05
R76715 out.n5286 out.n5285 0.05
R76716 out.n6574 out.n6573 0.05
R76717 out.n6557 out.n6556 0.05
R76718 out.n6555 out.n6554 0.05
R76719 out.n6548 out.n6547 0.05
R76720 out.n6545 out.n6544 0.05
R76721 out.n6542 out.n6541 0.05
R76722 out.n6653 out.n6643 0.05
R76723 out.n6636 out.n6489 0.05
R76724 out.n6683 out.n6682 0.05
R76725 out.n2128 out.n2127 0.05
R76726 out.n2131 out.n2130 0.05
R76727 out.n2140 out.n2139 0.05
R76728 out.n2150 out.n2149 0.05
R76729 out.n2006 out.n2005 0.05
R76730 out.n2031 out.n2029 0.05
R76731 out.n2022 out.n2021 0.05
R76732 out.n6285 out.n6284 0.05
R76733 out.n6343 out.n6342 0.05
R76734 out.n6334 out.n6333 0.05
R76735 out.n2060 out.n1868 0.05
R76736 out.n2042 out.n2041 0.05
R76737 out.n5987 out.n5977 0.05
R76738 out.n5973 out.n5936 0.05
R76739 out.n5965 out.n5937 0.05
R76740 out.n6089 out.n6079 0.05
R76741 out.n6075 out.n5901 0.05
R76742 out.n1572 out.n1571 0.05
R76743 out.n1575 out.n1574 0.05
R76744 out.n1582 out.n1581 0.05
R76745 out.n1592 out.n1591 0.05
R76746 out.n1816 out.n1815 0.05
R76747 out.n1818 out.n1817 0.05
R76748 out.n1820 out.n1819 0.05
R76749 out.n7312 out.n7303 0.05
R76750 out.n7302 out.n7301 0.05
R76751 out.n7300 out.n7299 0.05
R76752 out.n2340 out.n2339 0.05
R76753 out.n2348 out.n2347 0.05
R76754 out.n2350 out.n2349 0.05
R76755 out.n2540 out.n2538 0.05
R76756 out.n7116 out.n7115 0.05
R76757 out.n7631 out.n7630 0.05
R76758 out.n7611 out.n7610 0.05
R76759 out.n7609 out.n7608 0.05
R76760 out.n7608 out.n7607 0.05
R76761 out.n7607 out.n7606 0.05
R76762 out.n7596 out.n7595 0.05
R76763 out.n7703 out.n7702 0.05
R76764 out.n7701 out.n7700 0.05
R76765 out.n7700 out.n7699 0.05
R76766 out.n7699 out.n7698 0.05
R76767 out.n2691 out.n2689 0.05
R76768 out.n2665 out.n2664 0.05
R76769 out.n6640 out.n6482 0.05
R76770 out.n2669 out.n2645 0.05
R76771 out.n1320 out.n1319 0.05
R76772 out.n6546 out.n6524 0.05
R76773 out.n7605 out.n7575 0.05
R76774 out.n6560 out.n6559 0.05
R76775 out.n1110 out.n1109 0.05
R76776 out.n2555 out.n2428 0.05
R76777 out.n5974 out.n5935 0.05
R76778 out.n2578 out.n2577 0.05
R76779 out.n1376 out.n1375 0.05
R76780 out.n2220 out.n2219 0.05
R76781 out.n961 out.n960 0.05
R76782 out.n1906 out.n1905 0.05
R76783 out.n2782 out.n2781 0.049
R76784 out.n1178 out.n1177 0.049
R76785 out.n1686 out.n1685 0.049
R76786 out.n7614 out.n7613 0.049
R76787 out.n9460 out.n9459 0.049
R76788 out.n12340 out.n12339 0.049
R76789 out.n12262 out.n12261 0.049
R76790 out.n12251 out.n12250 0.049
R76791 out.n12240 out.n12239 0.049
R76792 out.n12121 out.n12111 0.049
R76793 out.n12160 out.n12159 0.049
R76794 out.n12152 out.n12151 0.049
R76795 out.n12141 out.n12140 0.049
R76796 out.n12036 out.n12035 0.049
R76797 out.n12030 out.n12029 0.049
R76798 out.n13529 out.n13528 0.049
R76799 out.n13518 out.n13517 0.049
R76800 out.n13394 out.n13382 0.049
R76801 out.n13415 out.n13414 0.049
R76802 out.n13984 out.n13983 0.049
R76803 out.n13973 out.n13972 0.049
R76804 out.n13849 out.n13837 0.049
R76805 out.n13870 out.n13869 0.049
R76806 out.n17312 out.n8879 0.049
R76807 out.n2882 out.n2881 0.049
R76808 out.n2907 out.n2905 0.049
R76809 out.n5779 out.n5773 0.049
R76810 out.n5708 out.n5707 0.049
R76811 out.n2918 out.n2917 0.049
R76812 out.n2920 out.n2919 0.049
R76813 out.n1469 out.n1468 0.049
R76814 out.n1471 out.n1470 0.049
R76815 out.n1487 out.n1486 0.049
R76816 out.n1489 out.n1488 0.049
R76817 out.n1491 out.n1490 0.049
R76818 out.n5533 out.n5527 0.049
R76819 out.n5526 out.n5520 0.049
R76820 out.n5464 out.n5463 0.049
R76821 out.n1505 out.n1504 0.049
R76822 out.n1507 out.n1506 0.049
R76823 out.n1265 out.n1263 0.049
R76824 out.n5254 out.n5253 0.049
R76825 out.n6575 out.n6498 0.049
R76826 out.n2008 out.n2007 0.049
R76827 out.n1786 out.n1785 0.049
R76828 out.n1811 out.n1809 0.049
R76829 out.n6913 out.n6907 0.049
R76830 out.n6842 out.n6841 0.049
R76831 out.n1822 out.n1821 0.049
R76832 out.n1824 out.n1823 0.049
R76833 out.n2316 out.n2315 0.049
R76834 out.n2318 out.n2317 0.049
R76835 out.n2334 out.n2333 0.049
R76836 out.n2336 out.n2335 0.049
R76837 out.n2338 out.n2337 0.049
R76838 out.n7391 out.n7385 0.049
R76839 out.n7384 out.n7378 0.049
R76840 out.n7322 out.n7321 0.049
R76841 out.n2352 out.n2351 0.049
R76842 out.n2354 out.n2353 0.049
R76843 out.n2515 out.n2514 0.049
R76844 out.n2522 out.n2521 0.049
R76845 out.n2525 out.n2523 0.049
R76846 out.n2535 out.n2534 0.049
R76847 out.n2538 out.n2537 0.049
R76848 out.n2537 out.n2536 0.049
R76849 out.n7139 out.n7127 0.049
R76850 out.n7126 out.n7116 0.049
R76851 out.n7112 out.n7104 0.049
R76852 out.n7160 out.n7159 0.049
R76853 out.n7151 out.n7150 0.049
R76854 out.n7233 out.n7223 0.049
R76855 out.n7223 out.n7222 0.049
R76856 out.n2583 out.n2397 0.049
R76857 out.n2554 out.n2553 0.049
R76858 out.n2564 out.n2563 0.049
R76859 out.n2571 out.n2570 0.049
R76860 out.n2573 out.n2572 0.049
R76861 out.n2575 out.n2574 0.049
R76862 out.n2582 out.n2581 0.049
R76863 out.n1520 out.n1519 0.049
R76864 out.n2367 out.n2366 0.049
R76865 out.n6568 out.n6567 0.049
R76866 out.n5295 out.n5294 0.049
R76867 out.n1479 out.n1478 0.048
R76868 out.n2326 out.n2325 0.048
R76869 out.n7149 out.n7148 0.048
R76870 out.n1481 out.n1480 0.048
R76871 out.n2328 out.n2327 0.048
R76872 out.n10142 out.n10139 0.048
R76873 out.n9453 out.n9452 0.048
R76874 out.n13086 out.n13085 0.048
R76875 out.n13205 out.n13204 0.048
R76876 out.n13116 out.n13115 0.048
R76877 out.n13105 out.n13104 0.048
R76878 out.n12976 out.n12975 0.048
R76879 out.n13006 out.n13005 0.048
R76880 out.n10868 out.n10858 0.048
R76881 out.n11801 out.n11800 0.048
R76882 out.n11920 out.n11919 0.048
R76883 out.n11831 out.n11830 0.048
R76884 out.n11820 out.n11819 0.048
R76885 out.n11691 out.n11690 0.048
R76886 out.n11721 out.n11720 0.048
R76887 out.n10534 out.n10533 0.048
R76888 out.n10653 out.n10652 0.048
R76889 out.n10564 out.n10563 0.048
R76890 out.n10553 out.n10552 0.048
R76891 out.n10424 out.n10423 0.048
R76892 out.n10454 out.n10453 0.048
R76893 out.n14528 out.n14527 0.048
R76894 out.n14526 out.n14525 0.048
R76895 out.n14524 out.n14523 0.048
R76896 out.n14508 out.n14507 0.048
R76897 out.n14505 out.n14504 0.048
R76898 out.n14496 out.n14495 0.048
R76899 out.n14475 out.n14474 0.048
R76900 out.n14428 out.n14427 0.048
R76901 out.n5149 out.n5148 0.048
R76902 out.n5102 out.n5101 0.048
R76903 out.n1039 out.n1038 0.048
R76904 out.n1046 out.n1045 0.048
R76905 out.n1057 out.n1056 0.048
R76906 out.n1059 out.n1058 0.048
R76907 out.n1061 out.n1060 0.048
R76908 out.n1094 out.n1093 0.048
R76909 out.n1101 out.n1100 0.048
R76910 out.n2922 out.n2921 0.048
R76911 out.n1247 out.n1246 0.048
R76912 out.n1260 out.n1259 0.048
R76913 out.n1263 out.n1262 0.048
R76914 out.n1269 out.n1268 0.048
R76915 out.n5264 out.n5254 0.048
R76916 out.n1299 out.n1298 0.048
R76917 out.n1306 out.n1305 0.048
R76918 out.n1313 out.n1312 0.048
R76919 out.n1315 out.n1314 0.048
R76920 out.n6575 out.n6574 0.048
R76921 out.n6677 out.n6676 0.048
R76922 out.n2149 out.n2148 0.048
R76923 out.n2005 out.n2004 0.048
R76924 out.n2007 out.n2006 0.048
R76925 out.n2010 out.n2008 0.048
R76926 out.n2020 out.n2019 0.048
R76927 out.n2023 out.n2022 0.048
R76928 out.n2029 out.n2028 0.048
R76929 out.n6320 out.n6308 0.048
R76930 out.n6307 out.n6297 0.048
R76931 out.n6293 out.n6285 0.048
R76932 out.n6425 out.n6415 0.048
R76933 out.n2041 out.n2040 0.048
R76934 out.n2043 out.n2042 0.048
R76935 out.n2050 out.n2049 0.048
R76936 out.n2051 out.n2050 0.048
R76937 out.n2052 out.n2051 0.048
R76938 out.n2054 out.n2053 0.048
R76939 out.n2059 out.n2058 0.048
R76940 out.n5977 out.n5976 0.048
R76941 out.n6079 out.n6078 0.048
R76942 out.n6103 out.n6102 0.048
R76943 out.n1826 out.n1825 0.048
R76944 out.n2523 out.n2522 0.048
R76945 out.n2551 out.n2550 0.048
R76946 out.n2557 out.n2556 0.048
R76947 out.n2572 out.n2571 0.048
R76948 out.n1500 out.n1499 0.048
R76949 out.n2347 out.n2346 0.048
R76950 out.n1134 out.n1130 0.048
R76951 out.n2057 out.n2056 0.048
R76952 out.n17312 out.n4 0.047
R76953 out.n6747 out.n6746 0.047
R76954 out.n5593 out.n5592 0.047
R76955 out.n7451 out.n7450 0.047
R76956 out.n13237 out.n13234 0.047
R76957 out.n13168 out.n13166 0.047
R76958 out.n13179 out.n13177 0.047
R76959 out.n13205 out.n13193 0.047
R76960 out.n13127 out.n13126 0.047
R76961 out.n13069 out.n13067 0.047
R76962 out.n13025 out.n13024 0.047
R76963 out.n13017 out.n13016 0.047
R76964 out.n12846 out.n12844 0.047
R76965 out.n12901 out.n12900 0.047
R76966 out.n12747 out.n12745 0.047
R76967 out.n12758 out.n12756 0.047
R76968 out.n12636 out.n12634 0.047
R76969 out.n12647 out.n12645 0.047
R76970 out.n12561 out.n12549 0.047
R76971 out.n12527 out.n12525 0.047
R76972 out.n12303 out.n12301 0.047
R76973 out.n12314 out.n12312 0.047
R76974 out.n12221 out.n12220 0.047
R76975 out.n12204 out.n12202 0.047
R76976 out.n12385 out.n12384 0.047
R76977 out.n13581 out.n13579 0.047
R76978 out.n13592 out.n13590 0.047
R76979 out.n13616 out.n13604 0.047
R76980 out.n13469 out.n13467 0.047
R76981 out.n13480 out.n13478 0.047
R76982 out.n13662 out.n13661 0.047
R76983 out.n13360 out.n13358 0.047
R76984 out.n11414 out.n11157 0.047
R76985 out.n11472 out.n11470 0.047
R76986 out.n11483 out.n11481 0.047
R76987 out.n11309 out.n11178 0.047
R76988 out.n11378 out.n11376 0.047
R76989 out.n11298 out.n11288 0.047
R76990 out.n10987 out.n10734 0.047
R76991 out.n11045 out.n11043 0.047
R76992 out.n11056 out.n11054 0.047
R76993 out.n10951 out.n10949 0.047
R76994 out.n11883 out.n11881 0.047
R76995 out.n11894 out.n11892 0.047
R76996 out.n11920 out.n11908 0.047
R76997 out.n11842 out.n11841 0.047
R76998 out.n11784 out.n11782 0.047
R76999 out.n11740 out.n11739 0.047
R77000 out.n11732 out.n11731 0.047
R77001 out.n11967 out.n11965 0.047
R77002 out.n11616 out.n11615 0.047
R77003 out.n14036 out.n14034 0.047
R77004 out.n14047 out.n14045 0.047
R77005 out.n14071 out.n14059 0.047
R77006 out.n13924 out.n13922 0.047
R77007 out.n13935 out.n13933 0.047
R77008 out.n13695 out.n13694 0.047
R77009 out.n13815 out.n13813 0.047
R77010 out.n10616 out.n10614 0.047
R77011 out.n10627 out.n10625 0.047
R77012 out.n10653 out.n10641 0.047
R77013 out.n10575 out.n10574 0.047
R77014 out.n10517 out.n10515 0.047
R77015 out.n10473 out.n10472 0.047
R77016 out.n10465 out.n10464 0.047
R77017 out.n10700 out.n10698 0.047
R77018 out.n10349 out.n10348 0.047
R77019 out.n14519 out.n14241 0.047
R77020 out.n14521 out.n14232 0.047
R77021 out.n14498 out.n14497 0.047
R77022 out.n14468 out.n14321 0.047
R77023 out.n14470 out.n14312 0.047
R77024 out.n14449 out.n14448 0.047
R77025 out.n14443 out.n14442 0.047
R77026 out.n14176 out.n14165 0.047
R77027 out.n14415 out.n14379 0.047
R77028 out.n14412 out.n14411 0.047
R77029 out.n14410 out.n14409 0.047
R77030 out.n5142 out.n5008 0.047
R77031 out.n5144 out.n4999 0.047
R77032 out.n5123 out.n5122 0.047
R77033 out.n5117 out.n5116 0.047
R77034 out.n1054 out.n1017 0.047
R77035 out.n1052 out.n1026 0.047
R77036 out.n5089 out.n5068 0.047
R77037 out.n5086 out.n5085 0.047
R77038 out.n5084 out.n5083 0.047
R77039 out.n1080 out.n1079 0.047
R77040 out.n1082 out.n1081 0.047
R77041 out.n1084 out.n1083 0.047
R77042 out.n1087 out.n1086 0.047
R77043 out.n5815 out.n5813 0.047
R77044 out.n5664 out.n5662 0.047
R77045 out.n2815 out.n2813 0.047
R77046 out.n2881 out.n2880 0.047
R77047 out.n2883 out.n2882 0.047
R77048 out.n2884 out.n2883 0.047
R77049 out.n2886 out.n2884 0.047
R77050 out.n2896 out.n2895 0.047
R77051 out.n2899 out.n2898 0.047
R77052 out.n2905 out.n2904 0.047
R77053 out.n5773 out.n5772 0.047
R77054 out.n5743 out.n5731 0.047
R77055 out.n5730 out.n5720 0.047
R77056 out.n5720 out.n5719 0.047
R77057 out.n5716 out.n5708 0.047
R77058 out.n5853 out.n5843 0.047
R77059 out.n2796 out.n2793 0.047
R77060 out.n2917 out.n2916 0.047
R77061 out.n2919 out.n2918 0.047
R77062 out.n2921 out.n2920 0.047
R77063 out.n2923 out.n2922 0.047
R77064 out.n2925 out.n2924 0.047
R77065 out.n2930 out.n2929 0.047
R77066 out.n5442 out.n5436 0.047
R77067 out.n5443 out.n5442 0.047
R77068 out.n1470 out.n1469 0.047
R77069 out.n1472 out.n1471 0.047
R77070 out.n1474 out.n1473 0.047
R77071 out.n1484 out.n1483 0.047
R77072 out.n1486 out.n1485 0.047
R77073 out.n1488 out.n1487 0.047
R77074 out.n1490 out.n1489 0.047
R77075 out.n5569 out.n5567 0.047
R77076 out.n5527 out.n5526 0.047
R77077 out.n5520 out.n5519 0.047
R77078 out.n5489 out.n5479 0.047
R77079 out.n5472 out.n5464 0.047
R77080 out.n1506 out.n1505 0.047
R77081 out.n1511 out.n1510 0.047
R77082 out.n5349 out.n5347 0.047
R77083 out.n1256 out.n1230 0.047
R77084 out.n1295 out.n1294 0.047
R77085 out.n1297 out.n1296 0.047
R77086 out.n1314 out.n1313 0.047
R77087 out.n6605 out.n6603 0.047
R77088 out.n6556 out.n6555 0.047
R77089 out.n6723 out.n6721 0.047
R77090 out.n6643 out.n6642 0.047
R77091 out.n2164 out.n2083 0.047
R77092 out.n2163 out.n2162 0.047
R77093 out.n2164 out.n2163 0.047
R77094 out.n6387 out.n6385 0.047
R77095 out.n6241 out.n6239 0.047
R77096 out.n1939 out.n1937 0.047
R77097 out.n2025 out.n2023 0.047
R77098 out.n6297 out.n6296 0.047
R77099 out.n6415 out.n6414 0.047
R77100 out.n1920 out.n1917 0.047
R77101 out.n2037 out.n2036 0.047
R77102 out.n2039 out.n2038 0.047
R77103 out.n6161 out.n6159 0.047
R77104 out.n6008 out.n6007 0.047
R77105 out.n6002 out.n6001 0.047
R77106 out.n6122 out.n6121 0.047
R77107 out.n6114 out.n6113 0.047
R77108 out.n1591 out.n1590 0.047
R77109 out.n6949 out.n6947 0.047
R77110 out.n6798 out.n6796 0.047
R77111 out.n1719 out.n1717 0.047
R77112 out.n1785 out.n1784 0.047
R77113 out.n1787 out.n1786 0.047
R77114 out.n1788 out.n1787 0.047
R77115 out.n1790 out.n1788 0.047
R77116 out.n1800 out.n1799 0.047
R77117 out.n1803 out.n1802 0.047
R77118 out.n1809 out.n1808 0.047
R77119 out.n6907 out.n6906 0.047
R77120 out.n6877 out.n6865 0.047
R77121 out.n6864 out.n6854 0.047
R77122 out.n6854 out.n6853 0.047
R77123 out.n6850 out.n6842 0.047
R77124 out.n6987 out.n6977 0.047
R77125 out.n1700 out.n1697 0.047
R77126 out.n1821 out.n1820 0.047
R77127 out.n1823 out.n1822 0.047
R77128 out.n1825 out.n1824 0.047
R77129 out.n1827 out.n1826 0.047
R77130 out.n1829 out.n1828 0.047
R77131 out.n1834 out.n1833 0.047
R77132 out.n7300 out.n7297 0.047
R77133 out.n7301 out.n7300 0.047
R77134 out.n2317 out.n2316 0.047
R77135 out.n2319 out.n2318 0.047
R77136 out.n2321 out.n2320 0.047
R77137 out.n2331 out.n2330 0.047
R77138 out.n2333 out.n2332 0.047
R77139 out.n2335 out.n2334 0.047
R77140 out.n2337 out.n2336 0.047
R77141 out.n7427 out.n7425 0.047
R77142 out.n7385 out.n7384 0.047
R77143 out.n7378 out.n7377 0.047
R77144 out.n7347 out.n7337 0.047
R77145 out.n7330 out.n7322 0.047
R77146 out.n2353 out.n2352 0.047
R77147 out.n2358 out.n2357 0.047
R77148 out.n7770 out.n7768 0.047
R77149 out.n7645 out.n7643 0.047
R77150 out.n7610 out.n7609 0.047
R77151 out.n7702 out.n7701 0.047
R77152 out.n2658 out.n2655 0.047
R77153 out.n2705 out.n2704 0.047
R77154 out.n2707 out.n2705 0.047
R77155 out.n2707 out.n2706 0.047
R77156 ldomc_0.out out.n2 0.047
R77157 out.n1321 out.n1320 0.047
R77158 out.n11307 out.n11306 0.047
R77159 out.n1482 out.n1481 0.046
R77160 out.n2329 out.n2328 0.046
R77161 out.n10877 out.n10876 0.046
R77162 out.n12340 out.n12328 0.046
R77163 out.n12111 out.n12110 0.046
R77164 out.n13500 out.n13499 0.046
R77165 out.n13382 out.n13381 0.046
R77166 out.n10968 out.n10967 0.046
R77167 out.n10858 out.n10857 0.046
R77168 out.n13955 out.n13954 0.046
R77169 out.n13837 out.n13836 0.046
R77170 out.n14467 out.n14466 0.046
R77171 out.n14429 out.n14428 0.046
R77172 out.n14414 out.n14413 0.046
R77173 out.n5141 out.n5140 0.046
R77174 out.n5103 out.n5102 0.046
R77175 out.n5088 out.n5087 0.046
R77176 out.n1058 out.n1057 0.046
R77177 out.n2901 out.n2899 0.046
R77178 out.n5843 out.n5842 0.046
R77179 out.n2913 out.n2912 0.046
R77180 out.n2915 out.n2914 0.046
R77181 out.n5445 out.n5444 0.046
R77182 out.n5441 out.n5440 0.046
R77183 out.n1468 out.n1467 0.046
R77184 out.n1492 out.n1491 0.046
R77185 out.n1502 out.n1501 0.046
R77186 out.n1504 out.n1503 0.046
R77187 out.n1805 out.n1803 0.046
R77188 out.n6977 out.n6976 0.046
R77189 out.n1817 out.n1816 0.046
R77190 out.n1819 out.n1818 0.046
R77191 out.n7303 out.n7302 0.046
R77192 out.n7299 out.n7298 0.046
R77193 out.n2315 out.n2314 0.046
R77194 out.n2339 out.n2338 0.046
R77195 out.n2349 out.n2348 0.046
R77196 out.n2351 out.n2350 0.046
R77197 out.n2537 out.n2535 0.046
R77198 out.n2583 out.n2582 0.046
R77199 out.n7630 out.n7629 0.046
R77200 out.n7726 out.n7725 0.046
R77201 out.n7717 out.n7716 0.046
R77202 out.n2689 out.n2688 0.046
R77203 out.n12130 out.n12129 0.046
R77204 out.n2928 out.n2927 0.046
R77205 out.n1832 out.n1831 0.046
R77206 out.n12569 out.n12568 0.046
R77207 out.n12995 out.n12994 0.046
R77208 out.n11710 out.n11709 0.046
R77209 out.n10443 out.n10442 0.046
R77210 out.n12161 out.n12160 0.046
R77211 out.n6090 out.n5894 0.046
R77212 out.n5314 out.n5313 0.046
R77213 out.n13402 out.n13401 0.046
R77214 out.n13857 out.n13856 0.046
R77215 out.n13435 out.n13434 0.046
R77216 out.n13890 out.n13889 0.046
R77217 out.n12722 out.n12721 0.046
R77218 out.n12602 out.n12601 0.046
R77219 out.n11445 out.n11444 0.046
R77220 out.n11335 out.n11334 0.046
R77221 out.n11018 out.n11017 0.045
R77222 out.n10908 out.n10907 0.045
R77223 out.n14509 out.n14508 0.045
R77224 out.n14450 out.n14449 0.045
R77225 out.n14395 out.n14394 0.045
R77226 out.n5124 out.n5123 0.045
R77227 out.n1047 out.n1046 0.045
R77228 out.n13026 out.n13025 0.045
R77229 out.n11741 out.n11740 0.045
R77230 out.n10474 out.n10473 0.045
R77231 out.n6123 out.n6122 0.045
R77232 out.n13141 out.n13140 0.045
R77233 out.n11856 out.n11855 0.045
R77234 out.n10589 out.n10588 0.045
R77235 out.n12276 out.n12275 0.045
R77236 out.n13556 out.n13555 0.045
R77237 out.n14011 out.n14010 0.045
R77238 out.n1480 out.n1479 0.045
R77239 out.n2327 out.n2326 0.045
R77240 out.n12782 out.n12770 0.045
R77241 out.n11395 out.n11394 0.045
R77242 out.n11288 out.n11287 0.045
R77243 out.n14520 out.n14519 0.045
R77244 out.n14471 out.n14470 0.045
R77245 out.n14469 out.n14468 0.045
R77246 out.n14436 out.n14435 0.045
R77247 out.n14175 out.n14174 0.045
R77248 out.n5145 out.n5144 0.045
R77249 out.n5143 out.n5142 0.045
R77250 out.n5110 out.n5109 0.045
R77251 out.n1051 out.n1050 0.045
R77252 out.n1473 out.n1472 0.045
R77253 out.n1510 out.n1509 0.045
R77254 out.n1262 out.n1260 0.045
R77255 out.n5265 out.n5264 0.045
R77256 out.n1316 out.n1315 0.045
R77257 out.n2320 out.n2319 0.045
R77258 out.n2357 out.n2356 0.045
R77259 out.n7127 out.n7126 0.045
R77260 out.n2574 out.n2573 0.045
R77261 out.n2685 out.n2684 0.045
R77262 out.n5755 out.n5754 0.044
R77263 out.n6332 out.n6331 0.044
R77264 out.n6889 out.n6888 0.044
R77265 out.n13001 out.n13000 0.044
R77266 out.n13058 out.n13056 0.044
R77267 out.n12954 out.n12952 0.044
R77268 out.n12136 out.n12135 0.044
R77269 out.n12193 out.n12191 0.044
R77270 out.n12089 out.n12087 0.044
R77271 out.n11367 out.n11365 0.044
R77272 out.n11266 out.n11264 0.044
R77273 out.n11082 out.n11070 0.044
R77274 out.n10883 out.n10882 0.044
R77275 out.n10940 out.n10938 0.044
R77276 out.n10836 out.n10834 0.044
R77277 out.n11716 out.n11715 0.044
R77278 out.n11773 out.n11771 0.044
R77279 out.n11669 out.n11667 0.044
R77280 out.n10449 out.n10448 0.044
R77281 out.n10506 out.n10504 0.044
R77282 out.n10402 out.n10400 0.044
R77283 out.n14525 out.n14524 0.044
R77284 out.n14518 out.n14517 0.044
R77285 out.n14494 out.n14493 0.044
R77286 out.n14474 out.n14473 0.044
R77287 out.n14434 out.n14433 0.044
R77288 out.n14432 out.n14431 0.044
R77289 out.n14413 out.n14386 0.044
R77290 out.n5148 out.n5147 0.044
R77291 out.n5108 out.n5107 0.044
R77292 out.n5106 out.n5105 0.044
R77293 out.n1017 out.n1014 0.044
R77294 out.n5087 out.n5075 0.044
R77295 out.n1053 out.n1052 0.044
R77296 out.n1078 out.n976 0.044
R77297 out.n2898 out.n2896 0.044
R77298 out.n2924 out.n2923 0.044
R77299 out.n2931 out.n2930 0.044
R77300 out.n5422 out.n5421 0.044
R77301 out.n1485 out.n1484 0.044
R77302 out.n5479 out.n5478 0.044
R77303 out.n1524 out.n1523 0.044
R77304 out.n5232 out.n5230 0.044
R77305 out.n5376 out.n5177 0.044
R77306 out.n1182 out.n1181 0.044
R77307 out.n6608 out.n6607 0.044
R77308 out.n2022 out.n2020 0.044
R77309 out.n6308 out.n6307 0.044
R77310 out.n2053 out.n2052 0.044
R77311 out.n2060 out.n2059 0.044
R77312 out.n6150 out.n6148 0.044
R77313 out.n6096 out.n6095 0.044
R77314 out.n6051 out.n6049 0.044
R77315 out.n1563 out.n1560 0.044
R77316 out.n5942 out.n5941 0.044
R77317 out.n1589 out.n1588 0.044
R77318 out.n1802 out.n1800 0.044
R77319 out.n1828 out.n1827 0.044
R77320 out.n1835 out.n1834 0.044
R77321 out.n7283 out.n7282 0.044
R77322 out.n2332 out.n2331 0.044
R77323 out.n7337 out.n7336 0.044
R77324 out.n2371 out.n2370 0.044
R77325 out.n7199 out.n7197 0.044
R77326 out.n7076 out.n7073 0.044
R77327 out.n7062 out.n7060 0.044
R77328 out.n2462 out.n2460 0.044
R77329 out.n2441 out.n2438 0.044
R77330 out.n10121 out.n10096 0.044
R77331 out.n7715 out.n7714 0.044
R77332 out.n12667 out.n12666 0.043
R77333 out.n12549 out.n12548 0.043
R77334 out.n11509 out.n11497 0.043
R77335 out.n5731 out.n5730 0.043
R77336 out.n1525 out.n1524 0.043
R77337 out.n6865 out.n6864 0.043
R77338 out.n2372 out.n2371 0.043
R77339 out.n2148 out.n2147 0.042
R77340 out.n1509 out.n1508 0.042
R77341 out.n2356 out.n2355 0.042
R77342 out.n9455 out.n9453 0.042
R77343 out.n12830 out.n12829 0.042
R77344 out.n12371 out.n12370 0.042
R77345 out.n11542 out.n11541 0.042
R77346 out.n11115 out.n11114 0.042
R77347 out.n11951 out.n11950 0.042
R77348 out.n10684 out.n10683 0.042
R77349 out.n1122 out.n1121 0.042
R77350 out.n6098 out.n6097 0.042
R77351 out.n10251 out.n10248 0.042
R77352 out.n5838 out.n5837 0.042
R77353 out.n6410 out.n6409 0.042
R77354 out.n6972 out.n6971 0.042
R77355 out.n7793 out.n7792 0.042
R77356 out.n2676 out.n2675 0.042
R77357 out.n6553 out.n6552 0.042
R77358 out.n1580 out.n1579 0.042
R77359 out.n1171 out.n1170 0.041
R77360 out.n2562 out.n2561 0.041
R77361 out.n14426 out.n14425 0.041
R77362 out.n5100 out.n5099 0.041
R77363 out.n14261 out.n14260 0.041
R77364 out.n957 out.n956 0.041
R77365 out.n1897 out.n1896 0.041
R77366 out.n1590 out.n1589 0.041
R77367 out.n2773 out.n2772 0.041
R77368 out.n1466 out.n1465 0.041
R77369 out.n1677 out.n1676 0.041
R77370 out.n2313 out.n2312 0.041
R77371 out.n10171 out.n10170 0.041
R77372 out.n10135 out.n10134 0.041
R77373 out.n12968 out.n12967 0.041
R77374 out.n12103 out.n12102 0.041
R77375 out.n11280 out.n11279 0.041
R77376 out.n10850 out.n10849 0.041
R77377 out.n11683 out.n11682 0.041
R77378 out.n10416 out.n10415 0.041
R77379 out.n1066 out.n1063 0.041
R77380 out.n5249 out.n5248 0.041
R77381 out.n2147 out.n2146 0.041
R77382 out.n6066 out.n6065 0.041
R77383 out.n7218 out.n7217 0.041
R77384 out.n11429 out.n11428 0.041
R77385 out.n11324 out.n11323 0.041
R77386 out.n11205 out.n11204 0.041
R77387 out.n1494 out.n1493 0.041
R77388 out.n2341 out.n2340 0.041
R77389 out.n12260 out.n12259 0.041
R77390 out.n12150 out.n12149 0.041
R77391 out.n12028 out.n12027 0.041
R77392 out.n11002 out.n11001 0.041
R77393 out.n10897 out.n10896 0.041
R77394 out.n10775 out.n10774 0.041
R77395 out.n10964 out.n10963 0.041
R77396 out.n11391 out.n11390 0.041
R77397 out.n12217 out.n12216 0.04
R77398 out.n12663 out.n12662 0.04
R77399 out.n13496 out.n13495 0.04
R77400 out.n13951 out.n13950 0.04
R77401 out.n13082 out.n13081 0.04
R77402 out.n11797 out.n11796 0.04
R77403 out.n10530 out.n10529 0.04
R77404 out.n13125 out.n13124 0.04
R77405 out.n13015 out.n13014 0.04
R77406 out.n12894 out.n12893 0.04
R77407 out.n11840 out.n11839 0.04
R77408 out.n11730 out.n11729 0.04
R77409 out.n11609 out.n11608 0.04
R77410 out.n10573 out.n10572 0.04
R77411 out.n10463 out.n10462 0.04
R77412 out.n10342 out.n10341 0.04
R77413 out.n6112 out.n6111 0.04
R77414 out.n6000 out.n5999 0.04
R77415 out.n10207 out.n10205 0.04
R77416 out.n12869 out.n12868 0.04
R77417 out.n13202 out.n13199 0.04
R77418 out.n13211 out.n13207 0.04
R77419 out.n12435 out.n12434 0.04
R77420 out.n12788 out.n12784 0.04
R77421 out.n12452 out.n12451 0.04
R77422 out.n12516 out.n12514 0.04
R77423 out.n12541 out.n12540 0.04
R77424 out.n12002 out.n12001 0.04
R77425 out.n12337 out.n12334 0.04
R77426 out.n12346 out.n12342 0.04
R77427 out.n13279 out.n13278 0.04
R77428 out.n13622 out.n13618 0.04
R77429 out.n13296 out.n13295 0.04
R77430 out.n13349 out.n13347 0.04
R77431 out.n13374 out.n13373 0.04
R77432 out.n11167 out.n11166 0.04
R77433 out.n11506 out.n11503 0.04
R77434 out.n11515 out.n11511 0.04
R77435 out.n10744 out.n10743 0.04
R77436 out.n11079 out.n11076 0.04
R77437 out.n11088 out.n11084 0.04
R77438 out.n11584 out.n11583 0.04
R77439 out.n11917 out.n11914 0.04
R77440 out.n11926 out.n11922 0.04
R77441 out.n13734 out.n13733 0.04
R77442 out.n14077 out.n14073 0.04
R77443 out.n13751 out.n13750 0.04
R77444 out.n13804 out.n13802 0.04
R77445 out.n13829 out.n13828 0.04
R77446 out.n10317 out.n10316 0.04
R77447 out.n10650 out.n10647 0.04
R77448 out.n10659 out.n10655 0.04
R77449 out.n14196 out.n14192 0.04
R77450 out.n14533 out.n14530 0.04
R77451 out.n14361 out.n14360 0.04
R77452 out.n14292 out.n14289 0.04
R77453 out.n14281 out.n14277 0.04
R77454 out.n5050 out.n5049 0.04
R77455 out.n4978 out.n4975 0.04
R77456 out.n4967 out.n4963 0.04
R77457 out.n5685 out.n5683 0.04
R77458 out.n5714 out.n5713 0.04
R77459 out.n5639 out.n5638 0.04
R77460 out.n2789 out.n2785 0.04
R77461 out.n1406 out.n1404 0.04
R77462 out.n5454 out.n5452 0.04
R77463 out.n5558 out.n5556 0.04
R77464 out.n5588 out.n5587 0.04
R77465 out.n5396 out.n5395 0.04
R77466 out.n1502 out.n1392 0.04
R77467 out.n1388 out.n1384 0.04
R77468 out.n1191 out.n1187 0.04
R77469 out.n5190 out.n5189 0.04
R77470 out.n6619 out.n6497 0.04
R77471 out.n6712 out.n6710 0.04
R77472 out.n6742 out.n6741 0.04
R77473 out.n6455 out.n6454 0.04
R77474 out.n2128 out.n2126 0.04
R77475 out.n2110 out.n2106 0.04
R77476 out.n6262 out.n6260 0.04
R77477 out.n6291 out.n6290 0.04
R77478 out.n6211 out.n6210 0.04
R77479 out.n1913 out.n1909 0.04
R77480 out.n5963 out.n5962 0.04
R77481 out.n5878 out.n5877 0.04
R77482 out.n6819 out.n6817 0.04
R77483 out.n6848 out.n6847 0.04
R77484 out.n6773 out.n6772 0.04
R77485 out.n1693 out.n1689 0.04
R77486 out.n2250 out.n2248 0.04
R77487 out.n7312 out.n7310 0.04
R77488 out.n7416 out.n7414 0.04
R77489 out.n7446 out.n7445 0.04
R77490 out.n7257 out.n7256 0.04
R77491 out.n2349 out.n2236 0.04
R77492 out.n2232 out.n2228 0.04
R77493 out.n7110 out.n7109 0.04
R77494 out.n7023 out.n7022 0.04
R77495 out.n7666 out.n7664 0.04
R77496 out.n7694 out.n7693 0.04
R77497 out.n7484 out.n7483 0.04
R77498 out.n2652 out.n2648 0.04
R77499 out.n14330 out.n14329 0.04
R77500 out.n5017 out.n5016 0.04
R77501 out.n2576 out.n2575 0.039
R77502 out.n10189 out.n10188 0.039
R77503 out.n10131 out.n10130 0.039
R77504 out.n10120 out.n10119 0.039
R77505 out.n12889 out.n12888 0.039
R77506 out.n12022 out.n12021 0.039
R77507 out.n11190 out.n11189 0.039
R77508 out.n10764 out.n10763 0.039
R77509 out.n11604 out.n11603 0.039
R77510 out.n10337 out.n10336 0.039
R77511 out.n984 out.n980 0.039
R77512 out.n5470 out.n5469 0.039
R77513 out.n6634 out.n6633 0.039
R77514 out.n6073 out.n6072 0.039
R77515 out.n7328 out.n7327 0.039
R77516 out.n5744 out.n5648 0.039
R77517 out.n6878 out.n6782 0.039
R77518 out.n7140 out.n7046 0.039
R77519 out.n1500 out.n1494 0.039
R77520 out.n2347 out.n2341 0.039
R77521 out.n6321 out.n6225 0.039
R77522 out.n1133 out.n1132 0.038
R77523 out.n9460 out.n9455 0.038
R77524 out.n2704 out.n2702 0.038
R77525 out.n12704 out.n12703 0.038
R77526 out.n10120 out.n10108 0.038
R77527 out.n1508 out.n1507 0.038
R77528 out.n2355 out.n2354 0.038
R77529 out.n11946 out.n11945 0.038
R77530 out.n10679 out.n10678 0.038
R77531 out.n9435 out.n9429 0.038
R77532 out.n7704 out.n7498 0.038
R77533 out.n13538 out.n13537 0.038
R77534 out.n13993 out.n13992 0.038
R77535 out.n12591 out.n12590 0.037
R77536 out.n12469 out.n12468 0.037
R77537 out.n5511 out.n5510 0.037
R77538 out.n7369 out.n7368 0.037
R77539 out.n13424 out.n13423 0.037
R77540 out.n13302 out.n13301 0.037
R77541 out.n13879 out.n13878 0.037
R77542 out.n13757 out.n13756 0.037
R77543 out.n6675 out.n6674 0.037
R77544 out.n12366 out.n12365 0.037
R77545 out.n1523 out.n1521 0.037
R77546 out.n2370 out.n2368 0.037
R77547 out.n1108 out.n1104 0.037
R77548 out.n2123 out.n2118 0.037
R77549 out.n9441 out.n9430 0.036
R77550 out.n2145 out.n2144 0.036
R77551 out.n9444 out.n9431 0.036
R77552 out.n9452 out.n9451 0.036
R77553 out.n13091 out.n13090 0.036
R77554 out.n13112 out.n13111 0.036
R77555 out.n12942 out.n12940 0.036
R77556 out.n12934 out.n12933 0.036
R77557 out.n12751 out.n12750 0.036
R77558 out.n12779 out.n12775 0.036
R77559 out.n12578 out.n12577 0.036
R77560 out.n12512 out.n12509 0.036
R77561 out.n12226 out.n12225 0.036
R77562 out.n12247 out.n12246 0.036
R77563 out.n12077 out.n12075 0.036
R77564 out.n12069 out.n12068 0.036
R77565 out.n13585 out.n13584 0.036
R77566 out.n13613 out.n13609 0.036
R77567 out.n13411 out.n13410 0.036
R77568 out.n13345 out.n13342 0.036
R77569 out.n11400 out.n11399 0.036
R77570 out.n11416 out.n11415 0.036
R77571 out.n11254 out.n11252 0.036
R77572 out.n11246 out.n11245 0.036
R77573 out.n10973 out.n10972 0.036
R77574 out.n10989 out.n10988 0.036
R77575 out.n10824 out.n10822 0.036
R77576 out.n10816 out.n10815 0.036
R77577 out.n11806 out.n11805 0.036
R77578 out.n11827 out.n11826 0.036
R77579 out.n11657 out.n11655 0.036
R77580 out.n11649 out.n11648 0.036
R77581 out.n14040 out.n14039 0.036
R77582 out.n14068 out.n14064 0.036
R77583 out.n13866 out.n13865 0.036
R77584 out.n13800 out.n13797 0.036
R77585 out.n10539 out.n10538 0.036
R77586 out.n10560 out.n10559 0.036
R77587 out.n10390 out.n10388 0.036
R77588 out.n10382 out.n10381 0.036
R77589 out.n14227 out.n14226 0.036
R77590 out.n14350 out.n14349 0.036
R77591 out.n14337 out.n14336 0.036
R77592 out.n5039 out.n5038 0.036
R77593 out.n5024 out.n5023 0.036
R77594 out.n1080 out.n970 0.036
R77595 out.n960 out.n959 0.036
R77596 out.n5676 out.n5675 0.036
R77597 out.n5669 out.n5666 0.036
R77598 out.n2812 out.n2808 0.036
R77599 out.n5434 out.n5431 0.036
R77600 out.n5447 out.n5446 0.036
R77601 out.n5554 out.n5551 0.036
R77602 out.n5592 out.n5591 0.036
R77603 out.n1230 out.n1226 0.036
R77604 out.n1177 out.n1176 0.036
R77605 out.n1293 out.n1186 0.036
R77606 out.n6601 out.n6598 0.036
R77607 out.n6492 out.n6491 0.036
R77608 out.n6708 out.n6705 0.036
R77609 out.n6253 out.n6252 0.036
R77610 out.n6246 out.n6243 0.036
R77611 out.n1936 out.n1932 0.036
R77612 out.n6039 out.n6037 0.036
R77613 out.n6031 out.n6030 0.036
R77614 out.n1558 out.n1554 0.036
R77615 out.n5949 out.n5947 0.036
R77616 out.n6810 out.n6809 0.036
R77617 out.n6803 out.n6800 0.036
R77618 out.n1716 out.n1712 0.036
R77619 out.n7295 out.n7292 0.036
R77620 out.n7305 out.n7304 0.036
R77621 out.n7412 out.n7409 0.036
R77622 out.n7450 out.n7449 0.036
R77623 out.n7147 out.n7146 0.036
R77624 out.n7081 out.n7079 0.036
R77625 out.n7067 out.n7064 0.036
R77626 out.n2435 out.n2431 0.036
R77627 out.n7657 out.n7656 0.036
R77628 out.n7650 out.n7647 0.036
R77629 out.n7582 out.n7581 0.036
R77630 out.n11108 out.n11107 0.036
R77631 out.n13638 out.n13637 0.036
R77632 out.n14093 out.n14092 0.036
R77633 out.n1477 out.n1474 0.036
R77634 out.n2324 out.n2321 0.036
R77635 out.n2166 out.n2164 0.036
R77636 out.n1528 out.n1525 0.036
R77637 out.n2375 out.n2372 0.036
R77638 out.n1369 out.n1368 0.035
R77639 out.n2213 out.n2212 0.035
R77640 out.n2162 out.n2160 0.035
R77641 out.n5490 out.n5407 0.035
R77642 out.n7348 out.n7268 0.035
R77643 out.n1085 out.n950 0.035
R77644 out.n2513 out.n2512 0.035
R77645 out.n2569 out.n2568 0.035
R77646 out.n5607 out.n5389 0.035
R77647 out.n7464 out.n7250 0.035
R77648 out.n11535 out.n11534 0.035
R77649 out.n9450 out.n9449 0.035
R77650 out.n12804 out.n12803 0.035
R77651 out.n1304 out.n1303 0.035
R77652 out.n2048 out.n2047 0.035
R77653 out.n14252 out.n14251 0.035
R77654 out.n2768 out.n2767 0.035
R77655 out.n1464 out.n1463 0.035
R77656 out.n1672 out.n1671 0.035
R77657 out.n2308 out.n2307 0.035
R77658 out.n6654 out.n6476 0.035
R77659 out.n2003 out.n2002 0.035
R77660 out.n5988 out.n5929 0.035
R77661 out.n2879 out.n2878 0.035
R77662 out.n1783 out.n1782 0.035
R77663 out.n6573 out.n6571 0.034
R77664 out.n5304 out.n5303 0.034
R77665 out.n7158 out.n7157 0.034
R77666 out.n9673 out 0.034
R77667 out.n9449 out.n9448 0.034
R77668 out.n9451 out.n9450 0.034
R77669 out.n1521 out.n1520 0.034
R77670 out.n2368 out.n2367 0.034
R77671 out.n13238 out.n13237 0.033
R77672 out.n11947 out.n11569 0.033
R77673 out.n10680 out.n10302 0.033
R77674 out.n11197 out.n11196 0.033
R77675 out.n5500 out.n5499 0.033
R77676 out.n7358 out.n7357 0.033
R77677 out.n12459 out.n12458 0.033
R77678 out.n5956 out.n5955 0.033
R77679 out.n10214 out.n10207 0.033
R77680 out.n5850 out.n5849 0.033
R77681 out.n2780 out.n2776 0.033
R77682 out.n2911 out.n2807 0.033
R77683 out.n5444 out.n5429 0.033
R77684 out.n1381 out.n1377 0.033
R77685 out.n6617 out.n6615 0.033
R77686 out.n6746 out.n6745 0.033
R77687 out.n2103 out.n2099 0.033
R77688 out.n6422 out.n6421 0.033
R77689 out.n1904 out.n1900 0.033
R77690 out.n2035 out.n1931 0.033
R77691 out.n6182 out.n6181 0.033
R77692 out.n5947 out.n5943 0.033
R77693 out.n6984 out.n6983 0.033
R77694 out.n1684 out.n1680 0.033
R77695 out.n1815 out.n1711 0.033
R77696 out.n7302 out.n7290 0.033
R77697 out.n2225 out.n2221 0.033
R77698 out.n7079 out.n7076 0.033
R77699 out.n2459 out.n2455 0.033
R77700 out.n2423 out.n2422 0.033
R77701 out.n2644 out.n2640 0.033
R77702 out.n2662 out.n2661 0.033
R77703 out.n5991 out.n5921 0.033
R77704 out.n1479 out.n1477 0.033
R77705 out.n2326 out.n2324 0.033
R77706 out.n7592 out.n7591 0.033
R77707 out.n6664 out.n6663 0.033
R77708 out.n6627 out.n6626 0.032
R77709 out.n1520 out.n1518 0.032
R77710 out.n2367 out.n2365 0.032
R77711 out.n1110 out.n1108 0.032
R77712 out.n2160 out.n2159 0.032
R77713 out.n2683 out.n2682 0.032
R77714 out.n1587 out.n1586 0.032
R77715 out.n10242 out.n10239 0.032
R77716 out.n10134 out.n10131 0.032
R77717 out.n7797 out.n7796 0.032
R77718 out.n2450 out.n2449 0.032
R77719 out.n12806 out.n12805 0.032
R77720 out.n5764 out.n5763 0.032
R77721 out.n6341 out.n6340 0.032
R77722 out.n6898 out.n6897 0.032
R77723 out.n13640 out.n13639 0.032
R77724 out.n14095 out.n14094 0.032
R77725 out.n1518 out.n1514 0.032
R77726 out.n2365 out.n2361 0.032
R77727 out.n13375 out.n13374 0.032
R77728 out.n13830 out.n13829 0.032
R77729 out.n12542 out.n12541 0.032
R77730 out.n7219 out.n7218 0.032
R77731 out.n14530 out.n14529 0.032
R77732 out.n5250 out.n5249 0.032
R77733 out.n6571 out.n6568 0.032
R77734 out.n5589 out.n5588 0.032
R77735 out.n7447 out.n7446 0.032
R77736 out.n6743 out.n6742 0.032
R77737 out.n1929 out.n1928 0.031
R77738 out.n1603 out.n1601 0.031
R77739 out.n5372 out.n5371 0.031
R77740 out.n11110 out.n11109 0.031
R77741 out.n14550 out.n14549 0.031
R77742 out.n7724 out.n7723 0.031
R77743 out.n7628 out.n7627 0.031
R77744 out.n2159 out.n2157 0.031
R77745 out.n11537 out.n11536 0.031
R77746 out.n12368 out.n12367 0.031
R77747 out.n12713 out.n12712 0.031
R77748 out.n5462 out.n5461 0.031
R77749 out.n7320 out.n7319 0.031
R77750 out.n10247 out.n10246 0.031
R77751 out.n10169 out.n10168 0.031
R77752 out.n13223 out.n13220 0.031
R77753 out.n13081 out.n13080 0.031
R77754 out.n12793 out.n12792 0.031
R77755 out.n12659 out.n12656 0.031
R77756 out.n12358 out.n12355 0.031
R77757 out.n12216 out.n12215 0.031
R77758 out.n13627 out.n13626 0.031
R77759 out.n13492 out.n13489 0.031
R77760 out.n11527 out.n11524 0.031
R77761 out.n11390 out.n11389 0.031
R77762 out.n11100 out.n11097 0.031
R77763 out.n10963 out.n10962 0.031
R77764 out.n11938 out.n11935 0.031
R77765 out.n11796 out.n11795 0.031
R77766 out.n14082 out.n14081 0.031
R77767 out.n13947 out.n13944 0.031
R77768 out.n10671 out.n10668 0.031
R77769 out.n10529 out.n10528 0.031
R77770 out.n14485 out.n14482 0.031
R77771 out.n14425 out.n14424 0.031
R77772 out.n5159 out.n5156 0.031
R77773 out.n5099 out.n5098 0.031
R77774 out.n6178 out.n6172 0.031
R77775 out.n2 out.n1 0.031
R77776 out.n11948 out.n11947 0.031
R77777 out.n10681 out.n10680 0.031
R77778 out.n2805 out.n2804 0.031
R77779 out.n1709 out.n1708 0.031
R77780 out.n13547 out.n13546 0.031
R77781 out.n14002 out.n14001 0.031
R77782 out.n12104 out.n12103 0.031
R77783 out.n10851 out.n10850 0.031
R77784 out.n11436 out.n11435 0.031
R77785 out.n11009 out.n11008 0.031
R77786 out.n11281 out.n11280 0.031
R77787 out.n1601 out.n1597 0.031
R77788 out.n9442 out.n9435 0.031
R77789 out.n1063 out.n1062 0.031
R77790 out.n6284 out.n6283 0.031
R77791 out.n6411 out.n6410 0.031
R77792 out.n12969 out.n12968 0.031
R77793 out.n11684 out.n11683 0.031
R77794 out.n10417 out.n10416 0.031
R77795 out.n5707 out.n5706 0.031
R77796 out.n5839 out.n5838 0.031
R77797 out.n6841 out.n6840 0.031
R77798 out.n6973 out.n6972 0.031
R77799 out.n6067 out.n6066 0.031
R77800 out.n10101 out.n10097 0.031
R77801 out.n7688 out.n7687 0.031
R77802 out.n7794 out.n7793 0.031
R77803 out.n2157 out.n2153 0.031
R77804 out.n12267 out.n12266 0.031
R77805 out.n2578 out.n2576 0.03
R77806 out.n13132 out.n13131 0.03
R77807 out.n11847 out.n11846 0.03
R77808 out.n10580 out.n10579 0.03
R77809 out.n5463 out.n5462 0.03
R77810 out.n7321 out.n7320 0.03
R77811 out.n10262 out.n10259 0.03
R77812 out.n10229 out.n10228 0.03
R77813 out.n10196 out.n10194 0.03
R77814 out.n10167 out.n10166 0.03
R77815 out.n10165 out.n10164 0.03
R77816 out.n10145 out.n10144 0.03
R77817 out.n13217 out.n13215 0.03
R77818 out.n13079 out.n13078 0.03
R77819 out.n12797 out.n12794 0.03
R77820 out.n12662 out.n12661 0.03
R77821 out.n12535 out.n12534 0.03
R77822 out.n12352 out.n12350 0.03
R77823 out.n12214 out.n12213 0.03
R77824 out.n13631 out.n13628 0.03
R77825 out.n13495 out.n13494 0.03
R77826 out.n13368 out.n13367 0.03
R77827 out.n11521 out.n11519 0.03
R77828 out.n11388 out.n11387 0.03
R77829 out.n11094 out.n11092 0.03
R77830 out.n10961 out.n10960 0.03
R77831 out.n11932 out.n11930 0.03
R77832 out.n11794 out.n11793 0.03
R77833 out.n14086 out.n14083 0.03
R77834 out.n13950 out.n13949 0.03
R77835 out.n13823 out.n13822 0.03
R77836 out.n10665 out.n10663 0.03
R77837 out.n10527 out.n10526 0.03
R77838 out.n14542 out.n14539 0.03
R77839 out.n14479 out.n14477 0.03
R77840 out.n14423 out.n14422 0.03
R77841 out.n5153 out.n5151 0.03
R77842 out.n5097 out.n5096 0.03
R77843 out.n5701 out.n5699 0.03
R77844 out.n5834 out.n5831 0.03
R77845 out.n5825 out.n5822 0.03
R77846 out.n5581 out.n5578 0.03
R77847 out.n5247 out.n5246 0.03
R77848 out.n5359 out.n5358 0.03
R77849 out.n5357 out.n5356 0.03
R77850 out.n5384 out.n5381 0.03
R77851 out.n5378 out.n5376 0.03
R77852 out.n1281 out.n1277 0.03
R77853 out.n6735 out.n6732 0.03
R77854 out.n6278 out.n6276 0.03
R77855 out.n6406 out.n6403 0.03
R77856 out.n6397 out.n6394 0.03
R77857 out.n6171 out.n6170 0.03
R77858 out.n6190 out.n6188 0.03
R77859 out.n6835 out.n6833 0.03
R77860 out.n6968 out.n6965 0.03
R77861 out.n6959 out.n6956 0.03
R77862 out.n7439 out.n7436 0.03
R77863 out.n7097 out.n7095 0.03
R77864 out.n7216 out.n7215 0.03
R77865 out.n7682 out.n7680 0.03
R77866 out.n7789 out.n7786 0.03
R77867 out.n7780 out.n7777 0.03
R77868 out.n14503 out.n14502 0.03
R77869 out.n1998 out.n1997 0.03
R77870 out.n14441 out.n14440 0.03
R77871 out.n5115 out.n5114 0.03
R77872 out.n1037 out.n1036 0.03
R77873 out.n2520 out.n2519 0.03
R77874 out.n2874 out.n2873 0.03
R77875 out.n1778 out.n1777 0.03
R77876 out.n1092 out.n1091 0.03
R77877 out.n1311 out.n1310 0.03
R77878 out.n7103 out.n7102 0.03
R77879 out.n2702 out.n2697 0.03
R77880 out.n1459 out.n1458 0.03
R77881 out.n2303 out.n2302 0.03
R77882 out.n5373 out.n5372 0.029
R77883 out.n11332 out.n11331 0.029
R77884 out.n11211 out.n11210 0.029
R77885 out.n10905 out.n10904 0.029
R77886 out.n10781 out.n10780 0.029
R77887 out.n7612 out.n7549 0.029
R77888 out.n6558 out.n6510 0.029
R77889 out.n2911 out.n2805 0.029
R77890 out.n1815 out.n1709 0.029
R77891 out.n12158 out.n12157 0.029
R77892 out.n12034 out.n12033 0.029
R77893 out.n1274 out.n1270 0.029
R77894 out.n10233 out.n10230 0.029
R77895 out.n10147 out.n10146 0.029
R77896 out.n10114 out.n10113 0.029
R77897 out.n10090 out.n10089 0.029
R77898 out.n13241 out.n13240 0.029
R77899 out.n13172 out.n13171 0.029
R77900 out.n13054 out.n13051 0.029
R77901 out.n12844 out.n12840 0.029
R77902 out.n12927 out.n12924 0.029
R77903 out.n12945 out.n12944 0.029
R77904 out.n12691 out.n12690 0.029
R77905 out.n12640 out.n12639 0.029
R77906 out.n12503 out.n12500 0.029
R77907 out.n12514 out.n12512 0.029
R77908 out.n11984 out.n11983 0.029
R77909 out.n12307 out.n12306 0.029
R77910 out.n12189 out.n12186 0.029
R77911 out.n12062 out.n12059 0.029
R77912 out.n12080 out.n12079 0.029
R77913 out.n13525 out.n13524 0.029
R77914 out.n13473 out.n13472 0.029
R77915 out.n13336 out.n13333 0.029
R77916 out.n13347 out.n13345 0.029
R77917 out.n11144 out.n11143 0.029
R77918 out.n11476 out.n11475 0.029
R77919 out.n11363 out.n11360 0.029
R77920 out.n11203 out.n11202 0.029
R77921 out.n11239 out.n11236 0.029
R77922 out.n11257 out.n11256 0.029
R77923 out.n10721 out.n10720 0.029
R77924 out.n11049 out.n11048 0.029
R77925 out.n10936 out.n10933 0.029
R77926 out.n10773 out.n10772 0.029
R77927 out.n10809 out.n10806 0.029
R77928 out.n10827 out.n10826 0.029
R77929 out.n11567 out.n11566 0.029
R77930 out.n11887 out.n11886 0.029
R77931 out.n11769 out.n11766 0.029
R77932 out.n11965 out.n11961 0.029
R77933 out.n11642 out.n11639 0.029
R77934 out.n11660 out.n11659 0.029
R77935 out.n13980 out.n13979 0.029
R77936 out.n13928 out.n13927 0.029
R77937 out.n13791 out.n13788 0.029
R77938 out.n13802 out.n13800 0.029
R77939 out.n10300 out.n10299 0.029
R77940 out.n10620 out.n10619 0.029
R77941 out.n10502 out.n10499 0.029
R77942 out.n10698 out.n10694 0.029
R77943 out.n10375 out.n10372 0.029
R77944 out.n10393 out.n10392 0.029
R77945 out.n14268 out.n14267 0.029
R77946 out.n14307 out.n14306 0.029
R77947 out.n14384 out.n14381 0.029
R77948 out.n4994 out.n4993 0.029
R77949 out.n5073 out.n5070 0.029
R77950 out.n956 out.n955 0.029
R77951 out.n964 out.n963 0.029
R77952 out.n5800 out.n5797 0.029
R77953 out.n5753 out.n5752 0.029
R77954 out.n5683 out.n5677 0.029
R77955 out.n5660 out.n5657 0.029
R77956 out.n5692 out.n5691 0.029
R77957 out.n2772 out.n2771 0.029
R77958 out.n2776 out.n2775 0.029
R77959 out.n1403 out.n1399 0.029
R77960 out.n1493 out.n1406 0.029
R77961 out.n1425 out.n1422 0.029
R77962 out.n5429 out.n5423 0.029
R77963 out.n5452 out.n5448 0.029
R77964 out.n5556 out.n5554 0.029
R77965 out.n5545 out.n5542 0.029
R77966 out.n1368 out.n1367 0.029
R77967 out.n1498 out.n1495 0.029
R77968 out.n5293 out.n5292 0.029
R77969 out.n5270 out.n5269 0.029
R77970 out.n5261 out.n5260 0.029
R77971 out.n5224 out.n5223 0.029
R77972 out.n5217 out.n5214 0.029
R77973 out.n1170 out.n1169 0.029
R77974 out.n6539 out.n6538 0.029
R77975 out.n6533 out.n6532 0.029
R77976 out.n6552 out.n6551 0.029
R77977 out.n6594 out.n6591 0.029
R77978 out.n6615 out.n6609 0.029
R77979 out.n6497 out.n6493 0.029
R77980 out.n6710 out.n6708 0.029
R77981 out.n6699 out.n6696 0.029
R77982 out.n2144 out.n2143 0.029
R77983 out.n6372 out.n6369 0.029
R77984 out.n6330 out.n6329 0.029
R77985 out.n6260 out.n6254 0.029
R77986 out.n6237 out.n6234 0.029
R77987 out.n6269 out.n6268 0.029
R77988 out.n1896 out.n1895 0.029
R77989 out.n1900 out.n1899 0.029
R77990 out.n6146 out.n6143 0.029
R77991 out.n6042 out.n6041 0.029
R77992 out.n6024 out.n6021 0.029
R77993 out.n5998 out.n5997 0.029
R77994 out.n1579 out.n1578 0.029
R77995 out.n1569 out.n1568 0.029
R77996 out.n6934 out.n6931 0.029
R77997 out.n6887 out.n6886 0.029
R77998 out.n6817 out.n6811 0.029
R77999 out.n6794 out.n6791 0.029
R78000 out.n6826 out.n6825 0.029
R78001 out.n1676 out.n1675 0.029
R78002 out.n1680 out.n1679 0.029
R78003 out.n2247 out.n2243 0.029
R78004 out.n2340 out.n2250 0.029
R78005 out.n2269 out.n2266 0.029
R78006 out.n2312 out.n2311 0.029
R78007 out.n7290 out.n7284 0.029
R78008 out.n7310 out.n7306 0.029
R78009 out.n7414 out.n7412 0.029
R78010 out.n7403 out.n7400 0.029
R78011 out.n2212 out.n2211 0.029
R78012 out.n2345 out.n2342 0.029
R78013 out.n7230 out.n7229 0.029
R78014 out.n7191 out.n7190 0.029
R78015 out.n7184 out.n7181 0.029
R78016 out.n7058 out.n7055 0.029
R78017 out.n2482 out.n2480 0.029
R78018 out.n2561 out.n2560 0.029
R78019 out.n2427 out.n2423 0.029
R78020 out.n2549 out.n2454 0.029
R78021 out.n7755 out.n7752 0.029
R78022 out.n7713 out.n7712 0.029
R78023 out.n7664 out.n7658 0.029
R78024 out.n7641 out.n7638 0.029
R78025 out.n7673 out.n7672 0.029
R78026 out.n2675 out.n2674 0.029
R78027 out.n2640 out.n2639 0.029
R78028 out.n13023 out.n13022 0.029
R78029 out.n12899 out.n12898 0.029
R78030 out.n11738 out.n11737 0.029
R78031 out.n11614 out.n11613 0.029
R78032 out.n10471 out.n10470 0.029
R78033 out.n10347 out.n10346 0.029
R78034 out.n6120 out.n6119 0.029
R78035 out.n6006 out.n6005 0.029
R78036 out.n7593 out.n7592 0.028
R78037 out.n2035 out.n1929 0.028
R78038 out.n10179 out.n10172 0.028
R78039 out.n6628 out.n6627 0.028
R78040 out.n5376 out.n5373 0.028
R78041 out.n1293 out.n1292 0.028
R78042 out.n12961 out.n12960 0.028
R78043 out.n12096 out.n12095 0.028
R78044 out.n11273 out.n11272 0.028
R78045 out.n10843 out.n10842 0.028
R78046 out.n11676 out.n11675 0.028
R78047 out.n10409 out.n10408 0.028
R78048 out.n1074 out.n1071 0.028
R78049 out.n5240 out.n5239 0.028
R78050 out.n6059 out.n6057 0.028
R78051 out.n7209 out.n7206 0.028
R78052 out.n5957 out.n5956 0.028
R78053 out.n2549 out.n2450 0.028
R78054 out.n12599 out.n12598 0.028
R78055 out.n12475 out.n12474 0.028
R78056 out.n5517 out.n5516 0.028
R78057 out.n7375 out.n7374 0.028
R78058 out.n1116 out.n1113 0.028
R78059 out.n7622 out.n7621 0.028
R78060 out.n13432 out.n13431 0.028
R78061 out.n13308 out.n13307 0.028
R78062 out.n13887 out.n13886 0.028
R78063 out.n13763 out.n13762 0.028
R78064 out.n2548 out.n2547 0.027
R78065 out.n6681 out.n6680 0.027
R78066 out.n6620 out.n6619 0.027
R78067 out.n7083 out.n7081 0.027
R78068 out.n1289 out.n1286 0.027
R78069 out.n7088 out.n7087 0.027
R78070 out.n2034 out.n2033 0.027
R78071 out.n6752 out.n6747 0.027
R78072 out.n5364 out.n5359 0.027
R78073 out.n12719 out.n12718 0.027
R78074 out.n11442 out.n11441 0.027
R78075 out.n11015 out.n11014 0.026
R78076 out.n5311 out.n5310 0.026
R78077 out.n2910 out.n2909 0.026
R78078 out.n1814 out.n1813 0.026
R78079 out.n1318 out.n1317 0.026
R78080 out.n5365 out.n5364 0.026
R78081 out.n7164 out.n7163 0.026
R78082 out.n5595 out.n5593 0.026
R78083 out.n7453 out.n7451 0.026
R78084 out.n12273 out.n12272 0.026
R78085 out.n13553 out.n13552 0.026
R78086 out.n14008 out.n14007 0.026
R78087 out.n13138 out.n13137 0.026
R78088 out.n11853 out.n11852 0.026
R78089 out.n10586 out.n10585 0.026
R78090 out.n10256 out.n10254 0.026
R78091 out.n10225 out.n10221 0.026
R78092 out.n10191 out.n10189 0.026
R78093 out.n10158 out.n10153 0.026
R78094 out.n5167 out.n5165 0.026
R78095 out.n1512 out.n1357 0.026
R78096 out.n2359 out.n2201 0.026
R78097 out.n2708 out.n2707 0.026
R78098 out.n2692 out.n2691 0.026
R78099 out.n7235 out.n7233 0.026
R78100 out.n3267 out.n3265 0.026
R78101 out.n3263 out.n3262 0.026
R78102 out.n3127 out.n3126 0.026
R78103 out.n14506 out.n14245 0.026
R78104 out.n14447 out.n14446 0.026
R78105 out.n5121 out.n5120 0.026
R78106 out.n1044 out.n1043 0.026
R78107 out.n1099 out.n1098 0.026
R78108 out.n1245 out.n1244 0.026
R78109 out.n5770 out.n5769 0.026
R78110 out.n6904 out.n6903 0.026
R78111 out.n7814 out.n7809 0.025
R78112 out.n5455 out.n5454 0.025
R78113 out.n7313 out.n7312 0.025
R78114 out.n2151 out.n2091 0.025
R78115 out.n12091 out.n12089 0.025
R78116 out.n7799 out.n7798 0.025
R78117 out.n10838 out.n10836 0.025
R78118 out.n6347 out.n6346 0.025
R78119 out.n7668 out.n7666 0.025
R78120 out.n7809 out.n7804 0.025
R78121 out.n11268 out.n11266 0.025
R78122 out.n1078 out.n1077 0.025
R78123 out.n5993 out.n5991 0.025
R78124 out.n5687 out.n5685 0.025
R78125 out.n6821 out.n6819 0.025
R78126 out.n12956 out.n12954 0.025
R78127 out.n11671 out.n11669 0.025
R78128 out.n10404 out.n10402 0.025
R78129 out.n1593 out.n1592 0.025
R78130 out.n6427 out.n6425 0.025
R78131 out.n12847 out.n12846 0.025
R78132 out.n11968 out.n11967 0.025
R78133 out.n10701 out.n10700 0.025
R78134 out.n6264 out.n6262 0.025
R78135 out.n5855 out.n5853 0.025
R78136 out.n6989 out.n6987 0.025
R78137 out.n10201 out.n10199 0.025
R78138 out.n12883 out.n12882 0.025
R78139 out.n13056 out.n13054 0.025
R78140 out.n12940 out.n12935 0.025
R78141 out.n12952 out.n12946 0.025
R78142 out.n12446 out.n12445 0.025
R78143 out.n12557 out.n12556 0.025
R78144 out.n12568 out.n12565 0.025
R78145 out.n12016 out.n12015 0.025
R78146 out.n12191 out.n12189 0.025
R78147 out.n12075 out.n12070 0.025
R78148 out.n12087 out.n12081 0.025
R78149 out.n13290 out.n13289 0.025
R78150 out.n13390 out.n13389 0.025
R78151 out.n13401 out.n13398 0.025
R78152 out.n11184 out.n11183 0.025
R78153 out.n11365 out.n11363 0.025
R78154 out.n11252 out.n11247 0.025
R78155 out.n11264 out.n11258 0.025
R78156 out.n10758 out.n10757 0.025
R78157 out.n10938 out.n10936 0.025
R78158 out.n10822 out.n10817 0.025
R78159 out.n10834 out.n10828 0.025
R78160 out.n11598 out.n11597 0.025
R78161 out.n11771 out.n11769 0.025
R78162 out.n11655 out.n11650 0.025
R78163 out.n11667 out.n11661 0.025
R78164 out.n13745 out.n13744 0.025
R78165 out.n13845 out.n13844 0.025
R78166 out.n13856 out.n13853 0.025
R78167 out.n10331 out.n10330 0.025
R78168 out.n10504 out.n10502 0.025
R78169 out.n10388 out.n10383 0.025
R78170 out.n10400 out.n10394 0.025
R78171 out.n14222 out.n14219 0.025
R78172 out.n14214 out.n14208 0.025
R78173 out.n14203 out.n14199 0.025
R78174 out.n14386 out.n14384 0.025
R78175 out.n991 out.n987 0.025
R78176 out.n5075 out.n5073 0.025
R78177 out.n5654 out.n5653 0.025
R78178 out.n2836 out.n2835 0.025
R78179 out.n2828 out.n2827 0.025
R78180 out.n2821 out.n2817 0.025
R78181 out.n1412 out.n1408 0.025
R78182 out.n1420 out.n1419 0.025
R78183 out.n5412 out.n5408 0.025
R78184 out.n5419 out.n5418 0.025
R78185 out.n1374 out.n1370 0.025
R78186 out.n1500 out.n1498 0.025
R78187 out.n5230 out.n5225 0.025
R78188 out.n1198 out.n1194 0.025
R78189 out.n1169 out.n1166 0.025
R78190 out.n6530 out.n6529 0.025
R78191 out.n6523 out.n6519 0.025
R78192 out.n6481 out.n6477 0.025
R78193 out.n6488 out.n6487 0.025
R78194 out.n2136 out.n2132 0.025
R78195 out.n2123 out.n2121 0.025
R78196 out.n6231 out.n6230 0.025
R78197 out.n1960 out.n1959 0.025
R78198 out.n1952 out.n1951 0.025
R78199 out.n1945 out.n1941 0.025
R78200 out.n6148 out.n6146 0.025
R78201 out.n5900 out.n5899 0.025
R78202 out.n6049 out.n6043 0.025
R78203 out.n6037 out.n6032 0.025
R78204 out.n5934 out.n5930 0.025
R78205 out.n5971 out.n5970 0.025
R78206 out.n1554 out.n1553 0.025
R78207 out.n6788 out.n6787 0.025
R78208 out.n1740 out.n1739 0.025
R78209 out.n1732 out.n1731 0.025
R78210 out.n1725 out.n1721 0.025
R78211 out.n2256 out.n2252 0.025
R78212 out.n2264 out.n2263 0.025
R78213 out.n7273 out.n7269 0.025
R78214 out.n7280 out.n7279 0.025
R78215 out.n2218 out.n2214 0.025
R78216 out.n2347 out.n2345 0.025
R78217 out.n7197 out.n7192 0.025
R78218 out.n7052 out.n7051 0.025
R78219 out.n7060 out.n7058 0.025
R78220 out.n2476 out.n2475 0.025
R78221 out.n2468 out.n2464 0.025
R78222 out.n2547 out.n2462 0.025
R78223 out.n2431 out.n2430 0.025
R78224 out.n7524 out.n7523 0.025
R78225 out.n7567 out.n7562 0.025
R78226 out.n7574 out.n7570 0.025
R78227 out.n7602 out.n7601 0.025
R78228 out.n9439 out.n9428 0.025
R78229 out.n6566 out.n6565 0.025
R78230 out.n1607 out.n1606 0.025
R78231 out.n5235 out.n5232 0.025
R78232 out.n2695 out.n2692 0.025
R78233 out.n7202 out.n7199 0.025
R78234 out.n7730 out.n7729 0.025
R78235 out.n7624 out.n7622 0.025
R78236 out.n2529 out.n2528 0.025
R78237 out.n5352 out.n5349 0.024
R78238 out.n1595 out.n1593 0.024
R78239 out.n2612 out.n2608 0.024
R78240 out.n1631 out.n1627 0.024
R78241 out.n7142 out.n7140 0.024
R78242 out.n12386 out.n12385 0.024
R78243 out.n7706 out.n7704 0.024
R78244 out.n6053 out.n6051 0.024
R78245 out.n1879 out.n1876 0.024
R78246 out.n7773 out.n7770 0.024
R78247 out.n5871 out.n5870 0.024
R78248 out.n11198 out.n11197 0.024
R78249 out.n3224 out.n3223 0.024
R78250 out.n6390 out.n6387 0.024
R78251 out.n5818 out.n5815 0.024
R78252 out.n6952 out.n6949 0.024
R78253 out.n2750 out.n2747 0.024
R78254 out.n1654 out.n1651 0.024
R78255 out.n6666 out.n6664 0.024
R78256 out.n13663 out.n13662 0.024
R78257 out.n13696 out.n13695 0.024
R78258 out.n6092 out.n6090 0.024
R78259 out.n12997 out.n12995 0.024
R78260 out.n11712 out.n11710 0.024
R78261 out.n10445 out.n10443 0.024
R78262 out.n2584 out.n2583 0.023
R78263 out.n1257 out.n1256 0.023
R78264 out.n12132 out.n12130 0.023
R78265 out.n2890 out.n2889 0.023
R78266 out.n2014 out.n2013 0.023
R78267 out.n1794 out.n1793 0.023
R78268 out.n2926 out.n2750 0.023
R78269 out.n1830 out.n1654 0.023
R78270 out.n6323 out.n6321 0.023
R78271 out.n9015 out.n8985 0.023
R78272 out.n16263 out.n16238 0.023
R78273 out.n16231 out.n16208 0.023
R78274 out.n17277 out.n17248 0.023
R78275 out.n16196 out.n16173 0.023
R78276 out.n16166 out.n16141 0.023
R78277 out.n16135 out.n16112 0.023
R78278 out.n16105 out.n16080 0.023
R78279 out.n16073 out.n15943 0.023
R78280 out.n15978 out.n15949 0.023
R78281 out.n15935 out.n15912 0.023
R78282 out.n16014 out.n15985 0.023
R78283 out.n15899 out.n15876 0.023
R78284 out.n15869 out.n15844 0.023
R78285 out.n15838 out.n15815 0.023
R78286 out.n15808 out.n15783 0.023
R78287 out.n15777 out.n15754 0.023
R78288 out.n15747 out.n15717 0.023
R78289 out.n15711 out.n15683 0.023
R78290 out.n15676 out.n15646 0.023
R78291 out.n15639 out.n15570 0.023
R78292 out.n15605 out.n15576 0.023
R78293 out.n15558 out.n15535 0.023
R78294 out.n15528 out.n15498 0.023
R78295 out.n15492 out.n15463 0.023
R78296 out.n15455 out.n15449 0.023
R78297 out.n16235 out.n16206 0.023
R78298 out.n15938 out.n15910 0.023
R78299 out.n15643 out.n15568 0.023
R78300 out.n15459 out.n15392 0.023
R78301 out.n15528 out.n15516 0.023
R78302 out.n15492 out.n15480 0.023
R78303 out.n15605 out.n15589 0.023
R78304 out.n15558 out.n15548 0.023
R78305 out.n15676 out.n15664 0.023
R78306 out.n15639 out.n15629 0.023
R78307 out.n15747 out.n15735 0.023
R78308 out.n15711 out.n15701 0.023
R78309 out.n15808 out.n15796 0.023
R78310 out.n15777 out.n15767 0.023
R78311 out.n15869 out.n15857 0.023
R78312 out.n15838 out.n15828 0.023
R78313 out.n16014 out.n15998 0.023
R78314 out.n15899 out.n15889 0.023
R78315 out.n15978 out.n15962 0.023
R78316 out.n15935 out.n15925 0.023
R78317 out.n16105 out.n16093 0.023
R78318 out.n16073 out.n16063 0.023
R78319 out.n16166 out.n16154 0.023
R78320 out.n16135 out.n16125 0.023
R78321 out.n17277 out.n17261 0.023
R78322 out.n16196 out.n16186 0.023
R78323 out.n16263 out.n16251 0.023
R78324 out.n16231 out.n16221 0.023
R78325 out.n9015 out.n9003 0.023
R78326 out.n14103 out.n13245 0.023
R78327 out.n9015 out.n9006 0.023
R78328 out.n9015 out.n9007 0.023
R78329 out.n15328 out.n15319 0.023
R78330 out.n15359 out.n15351 0.023
R78331 out.n15263 out.n15254 0.023
R78332 out.n15294 out.n15286 0.023
R78333 out.n15198 out.n15189 0.023
R78334 out.n15229 out.n15221 0.023
R78335 out.n15157 out.n15148 0.023
R78336 out.n8964 out.n8956 0.023
R78337 out.n15119 out.n15110 0.023
R78338 out.n8929 out.n8921 0.023
R78339 out.n15054 out.n15045 0.023
R78340 out.n15086 out.n15078 0.023
R78341 out.n14989 out.n14980 0.023
R78342 out.n15021 out.n15013 0.023
R78343 out.n14918 out.n14909 0.023
R78344 out.n14953 out.n14945 0.023
R78345 out.n14847 out.n14838 0.023
R78346 out.n14882 out.n14874 0.023
R78347 out.n14776 out.n14767 0.023
R78348 out.n14811 out.n14803 0.023
R78349 out.n14705 out.n14696 0.023
R78350 out.n14740 out.n14732 0.023
R78351 out.n14634 out.n14625 0.023
R78352 out.n14669 out.n14661 0.023
R78353 out.n14598 out.n14590 0.023
R78354 out.n15492 out.n15477 0.023
R78355 out.n9015 out.n8997 0.023
R78356 out.n14147 out.n14132 0.023
R78357 out.n9015 out.n9010 0.023
R78358 out.n14103 out.n11975 0.023
R78359 out.n14147 out.n14128 0.023
R78360 out.n14634 out.n14616 0.023
R78361 out.n14705 out.n14687 0.023
R78362 out.n14776 out.n14758 0.023
R78363 out.n14847 out.n14829 0.023
R78364 out.n14918 out.n14900 0.023
R78365 out.n14989 out.n14971 0.023
R78366 out.n15054 out.n15036 0.023
R78367 out.n15119 out.n15101 0.023
R78368 out.n15157 out.n15139 0.023
R78369 out.n15198 out.n15179 0.023
R78370 out.n15263 out.n15245 0.023
R78371 out.n15328 out.n15310 0.023
R78372 out.n9015 out.n8996 0.023
R78373 out.n9015 out.n8988 0.023
R78374 out.n9015 out.n8991 0.023
R78375 out.n15528 out.n15507 0.023
R78376 out.n15605 out.n15580 0.023
R78377 out.n15676 out.n15655 0.023
R78378 out.n15747 out.n15726 0.023
R78379 out.n15808 out.n15787 0.023
R78380 out.n15869 out.n15848 0.023
R78381 out.n16014 out.n15989 0.023
R78382 out.n15978 out.n15953 0.023
R78383 out.n16105 out.n16084 0.023
R78384 out.n16166 out.n16145 0.023
R78385 out.n17277 out.n17252 0.023
R78386 out.n9015 out.n8993 0.023
R78387 out.n16263 out.n16242 0.023
R78388 out.n15455 out.n15454 0.023
R78389 out.n9015 out.n9014 0.023
R78390 out.n17309 out.n8982 0.023
R78391 out.n17309 out.n9016 0.023
R78392 out.n7820 out.n7475 0.023
R78393 out.n7897 out.n7893 0.023
R78394 out.n7974 out.n7970 0.023
R78395 out.n8051 out.n8047 0.023
R78396 out.n8128 out.n8124 0.023
R78397 out.n8205 out.n8201 0.023
R78398 out.n8282 out.n8278 0.023
R78399 out.n8359 out.n8355 0.023
R78400 out.n8436 out.n8432 0.023
R78401 out.n8513 out.n8509 0.023
R78402 out.n8590 out.n8586 0.023
R78403 out.n8667 out.n8663 0.023
R78404 out.n8744 out.n8740 0.023
R78405 out.n8792 out.n8786 0.023
R78406 out.n3984 out.n3979 0.023
R78407 out.n3923 out.n3918 0.023
R78408 out.n3846 out.n3841 0.023
R78409 out.n3769 out.n3764 0.023
R78410 out.n3692 out.n3687 0.023
R78411 out.n3615 out.n3610 0.023
R78412 out.n3538 out.n3533 0.023
R78413 out.n3461 out.n3456 0.023
R78414 out.n3384 out.n3379 0.023
R78415 out.n3307 out.n3302 0.023
R78416 out.n3176 out.n3168 0.023
R78417 out.n3176 out.n3171 0.023
R78418 out.n3150 out.n3141 0.023
R78419 out.n2943 out.n2607 0.023
R78420 out.n7821 out.n5621 0.023
R78421 out.n7860 out.n7829 0.023
R78422 out.n7898 out.n7869 0.023
R78423 out.n7937 out.n7906 0.023
R78424 out.n7975 out.n7946 0.023
R78425 out.n8014 out.n7983 0.023
R78426 out.n8052 out.n8023 0.023
R78427 out.n8091 out.n8060 0.023
R78428 out.n8129 out.n8100 0.023
R78429 out.n8168 out.n8137 0.023
R78430 out.n8206 out.n8177 0.023
R78431 out.n8245 out.n8214 0.023
R78432 out.n8283 out.n8254 0.023
R78433 out.n8322 out.n8291 0.023
R78434 out.n8360 out.n8331 0.023
R78435 out.n8399 out.n8368 0.023
R78436 out.n8437 out.n8408 0.023
R78437 out.n8476 out.n8445 0.023
R78438 out.n8514 out.n8485 0.023
R78439 out.n8553 out.n8522 0.023
R78440 out.n8591 out.n8562 0.023
R78441 out.n8630 out.n8599 0.023
R78442 out.n8668 out.n8639 0.023
R78443 out.n8707 out.n8676 0.023
R78444 out.n8745 out.n8716 0.023
R78445 out.n8793 out.n8754 0.023
R78446 out.n8793 out.n8756 0.023
R78447 out.n3985 out.n3972 0.023
R78448 out.n3962 out.n3933 0.023
R78449 out.n3924 out.n3895 0.023
R78450 out.n3885 out.n3856 0.023
R78451 out.n3847 out.n3818 0.023
R78452 out.n3808 out.n3779 0.023
R78453 out.n3770 out.n3741 0.023
R78454 out.n3731 out.n3702 0.023
R78455 out.n3693 out.n3664 0.023
R78456 out.n3654 out.n3625 0.023
R78457 out.n3616 out.n3587 0.023
R78458 out.n3577 out.n3548 0.023
R78459 out.n3539 out.n3510 0.023
R78460 out.n3500 out.n3471 0.023
R78461 out.n3462 out.n3433 0.023
R78462 out.n3423 out.n3394 0.023
R78463 out.n3385 out.n3356 0.023
R78464 out.n3346 out.n3317 0.023
R78465 out.n3308 out.n3279 0.023
R78466 out.n3269 out.n3201 0.023
R78467 out.n3188 out.n3187 0.023
R78468 out.n3190 out.n3189 0.023
R78469 out.n3177 out.n3162 0.023
R78470 out.n3177 out.n3163 0.023
R78471 out.n3151 out.n3081 0.023
R78472 out.n3071 out.n3042 0.023
R78473 out.n3024 out.n2965 0.023
R78474 out.n56 out.n26 0.023
R78475 out.n2944 out.n1338 0.023
R78476 out.n2944 out.n1533 0.023
R78477 out.n2952 out.n1136 0.023
R78478 out.n2952 out.n1335 0.023
R78479 out.n3031 out.n2964 0.023
R78480 out.n3154 out.n3080 0.023
R78481 out.n3074 out.n3041 0.023
R78482 out.n3195 out.n3186 0.023
R78483 out.n3180 out.n3159 0.023
R78484 out.n3311 out.n3278 0.023
R78485 out.n3272 out.n3200 0.023
R78486 out.n3388 out.n3355 0.023
R78487 out.n3349 out.n3316 0.023
R78488 out.n3465 out.n3432 0.023
R78489 out.n3426 out.n3393 0.023
R78490 out.n3542 out.n3509 0.023
R78491 out.n3503 out.n3470 0.023
R78492 out.n3619 out.n3586 0.023
R78493 out.n3580 out.n3547 0.023
R78494 out.n3696 out.n3663 0.023
R78495 out.n3657 out.n3624 0.023
R78496 out.n3773 out.n3740 0.023
R78497 out.n3734 out.n3701 0.023
R78498 out.n3850 out.n3817 0.023
R78499 out.n3811 out.n3778 0.023
R78500 out.n3927 out.n3894 0.023
R78501 out.n3888 out.n3855 0.023
R78502 out.n3988 out.n3971 0.023
R78503 out.n3965 out.n3932 0.023
R78504 out.n8747 out.n8713 0.023
R78505 out.n8794 out.n8750 0.023
R78506 out.n8794 out.n8753 0.023
R78507 out.n8670 out.n8636 0.023
R78508 out.n8709 out.n8673 0.023
R78509 out.n8593 out.n8559 0.023
R78510 out.n8632 out.n8596 0.023
R78511 out.n8516 out.n8482 0.023
R78512 out.n8555 out.n8519 0.023
R78513 out.n8439 out.n8405 0.023
R78514 out.n8478 out.n8442 0.023
R78515 out.n8362 out.n8328 0.023
R78516 out.n8401 out.n8365 0.023
R78517 out.n8285 out.n8251 0.023
R78518 out.n8324 out.n8288 0.023
R78519 out.n8208 out.n8174 0.023
R78520 out.n8247 out.n8211 0.023
R78521 out.n8131 out.n8097 0.023
R78522 out.n8170 out.n8134 0.023
R78523 out.n8054 out.n8020 0.023
R78524 out.n8093 out.n8057 0.023
R78525 out.n7977 out.n7943 0.023
R78526 out.n8016 out.n7980 0.023
R78527 out.n7900 out.n7866 0.023
R78528 out.n7939 out.n7903 0.023
R78529 out.n7823 out.n5615 0.023
R78530 out.n7862 out.n7826 0.023
R78531 out.n6445 out.n6439 0.023
R78532 out.n2180 out.n1858 0.023
R78533 out.n2180 out.n2070 0.023
R78534 out.n3121 out.n3101 0.023
R78535 out.n3121 out.n3102 0.023
R78536 out.n3057 out.n3051 0.023
R78537 out.n3109 out.n3107 0.023
R78538 out.n3294 out.n3288 0.023
R78539 out.n3238 out.n3227 0.023
R78540 out.n3371 out.n3365 0.023
R78541 out.n3332 out.n3326 0.023
R78542 out.n3448 out.n3442 0.023
R78543 out.n3409 out.n3403 0.023
R78544 out.n3525 out.n3519 0.023
R78545 out.n3486 out.n3480 0.023
R78546 out.n3602 out.n3596 0.023
R78547 out.n3563 out.n3557 0.023
R78548 out.n3679 out.n3673 0.023
R78549 out.n3640 out.n3634 0.023
R78550 out.n3756 out.n3750 0.023
R78551 out.n3717 out.n3711 0.023
R78552 out.n3833 out.n3827 0.023
R78553 out.n3794 out.n3788 0.023
R78554 out.n3910 out.n3904 0.023
R78555 out.n3871 out.n3865 0.023
R78556 out.n907 out.n904 0.023
R78557 out.n3948 out.n3942 0.023
R78558 out.n6767 out.n6204 0.023
R78559 out.n6446 out.n6434 0.023
R78560 out.n2996 out.n2972 0.023
R78561 out.n8732 out.n8721 0.023
R78562 out.n8775 out.n8759 0.023
R78563 out.n8655 out.n8644 0.023
R78564 out.n8692 out.n8681 0.023
R78565 out.n8578 out.n8567 0.023
R78566 out.n8615 out.n8604 0.023
R78567 out.n8501 out.n8490 0.023
R78568 out.n8538 out.n8527 0.023
R78569 out.n8424 out.n8413 0.023
R78570 out.n8461 out.n8450 0.023
R78571 out.n8347 out.n8336 0.023
R78572 out.n8384 out.n8373 0.023
R78573 out.n8270 out.n8259 0.023
R78574 out.n8307 out.n8296 0.023
R78575 out.n8193 out.n8182 0.023
R78576 out.n8230 out.n8219 0.023
R78577 out.n8116 out.n8105 0.023
R78578 out.n8153 out.n8142 0.023
R78579 out.n8039 out.n8028 0.023
R78580 out.n8076 out.n8065 0.023
R78581 out.n7962 out.n7951 0.023
R78582 out.n7999 out.n7988 0.023
R78583 out.n7885 out.n7874 0.023
R78584 out.n7922 out.n7911 0.023
R78585 out.n7845 out.n7834 0.023
R78586 out.n7009 out.n6996 0.023
R78587 out.n2943 out.n2380 0.023
R78588 out.n3070 out.n3058 0.023
R78589 out.n3023 out.n2997 0.023
R78590 out.n3133 out.n3132 0.023
R78591 out.n3150 out.n3124 0.023
R78592 out.n3243 out.n3242 0.023
R78593 out.n3253 out.n3244 0.023
R78594 out.n3307 out.n3295 0.023
R78595 out.n3268 out.n3239 0.023
R78596 out.n3384 out.n3372 0.023
R78597 out.n3345 out.n3333 0.023
R78598 out.n3461 out.n3449 0.023
R78599 out.n3422 out.n3410 0.023
R78600 out.n3538 out.n3526 0.023
R78601 out.n3499 out.n3487 0.023
R78602 out.n3615 out.n3603 0.023
R78603 out.n3576 out.n3564 0.023
R78604 out.n3692 out.n3680 0.023
R78605 out.n3653 out.n3641 0.023
R78606 out.n3769 out.n3757 0.023
R78607 out.n3730 out.n3718 0.023
R78608 out.n3846 out.n3834 0.023
R78609 out.n3807 out.n3795 0.023
R78610 out.n3923 out.n3911 0.023
R78611 out.n3884 out.n3872 0.023
R78612 out.n3984 out.n3973 0.023
R78613 out.n3961 out.n3949 0.023
R78614 out.n8792 out.n8778 0.023
R78615 out.n7465 out.n7242 0.023
R78616 out.n3023 out.n3017 0.023
R78617 out.n3014 out.n3013 0.023
R78618 out.n8792 out.n8787 0.023
R78619 out.n8706 out.n8701 0.023
R78620 out.n8629 out.n8624 0.023
R78621 out.n8552 out.n8547 0.023
R78622 out.n8475 out.n8470 0.023
R78623 out.n8398 out.n8393 0.023
R78624 out.n8321 out.n8316 0.023
R78625 out.n8244 out.n8239 0.023
R78626 out.n8167 out.n8162 0.023
R78627 out.n8090 out.n8085 0.023
R78628 out.n8013 out.n8008 0.023
R78629 out.n7936 out.n7931 0.023
R78630 out.n7859 out.n7854 0.023
R78631 out.n3039 out.n2963 0.023
R78632 out.n2957 out.n1135 0.023
R78633 out.n5862 out.n5857 0.023
R78634 out.n2055 out.n1879 0.023
R78635 out.n10172 out.n10171 0.023
R78636 out.n6185 out.n6182 0.023
R78637 out.n13626 out.n13625 0.023
R78638 out.n14081 out.n14080 0.023
R78639 out.n1596 out.n1595 0.023
R78640 out.n12350 out.n12349 0.023
R78641 out.n11092 out.n11091 0.023
R78642 out.n12792 out.n12791 0.023
R78643 out.n11519 out.n11518 0.023
R78644 out.n14477 out.n14476 0.023
R78645 out.n5151 out.n5150 0.023
R78646 out.n5502 out.n5500 0.023
R78647 out.n7360 out.n7358 0.023
R78648 out.n6179 out.n6178 0.023
R78649 out.n12460 out.n12459 0.023
R78650 out.n13215 out.n13214 0.023
R78651 out.n11930 out.n11929 0.023
R78652 out.n10663 out.n10662 0.023
R78653 out.n2061 out.n2060 0.022
R78654 out.n2932 out.n2931 0.022
R78655 out.n1836 out.n1835 0.022
R78656 out.n2696 out.n2695 0.022
R78657 out.n10879 out.n10877 0.022
R78658 out.n13483 out.n13480 0.022
R78659 out.n13938 out.n13935 0.022
R78660 out.n5746 out.n5744 0.022
R78661 out.n6880 out.n6878 0.022
R78662 out.n12650 out.n12647 0.022
R78663 out.n14492 out.n14491 0.022
R78664 out.n13404 out.n13402 0.022
R78665 out.n13859 out.n13857 0.022
R78666 out.n11309 out.n11307 0.022
R78667 out.n10189 out.n10068 0.022
R78668 out.n10068 out.n10067 0.022
R78669 out.n10131 out.n10090 0.022
R78670 out.n10128 out.n10123 0.022
R78671 out.n13242 out.n13241 0.022
R78672 out.n13113 out.n13112 0.022
R78673 out.n13124 out.n13123 0.022
R78674 out.n13160 out.n13159 0.022
R78675 out.n13171 out.n13170 0.022
R78676 out.n12983 out.n12982 0.022
R78677 out.n12994 out.n12990 0.022
R78678 out.n13014 out.n13013 0.022
R78679 out.n13013 out.n13012 0.022
R78680 out.n13045 out.n13042 0.022
R78681 out.n13062 out.n13061 0.022
R78682 out.n13061 out.n13060 0.022
R78683 out.n12920 out.n12917 0.022
R78684 out.n12806 out.n12410 0.022
R78685 out.n12410 out.n12409 0.022
R78686 out.n12805 out.n12413 0.022
R78687 out.n12692 out.n12691 0.022
R78688 out.n12703 out.n12702 0.022
R78689 out.n12739 out.n12738 0.022
R78690 out.n12750 out.n12749 0.022
R78691 out.n12579 out.n12578 0.022
R78692 out.n12590 out.n12589 0.022
R78693 out.n12621 out.n12618 0.022
R78694 out.n12634 out.n12629 0.022
R78695 out.n12628 out.n12627 0.022
R78696 out.n12639 out.n12638 0.022
R78697 out.n12468 out.n12467 0.022
R78698 out.n12467 out.n12466 0.022
R78699 out.n12496 out.n12493 0.022
R78700 out.n12525 out.n12520 0.022
R78701 out.n12520 out.n12519 0.022
R78702 out.n12519 out.n12518 0.022
R78703 out.n12368 out.n11984 0.022
R78704 out.n12367 out.n11987 0.022
R78705 out.n11987 out.n11986 0.022
R78706 out.n12248 out.n12247 0.022
R78707 out.n12259 out.n12258 0.022
R78708 out.n12295 out.n12294 0.022
R78709 out.n12306 out.n12305 0.022
R78710 out.n12118 out.n12117 0.022
R78711 out.n12129 out.n12125 0.022
R78712 out.n12149 out.n12148 0.022
R78713 out.n12148 out.n12147 0.022
R78714 out.n12180 out.n12177 0.022
R78715 out.n12197 out.n12196 0.022
R78716 out.n12196 out.n12195 0.022
R78717 out.n12027 out.n12026 0.022
R78718 out.n12055 out.n12052 0.022
R78719 out.n13640 out.n13255 0.022
R78720 out.n13255 out.n13254 0.022
R78721 out.n13639 out.n13258 0.022
R78722 out.n13526 out.n13525 0.022
R78723 out.n13537 out.n13536 0.022
R78724 out.n13573 out.n13572 0.022
R78725 out.n13584 out.n13583 0.022
R78726 out.n13412 out.n13411 0.022
R78727 out.n13423 out.n13422 0.022
R78728 out.n13454 out.n13451 0.022
R78729 out.n13467 out.n13462 0.022
R78730 out.n13461 out.n13460 0.022
R78731 out.n13472 out.n13471 0.022
R78732 out.n13301 out.n13300 0.022
R78733 out.n13329 out.n13326 0.022
R78734 out.n13358 out.n13353 0.022
R78735 out.n13353 out.n13352 0.022
R78736 out.n13352 out.n13351 0.022
R78737 out.n11537 out.n11144 0.022
R78738 out.n11536 out.n11147 0.022
R78739 out.n11147 out.n11146 0.022
R78740 out.n11417 out.n11416 0.022
R78741 out.n11428 out.n11427 0.022
R78742 out.n11464 out.n11463 0.022
R78743 out.n11475 out.n11474 0.022
R78744 out.n11295 out.n11294 0.022
R78745 out.n11306 out.n11302 0.022
R78746 out.n11323 out.n11322 0.022
R78747 out.n11322 out.n11321 0.022
R78748 out.n11354 out.n11351 0.022
R78749 out.n11371 out.n11370 0.022
R78750 out.n11370 out.n11369 0.022
R78751 out.n11204 out.n11203 0.022
R78752 out.n11232 out.n11229 0.022
R78753 out.n11110 out.n10721 0.022
R78754 out.n11109 out.n10724 0.022
R78755 out.n10724 out.n10723 0.022
R78756 out.n10990 out.n10989 0.022
R78757 out.n11001 out.n11000 0.022
R78758 out.n11037 out.n11036 0.022
R78759 out.n11048 out.n11047 0.022
R78760 out.n10865 out.n10864 0.022
R78761 out.n10876 out.n10872 0.022
R78762 out.n10896 out.n10895 0.022
R78763 out.n10895 out.n10894 0.022
R78764 out.n10927 out.n10924 0.022
R78765 out.n10944 out.n10943 0.022
R78766 out.n10943 out.n10942 0.022
R78767 out.n10774 out.n10773 0.022
R78768 out.n10802 out.n10799 0.022
R78769 out.n11948 out.n11567 0.022
R78770 out.n11828 out.n11827 0.022
R78771 out.n11839 out.n11838 0.022
R78772 out.n11875 out.n11874 0.022
R78773 out.n11886 out.n11885 0.022
R78774 out.n11698 out.n11697 0.022
R78775 out.n11709 out.n11705 0.022
R78776 out.n11729 out.n11728 0.022
R78777 out.n11728 out.n11727 0.022
R78778 out.n11760 out.n11757 0.022
R78779 out.n11777 out.n11776 0.022
R78780 out.n11776 out.n11775 0.022
R78781 out.n11635 out.n11632 0.022
R78782 out.n14095 out.n13710 0.022
R78783 out.n13710 out.n13709 0.022
R78784 out.n14094 out.n13713 0.022
R78785 out.n13981 out.n13980 0.022
R78786 out.n13992 out.n13991 0.022
R78787 out.n14028 out.n14027 0.022
R78788 out.n14039 out.n14038 0.022
R78789 out.n13867 out.n13866 0.022
R78790 out.n13878 out.n13877 0.022
R78791 out.n13909 out.n13906 0.022
R78792 out.n13922 out.n13917 0.022
R78793 out.n13916 out.n13915 0.022
R78794 out.n13927 out.n13926 0.022
R78795 out.n13756 out.n13755 0.022
R78796 out.n13784 out.n13781 0.022
R78797 out.n13813 out.n13808 0.022
R78798 out.n13808 out.n13807 0.022
R78799 out.n13807 out.n13806 0.022
R78800 out.n10681 out.n10300 0.022
R78801 out.n10561 out.n10560 0.022
R78802 out.n10572 out.n10571 0.022
R78803 out.n10608 out.n10607 0.022
R78804 out.n10619 out.n10618 0.022
R78805 out.n10431 out.n10430 0.022
R78806 out.n10442 out.n10438 0.022
R78807 out.n10462 out.n10461 0.022
R78808 out.n10461 out.n10460 0.022
R78809 out.n10493 out.n10490 0.022
R78810 out.n10510 out.n10509 0.022
R78811 out.n10509 out.n10508 0.022
R78812 out.n10368 out.n10365 0.022
R78813 out.n14550 out.n14187 0.022
R78814 out.n14187 out.n14186 0.022
R78815 out.n14186 out.n14185 0.022
R78816 out.n14269 out.n14268 0.022
R78817 out.n14260 out.n14259 0.022
R78818 out.n14258 out.n14257 0.022
R78819 out.n14251 out.n14250 0.022
R78820 out.n14235 out.n14234 0.022
R78821 out.n14226 out.n14225 0.022
R78822 out.n14338 out.n14337 0.022
R78823 out.n14329 out.n14328 0.022
R78824 out.n14315 out.n14314 0.022
R78825 out.n14306 out.n14305 0.022
R78826 out.n14159 out.n14158 0.022
R78827 out.n14160 out.n14159 0.022
R78828 out.n14391 out.n14388 0.022
R78829 out.n14374 out.n14373 0.022
R78830 out.n14373 out.n14372 0.022
R78831 out.n5025 out.n5024 0.022
R78832 out.n5016 out.n5015 0.022
R78833 out.n5002 out.n5001 0.022
R78834 out.n4993 out.n4992 0.022
R78835 out.n1000 out.n995 0.022
R78836 out.n1009 out.n1006 0.022
R78837 out.n1020 out.n1019 0.022
R78838 out.n1021 out.n1020 0.022
R78839 out.n5080 out.n5077 0.022
R78840 out.n5063 out.n5062 0.022
R78841 out.n5062 out.n5061 0.022
R78842 out.n950 out.n949 0.022
R78843 out.n2736 out.n2735 0.022
R78844 out.n5813 out.n5808 0.022
R78845 out.n5807 out.n5806 0.022
R78846 out.n5791 out.n5788 0.022
R78847 out.n5754 out.n5753 0.022
R78848 out.n5662 out.n5660 0.022
R78849 out.n2878 out.n2877 0.022
R78850 out.n2909 out.n2815 0.022
R78851 out.n2767 out.n2766 0.022
R78852 out.n2785 out.n2784 0.022
R78853 out.n1404 out.n1403 0.022
R78854 out.n1433 out.n1431 0.022
R78855 out.n1463 out.n1462 0.022
R78856 out.n5436 out.n5434 0.022
R78857 out.n5567 out.n5562 0.022
R78858 out.n5562 out.n5561 0.022
R78859 out.n5561 out.n5560 0.022
R78860 out.n5538 out.n5535 0.022
R78861 out.n5510 out.n5509 0.022
R78862 out.n5509 out.n5508 0.022
R78863 out.n5341 out.n5340 0.022
R78864 out.n5334 out.n5331 0.022
R78865 out.n5303 out.n5302 0.022
R78866 out.n5294 out.n5293 0.022
R78867 out.n5208 out.n5205 0.022
R78868 out.n1234 out.n1231 0.022
R78869 out.n1226 out.n1225 0.022
R78870 out.n1207 out.n1206 0.022
R78871 out.n1156 out.n1154 0.022
R78872 out.n1303 out.n1302 0.022
R78873 out.n6538 out.n6534 0.022
R78874 out.n6514 out.n6513 0.022
R78875 out.n6587 out.n6584 0.022
R78876 out.n6603 out.n6601 0.022
R78877 out.n6721 out.n6716 0.022
R78878 out.n6716 out.n6715 0.022
R78879 out.n6715 out.n6714 0.022
R78880 out.n6692 out.n6689 0.022
R78881 out.n6674 out.n6673 0.022
R78882 out.n6673 out.n6672 0.022
R78883 out.n1865 out.n1864 0.022
R78884 out.n6385 out.n6380 0.022
R78885 out.n6379 out.n6378 0.022
R78886 out.n6363 out.n6360 0.022
R78887 out.n6331 out.n6330 0.022
R78888 out.n6239 out.n6237 0.022
R78889 out.n2002 out.n2001 0.022
R78890 out.n2033 out.n1939 0.022
R78891 out.n2047 out.n2046 0.022
R78892 out.n1909 out.n1908 0.022
R78893 out.n6154 out.n6153 0.022
R78894 out.n6153 out.n6152 0.022
R78895 out.n6137 out.n6134 0.022
R78896 out.n6111 out.n6110 0.022
R78897 out.n6110 out.n6109 0.022
R78898 out.n5894 out.n5893 0.022
R78899 out.n6086 out.n6085 0.022
R78900 out.n6017 out.n6014 0.022
R78901 out.n5999 out.n5998 0.022
R78902 out.n5983 out.n5978 0.022
R78903 out.n1586 out.n1585 0.022
R78904 out.n1640 out.n1639 0.022
R78905 out.n6947 out.n6942 0.022
R78906 out.n6941 out.n6940 0.022
R78907 out.n6925 out.n6922 0.022
R78908 out.n6888 out.n6887 0.022
R78909 out.n6796 out.n6794 0.022
R78910 out.n1782 out.n1781 0.022
R78911 out.n1813 out.n1719 0.022
R78912 out.n1671 out.n1670 0.022
R78913 out.n1689 out.n1688 0.022
R78914 out.n2248 out.n2247 0.022
R78915 out.n2277 out.n2275 0.022
R78916 out.n2307 out.n2306 0.022
R78917 out.n7297 out.n7295 0.022
R78918 out.n7425 out.n7420 0.022
R78919 out.n7420 out.n7419 0.022
R78920 out.n7419 out.n7418 0.022
R78921 out.n7396 out.n7393 0.022
R78922 out.n7368 out.n7367 0.022
R78923 out.n7367 out.n7366 0.022
R78924 out.n7175 out.n7172 0.022
R78925 out.n7157 out.n7156 0.022
R78926 out.n7148 out.n7147 0.022
R78927 out.n7122 out.n7117 0.022
R78928 out.n2512 out.n2511 0.022
R78929 out.n2502 out.n2500 0.022
R78930 out.n2488 out.n2486 0.022
R78931 out.n2412 out.n2410 0.022
R78932 out.n2568 out.n2567 0.022
R78933 out.n2626 out.n2625 0.022
R78934 out.n7768 out.n7763 0.022
R78935 out.n7762 out.n7761 0.022
R78936 out.n7746 out.n7743 0.022
R78937 out.n7714 out.n7713 0.022
R78938 out.n7643 out.n7641 0.022
R78939 out.n7530 out.n7527 0.022
R78940 out.n7593 out.n7584 0.022
R78941 out.n2682 out.n2681 0.022
R78942 out.n2648 out.n2647 0.022
R78943 out.n3165 out.n3164 0.022
R78944 out.n3215 out.n3212 0.022
R78945 out.n12571 out.n12569 0.022
R78946 out.n2960 out.n2959 0.022
R78947 out.n2697 out.n2696 0.022
R78948 out.n2075 out.n2074 0.021
R78949 out.n2171 out.n2170 0.021
R78950 out.n2990 out.n2989 0.021
R78951 out.n3232 out.n3231 0.021
R78952 out.n8773 out.n8772 0.021
R78953 out.n6765 out.n6764 0.021
R78954 out.n16268 out.n16267 0.021
R78955 out.n15166 out.n15165 0.021
R78956 out.n1597 out.n1596 0.021
R78957 out.n15432 out.n15431 0.021
R78958 out.n7461 out.n7460 0.021
R78959 out.n5603 out.n5602 0.021
R78960 out.n14549 out.n14548 0.021
R78961 out.n15941 out.n15371 0.021
R78962 out.n14131 out.n14130 0.021
R78963 out.n15446 out.n15445 0.021
R78964 out.n15346 out.n15344 0.021
R78965 out.n9000 out.n8998 0.021
R78966 out.n15281 out.n15279 0.021
R78967 out.n15314 out.n15312 0.021
R78968 out.n15216 out.n15214 0.021
R78969 out.n15249 out.n15247 0.021
R78970 out.n8950 out.n8948 0.021
R78971 out.n15183 out.n15181 0.021
R78972 out.n8913 out.n8911 0.021
R78973 out.n15143 out.n15141 0.021
R78974 out.n15073 out.n15071 0.021
R78975 out.n15105 out.n15103 0.021
R78976 out.n15008 out.n15006 0.021
R78977 out.n15040 out.n15038 0.021
R78978 out.n14940 out.n14938 0.021
R78979 out.n14975 out.n14973 0.021
R78980 out.n14869 out.n14867 0.021
R78981 out.n14904 out.n14902 0.021
R78982 out.n14798 out.n14796 0.021
R78983 out.n14833 out.n14831 0.021
R78984 out.n14727 out.n14725 0.021
R78985 out.n14762 out.n14760 0.021
R78986 out.n14656 out.n14654 0.021
R78987 out.n14691 out.n14689 0.021
R78988 out.n14583 out.n14581 0.021
R78989 out.n14620 out.n14618 0.021
R78990 out.n903 out.n902 0.021
R78991 out.n8724 out.n8723 0.021
R78992 out.n8763 out.n8762 0.021
R78993 out.n8647 out.n8646 0.021
R78994 out.n8684 out.n8683 0.021
R78995 out.n8570 out.n8569 0.021
R78996 out.n8607 out.n8606 0.021
R78997 out.n8493 out.n8492 0.021
R78998 out.n8530 out.n8529 0.021
R78999 out.n8416 out.n8415 0.021
R79000 out.n8453 out.n8452 0.021
R79001 out.n8339 out.n8338 0.021
R79002 out.n8376 out.n8375 0.021
R79003 out.n8262 out.n8261 0.021
R79004 out.n8299 out.n8298 0.021
R79005 out.n8185 out.n8184 0.021
R79006 out.n8222 out.n8221 0.021
R79007 out.n8108 out.n8107 0.021
R79008 out.n8145 out.n8144 0.021
R79009 out.n8031 out.n8030 0.021
R79010 out.n8068 out.n8067 0.021
R79011 out.n7954 out.n7953 0.021
R79012 out.n7991 out.n7990 0.021
R79013 out.n7877 out.n7876 0.021
R79014 out.n7914 out.n7913 0.021
R79015 out.n7837 out.n7836 0.021
R79016 out.n1857 out.n1853 0.021
R79017 out.n1852 out.n1845 0.021
R79018 out.n2984 out.n2977 0.021
R79019 out.n3048 out.n3047 0.021
R79020 out.n3100 out.n3094 0.021
R79021 out.n3093 out.n3092 0.021
R79022 out.n3218 out.n3216 0.021
R79023 out.n3224 out.n3208 0.021
R79024 out.n3285 out.n3284 0.021
R79025 out.n3323 out.n3322 0.021
R79026 out.n3362 out.n3361 0.021
R79027 out.n3400 out.n3399 0.021
R79028 out.n3439 out.n3438 0.021
R79029 out.n3477 out.n3476 0.021
R79030 out.n3516 out.n3515 0.021
R79031 out.n3554 out.n3553 0.021
R79032 out.n3593 out.n3592 0.021
R79033 out.n3631 out.n3630 0.021
R79034 out.n3670 out.n3669 0.021
R79035 out.n3708 out.n3707 0.021
R79036 out.n3747 out.n3746 0.021
R79037 out.n3785 out.n3784 0.021
R79038 out.n3824 out.n3823 0.021
R79039 out.n3862 out.n3861 0.021
R79040 out.n3901 out.n3900 0.021
R79041 out.n3939 out.n3938 0.021
R79042 out.n901 out.n900 0.021
R79043 out.n8761 out.n8760 0.021
R79044 out.n6203 out.n6199 0.021
R79045 out.n10709 out.n10708 0.021
R79046 out.n14117 out.n14116 0.021
R79047 out.n14112 out.n14111 0.021
R79048 out.n14602 out.n14601 0.021
R79049 out.n14639 out.n14638 0.021
R79050 out.n14673 out.n14672 0.021
R79051 out.n14710 out.n14709 0.021
R79052 out.n14744 out.n14743 0.021
R79053 out.n14781 out.n14780 0.021
R79054 out.n14815 out.n14814 0.021
R79055 out.n14852 out.n14851 0.021
R79056 out.n14886 out.n14885 0.021
R79057 out.n14923 out.n14922 0.021
R79058 out.n14957 out.n14956 0.021
R79059 out.n14994 out.n14993 0.021
R79060 out.n15025 out.n15024 0.021
R79061 out.n15059 out.n15058 0.021
R79062 out.n15090 out.n15089 0.021
R79063 out.n8899 out.n8898 0.021
R79064 out.n15128 out.n15127 0.021
R79065 out.n8936 out.n8935 0.021
R79066 out.n15168 out.n15167 0.021
R79067 out.n15202 out.n15201 0.021
R79068 out.n15234 out.n15233 0.021
R79069 out.n15267 out.n15266 0.021
R79070 out.n15299 out.n15298 0.021
R79071 out.n15332 out.n15331 0.021
R79072 out.n8984 out.n8983 0.021
R79073 out.n15396 out.n15394 0.021
R79074 out.n15444 out.n15443 0.021
R79075 out.n15348 out.n15347 0.021
R79076 out.n9002 out.n9001 0.021
R79077 out.n15283 out.n15282 0.021
R79078 out.n15316 out.n15315 0.021
R79079 out.n15218 out.n15217 0.021
R79080 out.n15251 out.n15250 0.021
R79081 out.n8952 out.n8951 0.021
R79082 out.n15185 out.n15184 0.021
R79083 out.n8915 out.n8914 0.021
R79084 out.n15145 out.n15144 0.021
R79085 out.n15075 out.n15074 0.021
R79086 out.n15107 out.n15106 0.021
R79087 out.n15010 out.n15009 0.021
R79088 out.n15042 out.n15041 0.021
R79089 out.n14942 out.n14941 0.021
R79090 out.n14977 out.n14976 0.021
R79091 out.n14871 out.n14870 0.021
R79092 out.n14906 out.n14905 0.021
R79093 out.n14800 out.n14799 0.021
R79094 out.n14835 out.n14834 0.021
R79095 out.n14729 out.n14728 0.021
R79096 out.n14764 out.n14763 0.021
R79097 out.n14658 out.n14657 0.021
R79098 out.n14693 out.n14692 0.021
R79099 out.n14585 out.n14584 0.021
R79100 out.n14622 out.n14621 0.021
R79101 out.n14134 out.n14133 0.021
R79102 out.n15482 out.n15481 0.021
R79103 out.n15448 out.n15447 0.021
R79104 out.n15550 out.n15549 0.021
R79105 out.n15518 out.n15517 0.021
R79106 out.n15631 out.n15630 0.021
R79107 out.n15595 out.n15594 0.021
R79108 out.n15703 out.n15702 0.021
R79109 out.n15666 out.n15665 0.021
R79110 out.n15769 out.n15768 0.021
R79111 out.n15737 out.n15736 0.021
R79112 out.n15830 out.n15829 0.021
R79113 out.n15798 out.n15797 0.021
R79114 out.n15891 out.n15890 0.021
R79115 out.n15859 out.n15858 0.021
R79116 out.n15927 out.n15926 0.021
R79117 out.n16004 out.n16003 0.021
R79118 out.n16065 out.n16064 0.021
R79119 out.n15968 out.n15967 0.021
R79120 out.n16127 out.n16126 0.021
R79121 out.n16095 out.n16094 0.021
R79122 out.n16188 out.n16187 0.021
R79123 out.n16156 out.n16155 0.021
R79124 out.n16223 out.n16222 0.021
R79125 out.n17267 out.n17266 0.021
R79126 out.n16253 out.n16252 0.021
R79127 out.n15513 out.n15512 0.021
R79128 out.n15545 out.n15544 0.021
R79129 out.n15586 out.n15585 0.021
R79130 out.n15626 out.n15625 0.021
R79131 out.n15661 out.n15660 0.021
R79132 out.n15698 out.n15697 0.021
R79133 out.n15732 out.n15731 0.021
R79134 out.n15764 out.n15763 0.021
R79135 out.n15793 out.n15792 0.021
R79136 out.n15825 out.n15824 0.021
R79137 out.n15854 out.n15853 0.021
R79138 out.n15886 out.n15885 0.021
R79139 out.n15995 out.n15994 0.021
R79140 out.n15922 out.n15921 0.021
R79141 out.n15959 out.n15958 0.021
R79142 out.n16060 out.n16059 0.021
R79143 out.n16090 out.n16089 0.021
R79144 out.n16122 out.n16121 0.021
R79145 out.n16151 out.n16150 0.021
R79146 out.n16183 out.n16182 0.021
R79147 out.n17258 out.n17257 0.021
R79148 out.n16218 out.n16217 0.021
R79149 out.n16248 out.n16247 0.021
R79150 out.n12397 out.n12394 0.021
R79151 out.n12827 out.n12824 0.021
R79152 out.n15487 out.n15485 0.021
R79153 out.n15523 out.n15521 0.021
R79154 out.n15554 out.n15553 0.021
R79155 out.n15600 out.n15598 0.021
R79156 out.n15635 out.n15634 0.021
R79157 out.n15671 out.n15669 0.021
R79158 out.n15707 out.n15706 0.021
R79159 out.n15742 out.n15740 0.021
R79160 out.n15773 out.n15772 0.021
R79161 out.n15803 out.n15801 0.021
R79162 out.n15834 out.n15833 0.021
R79163 out.n15864 out.n15862 0.021
R79164 out.n15895 out.n15894 0.021
R79165 out.n16009 out.n16007 0.021
R79166 out.n15931 out.n15930 0.021
R79167 out.n15973 out.n15971 0.021
R79168 out.n16069 out.n16068 0.021
R79169 out.n16100 out.n16098 0.021
R79170 out.n16131 out.n16130 0.021
R79171 out.n16161 out.n16159 0.021
R79172 out.n16192 out.n16191 0.021
R79173 out.n17272 out.n17270 0.021
R79174 out.n16227 out.n16226 0.021
R79175 out.n16258 out.n16256 0.021
R79176 out.n9009 out.n9008 0.021
R79177 out.n15354 out.n15353 0.021
R79178 out.n15322 out.n15321 0.021
R79179 out.n15289 out.n15288 0.021
R79180 out.n15257 out.n15256 0.021
R79181 out.n15224 out.n15223 0.021
R79182 out.n15192 out.n15191 0.021
R79183 out.n8959 out.n8958 0.021
R79184 out.n15151 out.n15150 0.021
R79185 out.n8924 out.n8923 0.021
R79186 out.n15113 out.n15112 0.021
R79187 out.n15081 out.n15080 0.021
R79188 out.n15048 out.n15047 0.021
R79189 out.n15016 out.n15015 0.021
R79190 out.n14983 out.n14982 0.021
R79191 out.n14948 out.n14947 0.021
R79192 out.n14912 out.n14911 0.021
R79193 out.n14877 out.n14876 0.021
R79194 out.n14841 out.n14840 0.021
R79195 out.n14806 out.n14805 0.021
R79196 out.n14770 out.n14769 0.021
R79197 out.n14735 out.n14734 0.021
R79198 out.n14699 out.n14698 0.021
R79199 out.n14664 out.n14663 0.021
R79200 out.n14628 out.n14627 0.021
R79201 out.n14593 out.n14592 0.021
R79202 out.n14141 out.n14139 0.021
R79203 out.n13674 out.n13671 0.021
R79204 out.n14579 out.n14578 0.021
R79205 out.n14652 out.n14651 0.021
R79206 out.n14723 out.n14722 0.021
R79207 out.n14794 out.n14793 0.021
R79208 out.n14865 out.n14864 0.021
R79209 out.n14936 out.n14935 0.021
R79210 out.n15004 out.n15003 0.021
R79211 out.n15069 out.n15068 0.021
R79212 out.n8909 out.n8908 0.021
R79213 out.n8946 out.n8945 0.021
R79214 out.n15212 out.n15211 0.021
R79215 out.n15277 out.n15276 0.021
R79216 out.n15342 out.n15341 0.021
R79217 out.n16240 out.n16239 0.021
R79218 out.n16210 out.n16209 0.021
R79219 out.n17250 out.n17249 0.021
R79220 out.n16175 out.n16174 0.021
R79221 out.n16143 out.n16142 0.021
R79222 out.n16114 out.n16113 0.021
R79223 out.n16082 out.n16081 0.021
R79224 out.n16052 out.n16051 0.021
R79225 out.n15951 out.n15950 0.021
R79226 out.n15914 out.n15913 0.021
R79227 out.n15987 out.n15986 0.021
R79228 out.n15878 out.n15877 0.021
R79229 out.n15846 out.n15845 0.021
R79230 out.n15817 out.n15816 0.021
R79231 out.n15785 out.n15784 0.021
R79232 out.n15756 out.n15755 0.021
R79233 out.n15724 out.n15723 0.021
R79234 out.n15690 out.n15689 0.021
R79235 out.n15653 out.n15652 0.021
R79236 out.n15618 out.n15617 0.021
R79237 out.n15578 out.n15577 0.021
R79238 out.n15537 out.n15536 0.021
R79239 out.n15505 out.n15504 0.021
R79240 out.n15470 out.n15469 0.021
R79241 out.n14122 out.n14121 0.021
R79242 out.n14610 out.n14609 0.021
R79243 out.n14681 out.n14680 0.021
R79244 out.n14752 out.n14751 0.021
R79245 out.n14823 out.n14822 0.021
R79246 out.n14894 out.n14893 0.021
R79247 out.n14965 out.n14964 0.021
R79248 out.n15030 out.n15029 0.021
R79249 out.n15095 out.n15094 0.021
R79250 out.n15133 out.n15132 0.021
R79251 out.n15173 out.n15172 0.021
R79252 out.n15239 out.n15238 0.021
R79253 out.n15304 out.n15303 0.021
R79254 out.n8990 out.n8989 0.021
R79255 out.n16213 out.n16212 0.021
R79256 out.n16178 out.n16177 0.021
R79257 out.n16117 out.n16116 0.021
R79258 out.n16055 out.n16054 0.021
R79259 out.n15917 out.n15916 0.021
R79260 out.n15881 out.n15880 0.021
R79261 out.n15820 out.n15819 0.021
R79262 out.n15759 out.n15758 0.021
R79263 out.n15693 out.n15692 0.021
R79264 out.n15621 out.n15620 0.021
R79265 out.n15540 out.n15539 0.021
R79266 out.n15473 out.n15472 0.021
R79267 out.n15442 out.n15441 0.021
R79268 out.n11136 out.n11133 0.021
R79269 out.n15435 out.n15434 0.021
R79270 out.n15337 out.n15336 0.021
R79271 out.n15272 out.n15271 0.021
R79272 out.n15207 out.n15206 0.021
R79273 out.n8941 out.n8940 0.021
R79274 out.n8904 out.n8903 0.021
R79275 out.n15064 out.n15063 0.021
R79276 out.n14999 out.n14998 0.021
R79277 out.n14931 out.n14930 0.021
R79278 out.n14860 out.n14859 0.021
R79279 out.n14789 out.n14788 0.021
R79280 out.n14718 out.n14717 0.021
R79281 out.n14647 out.n14646 0.021
R79282 out.n14574 out.n14573 0.021
R79283 out.n15491 out.n15490 0.021
R79284 out.n15527 out.n15526 0.021
R79285 out.n15557 out.n15556 0.021
R79286 out.n15604 out.n15603 0.021
R79287 out.n15638 out.n15637 0.021
R79288 out.n15675 out.n15674 0.021
R79289 out.n15710 out.n15709 0.021
R79290 out.n15746 out.n15745 0.021
R79291 out.n15776 out.n15775 0.021
R79292 out.n15807 out.n15806 0.021
R79293 out.n15837 out.n15836 0.021
R79294 out.n15868 out.n15867 0.021
R79295 out.n15898 out.n15897 0.021
R79296 out.n16013 out.n16012 0.021
R79297 out.n15934 out.n15933 0.021
R79298 out.n15977 out.n15976 0.021
R79299 out.n16072 out.n16071 0.021
R79300 out.n16104 out.n16103 0.021
R79301 out.n16134 out.n16133 0.021
R79302 out.n16165 out.n16164 0.021
R79303 out.n16195 out.n16194 0.021
R79304 out.n17276 out.n17275 0.021
R79305 out.n16230 out.n16229 0.021
R79306 out.n16262 out.n16261 0.021
R79307 out.n9013 out.n9011 0.021
R79308 out.n15357 out.n15356 0.021
R79309 out.n15326 out.n15324 0.021
R79310 out.n15292 out.n15291 0.021
R79311 out.n15261 out.n15259 0.021
R79312 out.n15227 out.n15226 0.021
R79313 out.n15196 out.n15194 0.021
R79314 out.n8962 out.n8961 0.021
R79315 out.n15155 out.n15153 0.021
R79316 out.n8927 out.n8926 0.021
R79317 out.n15117 out.n15115 0.021
R79318 out.n15084 out.n15083 0.021
R79319 out.n15052 out.n15050 0.021
R79320 out.n15019 out.n15018 0.021
R79321 out.n14987 out.n14985 0.021
R79322 out.n14951 out.n14950 0.021
R79323 out.n14916 out.n14914 0.021
R79324 out.n14880 out.n14879 0.021
R79325 out.n14845 out.n14843 0.021
R79326 out.n14809 out.n14808 0.021
R79327 out.n14774 out.n14772 0.021
R79328 out.n14738 out.n14737 0.021
R79329 out.n14703 out.n14701 0.021
R79330 out.n14667 out.n14666 0.021
R79331 out.n14632 out.n14630 0.021
R79332 out.n14596 out.n14595 0.021
R79333 out.n14145 out.n14143 0.021
R79334 out.n14101 out.n14098 0.021
R79335 out.n7857 out.n7856 0.021
R79336 out.n7934 out.n7933 0.021
R79337 out.n8011 out.n8010 0.021
R79338 out.n8088 out.n8087 0.021
R79339 out.n8165 out.n8164 0.021
R79340 out.n8242 out.n8241 0.021
R79341 out.n8319 out.n8318 0.021
R79342 out.n8396 out.n8395 0.021
R79343 out.n8473 out.n8472 0.021
R79344 out.n8550 out.n8549 0.021
R79345 out.n8627 out.n8626 0.021
R79346 out.n8704 out.n8703 0.021
R79347 out.n8791 out.n8790 0.021
R79348 out.n3960 out.n3959 0.021
R79349 out.n3883 out.n3882 0.021
R79350 out.n3806 out.n3805 0.021
R79351 out.n3729 out.n3728 0.021
R79352 out.n3652 out.n3651 0.021
R79353 out.n3575 out.n3574 0.021
R79354 out.n3498 out.n3497 0.021
R79355 out.n3421 out.n3420 0.021
R79356 out.n3344 out.n3343 0.021
R79357 out.n3267 out.n3266 0.021
R79358 out.n3069 out.n3068 0.021
R79359 out.n3022 out.n3021 0.021
R79360 out.n2942 out.n2941 0.021
R79361 out.n2971 out.n2966 0.021
R79362 out.n8767 out.n8766 0.021
R79363 out.n8765 out.n8764 0.021
R79364 out.n8726 out.n8725 0.021
R79365 out.n8686 out.n8685 0.021
R79366 out.n8649 out.n8648 0.021
R79367 out.n8609 out.n8608 0.021
R79368 out.n8572 out.n8571 0.021
R79369 out.n8532 out.n8531 0.021
R79370 out.n8495 out.n8494 0.021
R79371 out.n8455 out.n8454 0.021
R79372 out.n8418 out.n8417 0.021
R79373 out.n8378 out.n8377 0.021
R79374 out.n8341 out.n8340 0.021
R79375 out.n8301 out.n8300 0.021
R79376 out.n8264 out.n8263 0.021
R79377 out.n8224 out.n8223 0.021
R79378 out.n8187 out.n8186 0.021
R79379 out.n8147 out.n8146 0.021
R79380 out.n8110 out.n8109 0.021
R79381 out.n8070 out.n8069 0.021
R79382 out.n8033 out.n8032 0.021
R79383 out.n7993 out.n7992 0.021
R79384 out.n7956 out.n7955 0.021
R79385 out.n7916 out.n7915 0.021
R79386 out.n7879 out.n7878 0.021
R79387 out.n7839 out.n7838 0.021
R79388 out.n1620 out.n1613 0.021
R79389 out.n1626 out.n1622 0.021
R79390 out.n3083 out.n3082 0.021
R79391 out.n3044 out.n3043 0.021
R79392 out.n3089 out.n3087 0.021
R79393 out.n3281 out.n3280 0.021
R79394 out.n3203 out.n3202 0.021
R79395 out.n3358 out.n3357 0.021
R79396 out.n3319 out.n3318 0.021
R79397 out.n3435 out.n3434 0.021
R79398 out.n3396 out.n3395 0.021
R79399 out.n3512 out.n3511 0.021
R79400 out.n3473 out.n3472 0.021
R79401 out.n3589 out.n3588 0.021
R79402 out.n3550 out.n3549 0.021
R79403 out.n3666 out.n3665 0.021
R79404 out.n3627 out.n3626 0.021
R79405 out.n3743 out.n3742 0.021
R79406 out.n3704 out.n3703 0.021
R79407 out.n3820 out.n3819 0.021
R79408 out.n3781 out.n3780 0.021
R79409 out.n3897 out.n3896 0.021
R79410 out.n3858 out.n3857 0.021
R79411 out.n897 out.n896 0.021
R79412 out.n3935 out.n3934 0.021
R79413 out.n6197 out.n6194 0.021
R79414 out.n2387 out.n2383 0.021
R79415 out.n3127 out.n3125 0.021
R79416 out.n8780 out.n8779 0.021
R79417 out.n8736 out.n8735 0.021
R79418 out.n8696 out.n8695 0.021
R79419 out.n8659 out.n8658 0.021
R79420 out.n8619 out.n8618 0.021
R79421 out.n8582 out.n8581 0.021
R79422 out.n8542 out.n8541 0.021
R79423 out.n8505 out.n8504 0.021
R79424 out.n8465 out.n8464 0.021
R79425 out.n8428 out.n8427 0.021
R79426 out.n8388 out.n8387 0.021
R79427 out.n8351 out.n8350 0.021
R79428 out.n8311 out.n8310 0.021
R79429 out.n8274 out.n8273 0.021
R79430 out.n8234 out.n8233 0.021
R79431 out.n8197 out.n8196 0.021
R79432 out.n8157 out.n8156 0.021
R79433 out.n8120 out.n8119 0.021
R79434 out.n8080 out.n8079 0.021
R79435 out.n8043 out.n8042 0.021
R79436 out.n8003 out.n8002 0.021
R79437 out.n7966 out.n7965 0.021
R79438 out.n7926 out.n7925 0.021
R79439 out.n7889 out.n7888 0.021
R79440 out.n7849 out.n7848 0.021
R79441 out.n7468 out.n7016 0.021
R79442 out.n2606 out.n2605 0.021
R79443 out.n2600 out.n2593 0.021
R79444 out.n3061 out.n3060 0.021
R79445 out.n3006 out.n2999 0.021
R79446 out.n3138 out.n3137 0.021
R79447 out.n3129 out.n3128 0.021
R79448 out.n3250 out.n3249 0.021
R79449 out.n3255 out.n3241 0.021
R79450 out.n3336 out.n3335 0.021
R79451 out.n3298 out.n3297 0.021
R79452 out.n3413 out.n3412 0.021
R79453 out.n3375 out.n3374 0.021
R79454 out.n3490 out.n3489 0.021
R79455 out.n3452 out.n3451 0.021
R79456 out.n3567 out.n3566 0.021
R79457 out.n3529 out.n3528 0.021
R79458 out.n3644 out.n3643 0.021
R79459 out.n3606 out.n3605 0.021
R79460 out.n3721 out.n3720 0.021
R79461 out.n3683 out.n3682 0.021
R79462 out.n3798 out.n3797 0.021
R79463 out.n3760 out.n3759 0.021
R79464 out.n3875 out.n3874 0.021
R79465 out.n3837 out.n3836 0.021
R79466 out.n3952 out.n3951 0.021
R79467 out.n3914 out.n3913 0.021
R79468 out.n3975 out.n3974 0.021
R79469 out.n8739 out.n8738 0.021
R79470 out.n8785 out.n8784 0.021
R79471 out.n8782 out.n8781 0.021
R79472 out.n8662 out.n8661 0.021
R79473 out.n8700 out.n8699 0.021
R79474 out.n8585 out.n8584 0.021
R79475 out.n8623 out.n8622 0.021
R79476 out.n8508 out.n8507 0.021
R79477 out.n8546 out.n8545 0.021
R79478 out.n8431 out.n8430 0.021
R79479 out.n8469 out.n8468 0.021
R79480 out.n8354 out.n8353 0.021
R79481 out.n8392 out.n8391 0.021
R79482 out.n8277 out.n8276 0.021
R79483 out.n8315 out.n8314 0.021
R79484 out.n8200 out.n8199 0.021
R79485 out.n8238 out.n8237 0.021
R79486 out.n8123 out.n8122 0.021
R79487 out.n8161 out.n8160 0.021
R79488 out.n8046 out.n8045 0.021
R79489 out.n8084 out.n8083 0.021
R79490 out.n7969 out.n7968 0.021
R79491 out.n8007 out.n8006 0.021
R79492 out.n7892 out.n7891 0.021
R79493 out.n7930 out.n7929 0.021
R79494 out.n7474 out.n7473 0.021
R79495 out.n7853 out.n7852 0.021
R79496 out.n2723 out.n2722 0.021
R79497 out.n2715 out.n2714 0.021
R79498 out.n3147 out.n3146 0.021
R79499 out.n3149 out.n3148 0.021
R79500 out.n3066 out.n3065 0.021
R79501 out.n3306 out.n3305 0.021
R79502 out.n3263 out.n3261 0.021
R79503 out.n3383 out.n3382 0.021
R79504 out.n3341 out.n3340 0.021
R79505 out.n3460 out.n3459 0.021
R79506 out.n3418 out.n3417 0.021
R79507 out.n3537 out.n3536 0.021
R79508 out.n3495 out.n3494 0.021
R79509 out.n3614 out.n3613 0.021
R79510 out.n3572 out.n3571 0.021
R79511 out.n3691 out.n3690 0.021
R79512 out.n3649 out.n3648 0.021
R79513 out.n3768 out.n3767 0.021
R79514 out.n3726 out.n3725 0.021
R79515 out.n3845 out.n3844 0.021
R79516 out.n3803 out.n3802 0.021
R79517 out.n3922 out.n3921 0.021
R79518 out.n3880 out.n3879 0.021
R79519 out.n3983 out.n3982 0.021
R79520 out.n3957 out.n3956 0.021
R79521 out.n8789 out.n8788 0.021
R79522 out.n8742 out.n8741 0.021
R79523 out.n8665 out.n8664 0.021
R79524 out.n8588 out.n8587 0.021
R79525 out.n8511 out.n8510 0.021
R79526 out.n8434 out.n8433 0.021
R79527 out.n8357 out.n8356 0.021
R79528 out.n8280 out.n8279 0.021
R79529 out.n8203 out.n8202 0.021
R79530 out.n8126 out.n8125 0.021
R79531 out.n8049 out.n8048 0.021
R79532 out.n7972 out.n7971 0.021
R79533 out.n7895 out.n7894 0.021
R79534 out.n7818 out.n7817 0.021
R79535 out.n14576 out.n14575 0.021
R79536 out.n14649 out.n14648 0.021
R79537 out.n14720 out.n14719 0.021
R79538 out.n14791 out.n14790 0.021
R79539 out.n14862 out.n14861 0.021
R79540 out.n14933 out.n14932 0.021
R79541 out.n15001 out.n15000 0.021
R79542 out.n15066 out.n15065 0.021
R79543 out.n8906 out.n8905 0.021
R79544 out.n8943 out.n8942 0.021
R79545 out.n15209 out.n15208 0.021
R79546 out.n15274 out.n15273 0.021
R79547 out.n15339 out.n15338 0.021
R79548 out.n16245 out.n16244 0.021
R79549 out.n17255 out.n17254 0.021
R79550 out.n16148 out.n16147 0.021
R79551 out.n16087 out.n16086 0.021
R79552 out.n15956 out.n15955 0.021
R79553 out.n15992 out.n15991 0.021
R79554 out.n15851 out.n15850 0.021
R79555 out.n15790 out.n15789 0.021
R79556 out.n15729 out.n15728 0.021
R79557 out.n15658 out.n15657 0.021
R79558 out.n15583 out.n15582 0.021
R79559 out.n15510 out.n15509 0.021
R79560 out.n15438 out.n15437 0.021
R79561 out.n15476 out.n15475 0.021
R79562 out.n15543 out.n15542 0.021
R79563 out.n15624 out.n15623 0.021
R79564 out.n15696 out.n15695 0.021
R79565 out.n15762 out.n15761 0.021
R79566 out.n15823 out.n15822 0.021
R79567 out.n15884 out.n15883 0.021
R79568 out.n15920 out.n15919 0.021
R79569 out.n16058 out.n16057 0.021
R79570 out.n16120 out.n16119 0.021
R79571 out.n16181 out.n16180 0.021
R79572 out.n16216 out.n16215 0.021
R79573 out.n8995 out.n8994 0.021
R79574 out.n15308 out.n15307 0.021
R79575 out.n15243 out.n15242 0.021
R79576 out.n15177 out.n15176 0.021
R79577 out.n15137 out.n15136 0.021
R79578 out.n15099 out.n15098 0.021
R79579 out.n15034 out.n15033 0.021
R79580 out.n14969 out.n14968 0.021
R79581 out.n14898 out.n14897 0.021
R79582 out.n14827 out.n14826 0.021
R79583 out.n14756 out.n14755 0.021
R79584 out.n14685 out.n14684 0.021
R79585 out.n14614 out.n14613 0.021
R79586 out.n14126 out.n14125 0.021
R79587 out.n11559 out.n11556 0.021
R79588 out.n2056 out.n2055 0.021
R79589 out.n6164 out.n6161 0.021
R79590 out.n2579 out.n2578 0.02
R79591 out.n2883 out.n2874 0.02
R79592 out.n1787 out.n1778 0.02
R79593 out.n11381 out.n11378 0.02
R79594 out.n6726 out.n6723 0.02
R79595 out.n10954 out.n10951 0.02
R79596 out.n14416 out.n14415 0.02
R79597 out.n5090 out.n5089 0.02
R79598 out.n2927 out.n2926 0.02
R79599 out.n1831 out.n1830 0.02
R79600 out.n6560 out.n6558 0.02
R79601 out.n1472 out.n1459 0.02
R79602 out.n2319 out.n2303 0.02
R79603 out.n5572 out.n5569 0.02
R79604 out.n7430 out.n7427 0.02
R79605 out.n2921 out.n2768 0.02
R79606 out.n1470 out.n1464 0.02
R79607 out.n1825 out.n1672 0.02
R79608 out.n2317 out.n2308 0.02
R79609 out.n13072 out.n13069 0.02
R79610 out.n11787 out.n11784 0.02
R79611 out.n10520 out.n10517 0.02
R79612 out.n12207 out.n12204 0.02
R79613 out.n14505 out.n14503 0.02
R79614 out.n2007 out.n1998 0.02
R79615 out.n2686 out.n2685 0.02
R79616 out.n2881 out.n2879 0.02
R79617 out.n1785 out.n1783 0.02
R79618 out.n5610 out.n5608 0.02
R79619 out.n3026 out.n3025 0.02
R79620 out.n3028 out.n3027 0.02
R79621 out.n3001 out.n3000 0.02
R79622 out.n3004 out.n3002 0.02
R79623 out.n7466 out.n7017 0.02
R79624 out.n7732 out.n7730 0.02
R79625 out.n1094 out.n1092 0.02
R79626 out.n1313 out.n1311 0.02
R79627 out.n13361 out.n13360 0.02
R79628 out.n13816 out.n13815 0.02
R79629 out.n1306 out.n1304 0.02
R79630 out.n2050 out.n2048 0.02
R79631 out.n14458 out.n14457 0.02
R79632 out.n5132 out.n5131 0.02
R79633 out.n7169 out.n7168 0.02
R79634 out.n2963 out.n2962 0.02
R79635 out.n14508 out.n14506 0.02
R79636 out.n14451 out.n14450 0.02
R79637 out.n14449 out.n14447 0.02
R79638 out.n14396 out.n14395 0.02
R79639 out.n5125 out.n5124 0.02
R79640 out.n5123 out.n5121 0.02
R79641 out.n1046 out.n1044 0.02
R79642 out.n1101 out.n1099 0.02
R79643 out.n1247 out.n1245 0.02
R79644 out.n6350 out.n6349 0.02
R79645 out.n1323 out.n1322 0.02
R79646 out.n12528 out.n12527 0.02
R79647 out.n2005 out.n2003 0.02
R79648 out.n14443 out.n14441 0.02
R79649 out.n14403 out.n14402 0.02
R79650 out.n5117 out.n5115 0.02
R79651 out.n1039 out.n1037 0.02
R79652 out.n2522 out.n2520 0.02
R79653 out.n1087 out.n1085 0.02
R79654 out.n2515 out.n2513 0.02
R79655 out.n2571 out.n2569 0.02
R79656 out.n7167 out.n7166 0.02
R79657 out.n2153 out.n2151 0.019
R79658 out.n14498 out.n14252 0.019
R79659 out.n2919 out.n2773 0.019
R79660 out.n1468 out.n1466 0.019
R79661 out.n1823 out.n1677 0.019
R79662 out.n2315 out.n2313 0.019
R79663 out.n7614 out.n7612 0.019
R79664 out.n7799 out.n7797 0.019
R79665 out.n6192 out.n5868 0.019
R79666 out.n6568 out.n6566 0.019
R79667 out.n8868 out.n8867 0.019
R79668 out.n8862 out.n8861 0.019
R79669 out.n8865 out.n8864 0.019
R79670 out.n8856 out.n8855 0.019
R79671 out.n8859 out.n8858 0.019
R79672 out.n8850 out.n8849 0.019
R79673 out.n8853 out.n8852 0.019
R79674 out.n8841 out.n8840 0.019
R79675 out.n8835 out.n8834 0.019
R79676 out.n8838 out.n8837 0.019
R79677 out.n8829 out.n8828 0.019
R79678 out.n8832 out.n8831 0.019
R79679 out.n8824 out.n8823 0.019
R79680 out.n8821 out.n8820 0.019
R79681 out.n8813 out.n8812 0.019
R79682 out.n8816 out.n8815 0.019
R79683 out.n8807 out.n8806 0.019
R79684 out.n8810 out.n8809 0.019
R79685 out.n8801 out.n8800 0.019
R79686 out.n8804 out.n8803 0.019
R79687 out.n4908 out.n4907 0.019
R79688 out.n8798 out.n8797 0.019
R79689 out.n4898 out.n4897 0.019
R79690 out.n4901 out.n4900 0.019
R79691 out.n4892 out.n4891 0.019
R79692 out.n4895 out.n4894 0.019
R79693 out.n4885 out.n4884 0.019
R79694 out.n4877 out.n4876 0.019
R79695 out.n4880 out.n4879 0.019
R79696 out.n4874 out.n4873 0.019
R79697 out.n4866 out.n4865 0.019
R79698 out.n4869 out.n4868 0.019
R79699 out.n4863 out.n4862 0.019
R79700 out.n4855 out.n4854 0.019
R79701 out.n4858 out.n4857 0.019
R79702 out.n4849 out.n4848 0.019
R79703 out.n4852 out.n4851 0.019
R79704 out.n4843 out.n4842 0.019
R79705 out.n4846 out.n4845 0.019
R79706 out.n4840 out.n4839 0.019
R79707 out.n14496 out.n14261 0.019
R79708 out.n1084 out.n957 0.019
R79709 out.n2043 out.n1897 0.019
R79710 out.n15389 out.n15388 0.019
R79711 out.n6576 out.n6575 0.019
R79712 out.n6686 out.n6685 0.019
R79713 out.n6011 out.n6010 0.019
R79714 out.n7735 out.n7734 0.019
R79715 out.n10017 out.n10016 0.019
R79716 out.n77 out.n76 0.019
R79717 out.n137 out.n136 0.019
R79718 out.n333 out.n332 0.019
R79719 out.n399 out.n398 0.019
R79720 out.n461 out.n460 0.019
R79721 out.n589 out.n588 0.019
R79722 out.n781 out.n780 0.019
R79723 out.n4931 out.n4930 0.019
R79724 out.n4299 out.n4298 0.019
R79725 out.n4367 out.n4366 0.019
R79726 out.n4432 out.n4431 0.019
R79727 out.n4494 out.n4493 0.019
R79728 out.n4559 out.n4558 0.019
R79729 out.n4823 out.n4822 0.019
R79730 out.n6583 out.n6582 0.019
R79731 out.n7742 out.n7741 0.019
R79732 out.n6760 out.n6759 0.019
R79733 out.n6684 out.n6683 0.019
R79734 out.n6124 out.n6123 0.019
R79735 out.n6009 out.n6008 0.019
R79736 out.n13149 out.n13148 0.019
R79737 out.n11864 out.n11863 0.019
R79738 out.n10597 out.n10596 0.019
R79739 out.n7633 out.n7632 0.019
R79740 out out.n17311 0.019
R79741 out.n9412 out.n9411 0.019
R79742 out.n9044 out.n9043 0.019
R79743 out.n1299 out.n1171 0.019
R79744 out.n2564 out.n2562 0.019
R79745 out.n6349 out.n6347 0.019
R79746 out.n5990 out.n5988 0.019
R79747 out.n13134 out.n13132 0.019
R79748 out.n13034 out.n13033 0.019
R79749 out.n12909 out.n12908 0.019
R79750 out.n11849 out.n11847 0.019
R79751 out.n11749 out.n11748 0.019
R79752 out.n11624 out.n11623 0.019
R79753 out.n10582 out.n10580 0.019
R79754 out.n10482 out.n10481 0.019
R79755 out.n10357 out.n10356 0.019
R79756 out.n6126 out.n6125 0.019
R79757 out.n14510 out.n14509 0.019
R79758 out.n13041 out.n13040 0.019
R79759 out.n12916 out.n12915 0.019
R79760 out.n11756 out.n11755 0.019
R79761 out.n11631 out.n11630 0.019
R79762 out.n10489 out.n10488 0.019
R79763 out.n10364 out.n10363 0.019
R79764 out.n6688 out.n6687 0.019
R79765 out.n6013 out.n6012 0.019
R79766 out.n6133 out.n6132 0.019
R79767 out.n13142 out.n13141 0.019
R79768 out.n13140 out.n13138 0.019
R79769 out.n13027 out.n13026 0.019
R79770 out.n12902 out.n12901 0.019
R79771 out.n11857 out.n11856 0.019
R79772 out.n11855 out.n11853 0.019
R79773 out.n11742 out.n11741 0.019
R79774 out.n11617 out.n11616 0.019
R79775 out.n10590 out.n10589 0.019
R79776 out.n10588 out.n10586 0.019
R79777 out.n10475 out.n10474 0.019
R79778 out.n10350 out.n10349 0.019
R79779 out.n7733 out.n7732 0.019
R79780 out.n2532 out.n2531 0.019
R79781 out.n13443 out.n13442 0.019
R79782 out.n13898 out.n13897 0.019
R79783 out.n6656 out.n6654 0.019
R79784 out.n10007 out.n10004 0.019
R79785 out.n10036 out.n10032 0.019
R79786 out.n16274 out.n16271 0.019
R79787 out.n10030 out.n10027 0.019
R79788 out.n16279 out.n16276 0.019
R79789 out.n10025 out.n10022 0.019
R79790 out.n10020 out.n10017 0.019
R79791 out.n16284 out.n16283 0.019
R79792 out.n4746 out.n4745 0.019
R79793 out.n4680 out.n4679 0.019
R79794 out.n4619 out.n4618 0.019
R79795 out.n4617 out.n4616 0.019
R79796 out.n4551 out.n4550 0.019
R79797 out.n4549 out.n4548 0.019
R79798 out.n4487 out.n4486 0.019
R79799 out.n4423 out.n4422 0.019
R79800 out.n4421 out.n4420 0.019
R79801 out.n4359 out.n4358 0.019
R79802 out.n4357 out.n4356 0.019
R79803 out.n4292 out.n4291 0.019
R79804 out.n4228 out.n4227 0.019
R79805 out.n4166 out.n4165 0.019
R79806 out.n4164 out.n4163 0.019
R79807 out.n4103 out.n4102 0.019
R79808 out.n4036 out.n4035 0.019
R79809 out.n836 out.n835 0.019
R79810 out.n715 out.n714 0.019
R79811 out.n581 out.n580 0.019
R79812 out.n579 out.n578 0.019
R79813 out.n390 out.n389 0.019
R79814 out.n324 out.n323 0.019
R79815 out.n128 out.n127 0.019
R79816 out.n68 out.n67 0.019
R79817 out.n66 out.n65 0.019
R79818 out.n30 out.n29 0.019
R79819 out.n4779 out.n4778 0.019
R79820 out.n4781 out.n4780 0.019
R79821 out.n4716 out.n4715 0.019
R79822 out.n4718 out.n4717 0.019
R79823 out.n4651 out.n4650 0.019
R79824 out.n4653 out.n4652 0.019
R79825 out.n4586 out.n4585 0.019
R79826 out.n4588 out.n4587 0.019
R79827 out.n4521 out.n4520 0.019
R79828 out.n4523 out.n4522 0.019
R79829 out.n4459 out.n4458 0.019
R79830 out.n4461 out.n4460 0.019
R79831 out.n4393 out.n4392 0.019
R79832 out.n4395 out.n4394 0.019
R79833 out.n4329 out.n4328 0.019
R79834 out.n4331 out.n4330 0.019
R79835 out.n4264 out.n4263 0.019
R79836 out.n4266 out.n4265 0.019
R79837 out.n4198 out.n4197 0.019
R79838 out.n4200 out.n4199 0.019
R79839 out.n4132 out.n4131 0.019
R79840 out.n4134 out.n4133 0.019
R79841 out.n4070 out.n4069 0.019
R79842 out.n4072 out.n4071 0.019
R79843 out.n4005 out.n4004 0.019
R79844 out.n4007 out.n4006 0.019
R79845 out.n4919 out.n4918 0.019
R79846 out.n875 out.n874 0.019
R79847 out.n807 out.n806 0.019
R79848 out.n809 out.n808 0.019
R79849 out.n744 out.n743 0.019
R79850 out.n746 out.n745 0.019
R79851 out.n682 out.n681 0.019
R79852 out.n684 out.n683 0.019
R79853 out.n617 out.n616 0.019
R79854 out.n619 out.n618 0.019
R79855 out.n552 out.n551 0.019
R79856 out.n554 out.n553 0.019
R79857 out.n490 out.n489 0.019
R79858 out.n492 out.n491 0.019
R79859 out.n424 out.n423 0.019
R79860 out.n426 out.n425 0.019
R79861 out.n360 out.n359 0.019
R79862 out.n362 out.n361 0.019
R79863 out.n291 out.n290 0.019
R79864 out.n293 out.n292 0.019
R79865 out.n230 out.n229 0.019
R79866 out.n232 out.n231 0.019
R79867 out.n164 out.n163 0.019
R79868 out.n166 out.n165 0.019
R79869 out.n100 out.n99 0.019
R79870 out.n102 out.n101 0.019
R79871 out.n25 out.n24 0.019
R79872 out.n9 out.n8 0.019
R79873 out.n58 out.n57 0.019
R79874 out.n91 out.n90 0.019
R79875 out.n121 out.n120 0.019
R79876 out.n152 out.n151 0.019
R79877 out.n187 out.n186 0.019
R79878 out.n217 out.n216 0.019
R79879 out.n253 out.n252 0.019
R79880 out.n277 out.n276 0.019
R79881 out.n315 out.n314 0.019
R79882 out.n347 out.n346 0.019
R79883 out.n383 out.n382 0.019
R79884 out.n412 out.n411 0.019
R79885 out.n446 out.n445 0.019
R79886 out.n476 out.n475 0.019
R79887 out.n513 out.n512 0.019
R79888 out.n537 out.n536 0.019
R79889 out.n574 out.n573 0.019
R79890 out.n605 out.n604 0.019
R79891 out.n640 out.n639 0.019
R79892 out.n668 out.n667 0.019
R79893 out.n707 out.n706 0.019
R79894 out.n732 out.n731 0.019
R79895 out.n770 out.n769 0.019
R79896 out.n795 out.n794 0.019
R79897 out.n830 out.n829 0.019
R79898 out.n862 out.n861 0.019
R79899 out.n867 out.n866 0.019
R79900 out.n4910 out.n4909 0.019
R79901 out.n4028 out.n4027 0.019
R79902 out.n4058 out.n4057 0.019
R79903 out.n4094 out.n4093 0.019
R79904 out.n4123 out.n4122 0.019
R79905 out.n4157 out.n4156 0.019
R79906 out.n4187 out.n4186 0.019
R79907 out.n4221 out.n4220 0.019
R79908 out.n4251 out.n4250 0.019
R79909 out.n4284 out.n4283 0.019
R79910 out.n4317 out.n4316 0.019
R79911 out.n4351 out.n4350 0.019
R79912 out.n4382 out.n4381 0.019
R79913 out.n4416 out.n4415 0.019
R79914 out.n4445 out.n4444 0.019
R79915 out.n4480 out.n4479 0.019
R79916 out.n4510 out.n4509 0.019
R79917 out.n4543 out.n4542 0.019
R79918 out.n4574 out.n4573 0.019
R79919 out.n4611 out.n4610 0.019
R79920 out.n4640 out.n4639 0.019
R79921 out.n4675 out.n4674 0.019
R79922 out.n4702 out.n4701 0.019
R79923 out.n4739 out.n4738 0.019
R79924 out.n4767 out.n4766 0.019
R79925 out.n4804 out.n4803 0.019
R79926 out.n174 out.n173 0.019
R79927 out.n241 out.n240 0.019
R79928 out.n499 out.n498 0.019
R79929 out.n627 out.n626 0.019
R79930 out.n693 out.n692 0.019
R79931 out.n815 out.n814 0.019
R79932 out.n4015 out.n4014 0.019
R79933 out.n4081 out.n4080 0.019
R79934 out.n4142 out.n4141 0.019
R79935 out.n4208 out.n4207 0.019
R79936 out.n4597 out.n4596 0.019
R79937 out.n4662 out.n4661 0.019
R79938 out.n4726 out.n4725 0.019
R79939 out.n335 out.n334 0.019
R79940 out.n306 out.n304 0.019
R79941 out.n591 out.n590 0.019
R79942 out.n564 out.n562 0.019
R79943 out.n697 out.n696 0.019
R79944 out.n757 out.n755 0.019
R79945 out.n847 out.n846 0.019
R79946 out.n820 out.n818 0.019
R79947 out.n893 out.n892 0.019
R79948 out.n913 out.n912 0.019
R79949 out.n4146 out.n4145 0.019
R79950 out.n4301 out.n4300 0.019
R79951 out.n4341 out.n4339 0.019
R79952 out.n4561 out.n4560 0.019
R79953 out.n4534 out.n4532 0.019
R79954 out.n4601 out.n4600 0.019
R79955 out.n55 out.n54 0.019
R79956 out.n84 out.n83 0.019
R79957 out.n143 out.n142 0.019
R79958 out.n183 out.n182 0.019
R79959 out.n208 out.n207 0.019
R79960 out.n249 out.n248 0.019
R79961 out.n270 out.n269 0.019
R79962 out.n340 out.n339 0.019
R79963 out.n378 out.n377 0.019
R79964 out.n405 out.n404 0.019
R79965 out.n441 out.n440 0.019
R79966 out.n467 out.n466 0.019
R79967 out.n509 out.n508 0.019
R79968 out.n570 out.n569 0.019
R79969 out.n597 out.n596 0.019
R79970 out.n635 out.n634 0.019
R79971 out.n659 out.n658 0.019
R79972 out.n703 out.n702 0.019
R79973 out.n765 out.n764 0.019
R79974 out.n825 out.n824 0.019
R79975 out.n853 out.n852 0.019
R79976 out.n4938 out.n4937 0.019
R79977 out.n4023 out.n4022 0.019
R79978 out.n4050 out.n4049 0.019
R79979 out.n4089 out.n4088 0.019
R79980 out.n4116 out.n4115 0.019
R79981 out.n4152 out.n4151 0.019
R79982 out.n4216 out.n4215 0.019
R79983 out.n4243 out.n4242 0.019
R79984 out.n4279 out.n4278 0.019
R79985 out.n4308 out.n4307 0.019
R79986 out.n4374 out.n4373 0.019
R79987 out.n4411 out.n4410 0.019
R79988 out.n4475 out.n4474 0.019
R79989 out.n4501 out.n4500 0.019
R79990 out.n4566 out.n4565 0.019
R79991 out.n4606 out.n4605 0.019
R79992 out.n4633 out.n4632 0.019
R79993 out.n4670 out.n4669 0.019
R79994 out.n4695 out.n4694 0.019
R79995 out.n4734 out.n4733 0.019
R79996 out.n4759 out.n4758 0.019
R79997 out.n4829 out.n4828 0.019
R79998 out.n11 out.n10 0.019
R79999 out.n280 out.n279 0.019
R80000 out.n349 out.n348 0.019
R80001 out.n351 out.n350 0.019
R80002 out.n540 out.n539 0.019
R80003 out.n670 out.n669 0.019
R80004 out.n3996 out.n3995 0.019
R80005 out.n4060 out.n4059 0.019
R80006 out.n4190 out.n4189 0.019
R80007 out.n4253 out.n4252 0.019
R80008 out.n4319 out.n4318 0.019
R80009 out.n4447 out.n4446 0.019
R80010 out.n4576 out.n4575 0.019
R80011 out.n7635 out.n7634 0.019
R80012 out.n2017 out.n2016 0.019
R80013 out.n12169 out.n12168 0.019
R80014 out.n12044 out.n12043 0.019
R80015 out.n13318 out.n13317 0.019
R80016 out.n13773 out.n13772 0.019
R80017 out.n1514 out.n1512 0.019
R80018 out.n2361 out.n2359 0.019
R80019 out.n17184 out.n17183 0.019
R80020 out.n17082 out.n17081 0.019
R80021 out.n17047 out.n17046 0.019
R80022 out.n17016 out.n17015 0.019
R80023 out.n16983 out.n16982 0.019
R80024 out.n16950 out.n16949 0.019
R80025 out.n16915 out.n16914 0.019
R80026 out.n16884 out.n16883 0.019
R80027 out.n16851 out.n16850 0.019
R80028 out.n16818 out.n16817 0.019
R80029 out.n16785 out.n16784 0.019
R80030 out.n16752 out.n16751 0.019
R80031 out.n16717 out.n16716 0.019
R80032 out.n16686 out.n16685 0.019
R80033 out.n16651 out.n16650 0.019
R80034 out.n16620 out.n16619 0.019
R80035 out.n16587 out.n16586 0.019
R80036 out.n16554 out.n16553 0.019
R80037 out.n16519 out.n16518 0.019
R80038 out.n16490 out.n16489 0.019
R80039 out.n16453 out.n16452 0.019
R80040 out.n16424 out.n16423 0.019
R80041 out.n16387 out.n16386 0.019
R80042 out.n16356 out.n16355 0.019
R80043 out.n16321 out.n16320 0.019
R80044 out.n16290 out.n16289 0.019
R80045 out.n10003 out.n10002 0.019
R80046 out.n9966 out.n9965 0.019
R80047 out.n9058 out.n9057 0.019
R80048 out.n9928 out.n9927 0.019
R80049 out.n9894 out.n9893 0.019
R80050 out.n9862 out.n9861 0.019
R80051 out.n9091 out.n9090 0.019
R80052 out.n9823 out.n9822 0.019
R80053 out.n9125 out.n9124 0.019
R80054 out.n9787 out.n9786 0.019
R80055 out.n9159 out.n9158 0.019
R80056 out.n9751 out.n9750 0.019
R80057 out.n9193 out.n9192 0.019
R80058 out.n9715 out.n9714 0.019
R80059 out.n9227 out.n9226 0.019
R80060 out.n9679 out.n9678 0.019
R80061 out.n9261 out.n9260 0.019
R80062 out.n9623 out.n9622 0.019
R80063 out.n9294 out.n9293 0.019
R80064 out.n9584 out.n9583 0.019
R80065 out.n9328 out.n9327 0.019
R80066 out.n9548 out.n9547 0.019
R80067 out.n9362 out.n9361 0.019
R80068 out.n9512 out.n9511 0.019
R80069 out.n9395 out.n9394 0.019
R80070 out.n9471 out.n9470 0.019
R80071 out.n9409 out.n9408 0.019
R80072 out.n9524 out.n9523 0.019
R80073 out.n9377 out.n9376 0.019
R80074 out.n9560 out.n9559 0.019
R80075 out.n9343 out.n9342 0.019
R80076 out.n9596 out.n9595 0.019
R80077 out.n9309 out.n9308 0.019
R80078 out.n9635 out.n9634 0.019
R80079 out.n9276 out.n9275 0.019
R80080 out.n9691 out.n9690 0.019
R80081 out.n9242 out.n9241 0.019
R80082 out.n9727 out.n9726 0.019
R80083 out.n9208 out.n9207 0.019
R80084 out.n9763 out.n9762 0.019
R80085 out.n9174 out.n9173 0.019
R80086 out.n9799 out.n9798 0.019
R80087 out.n9140 out.n9139 0.019
R80088 out.n9835 out.n9834 0.019
R80089 out.n9106 out.n9105 0.019
R80090 out.n9874 out.n9873 0.019
R80091 out.n9909 out.n9908 0.019
R80092 out.n9940 out.n9939 0.019
R80093 out.n9073 out.n9072 0.019
R80094 out.n9978 out.n9977 0.019
R80095 out.n9039 out.n9038 0.019
R80096 out.n16305 out.n16304 0.019
R80097 out.n16333 out.n16332 0.019
R80098 out.n16371 out.n16370 0.019
R80099 out.n16399 out.n16398 0.019
R80100 out.n16439 out.n16438 0.019
R80101 out.n16465 out.n16464 0.019
R80102 out.n16505 out.n16504 0.019
R80103 out.n16531 out.n16530 0.019
R80104 out.n16569 out.n16568 0.019
R80105 out.n16599 out.n16598 0.019
R80106 out.n16635 out.n16634 0.019
R80107 out.n16663 out.n16662 0.019
R80108 out.n16701 out.n16700 0.019
R80109 out.n16729 out.n16728 0.019
R80110 out.n16767 out.n16766 0.019
R80111 out.n16797 out.n16796 0.019
R80112 out.n16833 out.n16832 0.019
R80113 out.n16863 out.n16862 0.019
R80114 out.n16899 out.n16898 0.019
R80115 out.n16927 out.n16926 0.019
R80116 out.n16965 out.n16964 0.019
R80117 out.n16995 out.n16994 0.019
R80118 out.n17031 out.n17030 0.019
R80119 out.n17059 out.n17058 0.019
R80120 out.n17097 out.n17096 0.019
R80121 out.n17123 out.n17122 0.019
R80122 out.n17175 out.n17174 0.019
R80123 out.n9416 out.n9415 0.019
R80124 out.n9531 out.n9530 0.019
R80125 out.n9384 out.n9383 0.019
R80126 out.n9567 out.n9566 0.019
R80127 out.n9350 out.n9349 0.019
R80128 out.n9603 out.n9602 0.019
R80129 out.n9316 out.n9315 0.019
R80130 out.n9642 out.n9641 0.019
R80131 out.n9283 out.n9282 0.019
R80132 out.n9698 out.n9697 0.019
R80133 out.n9249 out.n9248 0.019
R80134 out.n9734 out.n9733 0.019
R80135 out.n9215 out.n9214 0.019
R80136 out.n9770 out.n9769 0.019
R80137 out.n9181 out.n9180 0.019
R80138 out.n9806 out.n9805 0.019
R80139 out.n9147 out.n9146 0.019
R80140 out.n9842 out.n9841 0.019
R80141 out.n9113 out.n9112 0.019
R80142 out.n9881 out.n9880 0.019
R80143 out.n9916 out.n9915 0.019
R80144 out.n9949 out.n9948 0.019
R80145 out.n9078 out.n9077 0.019
R80146 out.n9985 out.n9984 0.019
R80147 out.n9047 out.n9046 0.019
R80148 out.n16312 out.n16311 0.019
R80149 out.n16340 out.n16339 0.019
R80150 out.n16378 out.n16377 0.019
R80151 out.n16408 out.n16407 0.019
R80152 out.n16444 out.n16443 0.019
R80153 out.n16474 out.n16473 0.019
R80154 out.n16510 out.n16509 0.019
R80155 out.n16538 out.n16537 0.019
R80156 out.n16578 out.n16577 0.019
R80157 out.n16604 out.n16603 0.019
R80158 out.n16642 out.n16641 0.019
R80159 out.n16670 out.n16669 0.019
R80160 out.n16708 out.n16707 0.019
R80161 out.n16736 out.n16735 0.019
R80162 out.n16776 out.n16775 0.019
R80163 out.n16802 out.n16801 0.019
R80164 out.n16842 out.n16841 0.019
R80165 out.n16868 out.n16867 0.019
R80166 out.n16906 out.n16905 0.019
R80167 out.n16934 out.n16933 0.019
R80168 out.n16974 out.n16973 0.019
R80169 out.n17000 out.n16999 0.019
R80170 out.n17038 out.n17037 0.019
R80171 out.n17066 out.n17065 0.019
R80172 out.n17104 out.n17103 0.019
R80173 out.n17132 out.n17131 0.019
R80174 out.n17170 out.n17169 0.019
R80175 out.n9406 out.n9405 0.019
R80176 out.n9521 out.n9520 0.019
R80177 out.n9374 out.n9373 0.019
R80178 out.n9557 out.n9556 0.019
R80179 out.n9340 out.n9339 0.019
R80180 out.n9593 out.n9592 0.019
R80181 out.n9306 out.n9305 0.019
R80182 out.n9632 out.n9631 0.019
R80183 out.n9273 out.n9272 0.019
R80184 out.n9688 out.n9687 0.019
R80185 out.n9239 out.n9238 0.019
R80186 out.n9724 out.n9723 0.019
R80187 out.n9205 out.n9204 0.019
R80188 out.n9760 out.n9759 0.019
R80189 out.n9171 out.n9170 0.019
R80190 out.n9796 out.n9795 0.019
R80191 out.n9137 out.n9136 0.019
R80192 out.n9832 out.n9831 0.019
R80193 out.n9103 out.n9102 0.019
R80194 out.n9871 out.n9870 0.019
R80195 out.n9906 out.n9905 0.019
R80196 out.n9937 out.n9936 0.019
R80197 out.n9070 out.n9069 0.019
R80198 out.n9975 out.n9974 0.019
R80199 out.n9035 out.n9034 0.019
R80200 out.n16302 out.n16301 0.019
R80201 out.n16330 out.n16329 0.019
R80202 out.n16368 out.n16367 0.019
R80203 out.n16396 out.n16395 0.019
R80204 out.n16436 out.n16435 0.019
R80205 out.n16462 out.n16461 0.019
R80206 out.n16502 out.n16501 0.019
R80207 out.n16528 out.n16527 0.019
R80208 out.n16566 out.n16565 0.019
R80209 out.n16596 out.n16595 0.019
R80210 out.n16632 out.n16631 0.019
R80211 out.n16660 out.n16659 0.019
R80212 out.n16698 out.n16697 0.019
R80213 out.n16726 out.n16725 0.019
R80214 out.n16764 out.n16763 0.019
R80215 out.n16794 out.n16793 0.019
R80216 out.n16830 out.n16829 0.019
R80217 out.n16860 out.n16859 0.019
R80218 out.n16896 out.n16895 0.019
R80219 out.n16924 out.n16923 0.019
R80220 out.n16962 out.n16961 0.019
R80221 out.n16992 out.n16991 0.019
R80222 out.n17028 out.n17027 0.019
R80223 out.n17056 out.n17055 0.019
R80224 out.n17094 out.n17093 0.019
R80225 out.n17120 out.n17119 0.019
R80226 out.n17168 out.n17167 0.019
R80227 out.n9419 out.n9418 0.019
R80228 out.n9535 out.n9533 0.019
R80229 out.n9387 out.n9386 0.019
R80230 out.n9571 out.n9569 0.019
R80231 out.n9353 out.n9352 0.019
R80232 out.n9607 out.n9605 0.019
R80233 out.n9319 out.n9318 0.019
R80234 out.n9646 out.n9644 0.019
R80235 out.n9286 out.n9285 0.019
R80236 out.n9702 out.n9700 0.019
R80237 out.n9252 out.n9251 0.019
R80238 out.n9738 out.n9736 0.019
R80239 out.n9218 out.n9217 0.019
R80240 out.n9774 out.n9772 0.019
R80241 out.n9184 out.n9183 0.019
R80242 out.n9810 out.n9808 0.019
R80243 out.n9150 out.n9149 0.019
R80244 out.n9846 out.n9844 0.019
R80245 out.n9116 out.n9115 0.019
R80246 out.n9885 out.n9883 0.019
R80247 out.n9919 out.n9918 0.019
R80248 out.n9953 out.n9951 0.019
R80249 out.n9081 out.n9080 0.019
R80250 out.n9989 out.n9987 0.019
R80251 out.n9049 out.n9048 0.019
R80252 out.n16315 out.n16314 0.019
R80253 out.n16344 out.n16342 0.019
R80254 out.n16381 out.n16380 0.019
R80255 out.n16412 out.n16410 0.019
R80256 out.n16447 out.n16446 0.019
R80257 out.n16478 out.n16476 0.019
R80258 out.n16513 out.n16512 0.019
R80259 out.n16542 out.n16540 0.019
R80260 out.n16581 out.n16580 0.019
R80261 out.n16608 out.n16606 0.019
R80262 out.n16645 out.n16644 0.019
R80263 out.n16674 out.n16672 0.019
R80264 out.n16711 out.n16710 0.019
R80265 out.n16740 out.n16738 0.019
R80266 out.n16779 out.n16778 0.019
R80267 out.n16806 out.n16804 0.019
R80268 out.n16845 out.n16844 0.019
R80269 out.n16872 out.n16870 0.019
R80270 out.n16909 out.n16908 0.019
R80271 out.n16938 out.n16936 0.019
R80272 out.n16977 out.n16976 0.019
R80273 out.n17004 out.n17002 0.019
R80274 out.n17041 out.n17040 0.019
R80275 out.n17070 out.n17068 0.019
R80276 out.n17107 out.n17106 0.019
R80277 out.n17136 out.n17134 0.019
R80278 out.n17166 out.n17165 0.019
R80279 out.n17155 out.n17154 0.019
R80280 out.n17117 out.n17116 0.019
R80281 out.n17085 out.n17084 0.019
R80282 out.n17053 out.n17052 0.019
R80283 out.n17019 out.n17018 0.019
R80284 out.n16989 out.n16988 0.019
R80285 out.n16953 out.n16952 0.019
R80286 out.n16921 out.n16920 0.019
R80287 out.n16887 out.n16886 0.019
R80288 out.n16857 out.n16856 0.019
R80289 out.n16821 out.n16820 0.019
R80290 out.n16791 out.n16790 0.019
R80291 out.n16755 out.n16754 0.019
R80292 out.n16723 out.n16722 0.019
R80293 out.n16689 out.n16688 0.019
R80294 out.n16657 out.n16656 0.019
R80295 out.n16623 out.n16622 0.019
R80296 out.n16593 out.n16592 0.019
R80297 out.n16557 out.n16556 0.019
R80298 out.n16525 out.n16524 0.019
R80299 out.n16493 out.n16492 0.019
R80300 out.n16459 out.n16458 0.019
R80301 out.n16427 out.n16426 0.019
R80302 out.n16393 out.n16392 0.019
R80303 out.n16359 out.n16358 0.019
R80304 out.n16327 out.n16326 0.019
R80305 out.n16293 out.n16292 0.019
R80306 out.n9031 out.n9030 0.019
R80307 out.n9025 out.n9024 0.019
R80308 out.n9972 out.n9971 0.019
R80309 out.n9061 out.n9060 0.019
R80310 out.n9934 out.n9933 0.019
R80311 out.n9897 out.n9896 0.019
R80312 out.n9868 out.n9867 0.019
R80313 out.n9094 out.n9093 0.019
R80314 out.n9829 out.n9828 0.019
R80315 out.n9128 out.n9127 0.019
R80316 out.n9793 out.n9792 0.019
R80317 out.n9162 out.n9161 0.019
R80318 out.n9757 out.n9756 0.019
R80319 out.n9196 out.n9195 0.019
R80320 out.n9721 out.n9720 0.019
R80321 out.n9230 out.n9229 0.019
R80322 out.n9685 out.n9684 0.019
R80323 out.n9264 out.n9263 0.019
R80324 out.n9629 out.n9628 0.019
R80325 out.n9297 out.n9296 0.019
R80326 out.n9590 out.n9589 0.019
R80327 out.n9331 out.n9330 0.019
R80328 out.n9554 out.n9553 0.019
R80329 out.n9365 out.n9364 0.019
R80330 out.n9518 out.n9517 0.019
R80331 out.n17164 out.n17163 0.019
R80332 out.n17113 out.n17112 0.019
R80333 out.n17092 out.n17091 0.019
R80334 out.n17049 out.n17048 0.019
R80335 out.n17026 out.n17025 0.019
R80336 out.n16985 out.n16984 0.019
R80337 out.n16960 out.n16959 0.019
R80338 out.n16917 out.n16916 0.019
R80339 out.n16894 out.n16893 0.019
R80340 out.n16853 out.n16852 0.019
R80341 out.n16828 out.n16827 0.019
R80342 out.n16787 out.n16786 0.019
R80343 out.n16762 out.n16761 0.019
R80344 out.n16719 out.n16718 0.019
R80345 out.n16696 out.n16695 0.019
R80346 out.n16653 out.n16652 0.019
R80347 out.n16630 out.n16629 0.019
R80348 out.n16589 out.n16588 0.019
R80349 out.n16564 out.n16563 0.019
R80350 out.n16521 out.n16520 0.019
R80351 out.n16500 out.n16499 0.019
R80352 out.n16455 out.n16454 0.019
R80353 out.n16434 out.n16433 0.019
R80354 out.n16389 out.n16388 0.019
R80355 out.n16366 out.n16365 0.019
R80356 out.n16323 out.n16322 0.019
R80357 out.n16300 out.n16299 0.019
R80358 out.n9033 out.n9032 0.019
R80359 out.n9968 out.n9967 0.019
R80360 out.n9068 out.n9067 0.019
R80361 out.n9930 out.n9929 0.019
R80362 out.n9904 out.n9903 0.019
R80363 out.n9864 out.n9863 0.019
R80364 out.n9101 out.n9100 0.019
R80365 out.n9825 out.n9824 0.019
R80366 out.n9135 out.n9134 0.019
R80367 out.n9789 out.n9788 0.019
R80368 out.n9169 out.n9168 0.019
R80369 out.n9753 out.n9752 0.019
R80370 out.n9203 out.n9202 0.019
R80371 out.n9717 out.n9716 0.019
R80372 out.n9237 out.n9236 0.019
R80373 out.n9681 out.n9680 0.019
R80374 out.n9271 out.n9270 0.019
R80375 out.n9625 out.n9624 0.019
R80376 out.n9304 out.n9303 0.019
R80377 out.n9586 out.n9585 0.019
R80378 out.n9338 out.n9337 0.019
R80379 out.n9550 out.n9549 0.019
R80380 out.n9372 out.n9371 0.019
R80381 out.n9401 out.n9400 0.019
R80382 out.n9404 out.n9403 0.019
R80383 out.n9370 out.n9369 0.019
R80384 out.n9368 out.n9367 0.019
R80385 out.n9336 out.n9335 0.019
R80386 out.n9334 out.n9333 0.019
R80387 out.n9302 out.n9301 0.019
R80388 out.n9300 out.n9299 0.019
R80389 out.n9269 out.n9268 0.019
R80390 out.n9267 out.n9266 0.019
R80391 out.n9235 out.n9234 0.019
R80392 out.n9233 out.n9232 0.019
R80393 out.n9201 out.n9200 0.019
R80394 out.n9199 out.n9198 0.019
R80395 out.n9167 out.n9166 0.019
R80396 out.n9165 out.n9164 0.019
R80397 out.n9133 out.n9132 0.019
R80398 out.n9131 out.n9130 0.019
R80399 out.n9099 out.n9098 0.019
R80400 out.n9097 out.n9096 0.019
R80401 out.n9902 out.n9901 0.019
R80402 out.n9900 out.n9899 0.019
R80403 out.n9066 out.n9065 0.019
R80404 out.n9064 out.n9063 0.019
R80405 out.n9028 out.n9027 0.019
R80406 out.n16298 out.n16297 0.019
R80407 out.n16296 out.n16295 0.019
R80408 out.n16364 out.n16363 0.019
R80409 out.n16362 out.n16361 0.019
R80410 out.n16432 out.n16431 0.019
R80411 out.n16430 out.n16429 0.019
R80412 out.n16498 out.n16497 0.019
R80413 out.n16496 out.n16495 0.019
R80414 out.n16562 out.n16561 0.019
R80415 out.n16560 out.n16559 0.019
R80416 out.n16628 out.n16627 0.019
R80417 out.n16626 out.n16625 0.019
R80418 out.n16694 out.n16693 0.019
R80419 out.n16692 out.n16691 0.019
R80420 out.n16760 out.n16759 0.019
R80421 out.n16758 out.n16757 0.019
R80422 out.n16826 out.n16825 0.019
R80423 out.n16824 out.n16823 0.019
R80424 out.n16892 out.n16891 0.019
R80425 out.n16890 out.n16889 0.019
R80426 out.n16958 out.n16957 0.019
R80427 out.n16956 out.n16955 0.019
R80428 out.n17024 out.n17023 0.019
R80429 out.n17022 out.n17021 0.019
R80430 out.n17090 out.n17089 0.019
R80431 out.n17088 out.n17087 0.019
R80432 out.n17159 out.n17158 0.019
R80433 out.n9487 out.n9486 0.019
R80434 out.n9516 out.n9515 0.019
R80435 out.n9397 out.n9396 0.019
R80436 out.n9538 out.n9537 0.019
R80437 out.n9421 out.n9420 0.019
R80438 out.n9389 out.n9388 0.019
R80439 out.n9574 out.n9573 0.019
R80440 out.n9355 out.n9354 0.019
R80441 out.n9610 out.n9609 0.019
R80442 out.n9321 out.n9320 0.019
R80443 out.n9649 out.n9648 0.019
R80444 out.n9288 out.n9287 0.019
R80445 out.n9705 out.n9704 0.019
R80446 out.n9254 out.n9253 0.019
R80447 out.n9741 out.n9740 0.019
R80448 out.n9220 out.n9219 0.019
R80449 out.n9777 out.n9776 0.019
R80450 out.n9186 out.n9185 0.019
R80451 out.n9813 out.n9812 0.019
R80452 out.n9152 out.n9151 0.019
R80453 out.n9849 out.n9848 0.019
R80454 out.n9118 out.n9117 0.019
R80455 out.n9888 out.n9887 0.019
R80456 out.n9921 out.n9920 0.019
R80457 out.n9956 out.n9955 0.019
R80458 out.n9083 out.n9082 0.019
R80459 out.n9992 out.n9991 0.019
R80460 out.n9051 out.n9050 0.019
R80461 out.n16317 out.n16316 0.019
R80462 out.n16347 out.n16346 0.019
R80463 out.n16383 out.n16382 0.019
R80464 out.n16415 out.n16414 0.019
R80465 out.n16449 out.n16448 0.019
R80466 out.n16481 out.n16480 0.019
R80467 out.n16515 out.n16514 0.019
R80468 out.n16545 out.n16544 0.019
R80469 out.n16583 out.n16582 0.019
R80470 out.n16611 out.n16610 0.019
R80471 out.n16647 out.n16646 0.019
R80472 out.n16677 out.n16676 0.019
R80473 out.n16713 out.n16712 0.019
R80474 out.n16743 out.n16742 0.019
R80475 out.n16781 out.n16780 0.019
R80476 out.n16809 out.n16808 0.019
R80477 out.n16847 out.n16846 0.019
R80478 out.n16875 out.n16874 0.019
R80479 out.n16911 out.n16910 0.019
R80480 out.n16941 out.n16940 0.019
R80481 out.n16979 out.n16978 0.019
R80482 out.n17007 out.n17006 0.019
R80483 out.n17043 out.n17042 0.019
R80484 out.n17073 out.n17072 0.019
R80485 out.n17109 out.n17108 0.019
R80486 out.n17140 out.n17139 0.019
R80487 out.n17138 out.n17137 0.019
R80488 out.n4774 out.n4773 0.019
R80489 out.n4710 out.n4709 0.019
R80490 out.n4712 out.n4711 0.019
R80491 out.n4454 out.n4453 0.019
R80492 out.n4259 out.n4258 0.019
R80493 out.n4261 out.n4260 0.019
R80494 out.n4066 out.n4065 0.019
R80495 out.n4000 out.n3999 0.019
R80496 out.n4002 out.n4001 0.019
R80497 out.n4917 out.n4916 0.019
R80498 out.n871 out.n870 0.019
R80499 out.n803 out.n802 0.019
R80500 out.n738 out.n737 0.019
R80501 out.n676 out.n675 0.019
R80502 out.n678 out.n677 0.019
R80503 out.n612 out.n611 0.019
R80504 out.n547 out.n546 0.019
R80505 out.n483 out.n482 0.019
R80506 out.n485 out.n484 0.019
R80507 out.n419 out.n418 0.019
R80508 out.n355 out.n354 0.019
R80509 out.n286 out.n285 0.019
R80510 out.n288 out.n287 0.019
R80511 out.n224 out.n223 0.019
R80512 out.n226 out.n225 0.019
R80513 out.n159 out.n158 0.019
R80514 out.n161 out.n160 0.019
R80515 out.n80 out.n79 0.019
R80516 out.n51 out.n50 0.019
R80517 out.n43 out.n42 0.019
R80518 out.n140 out.n139 0.019
R80519 out.n114 out.n113 0.019
R80520 out.n205 out.n204 0.019
R80521 out.n180 out.n179 0.019
R80522 out.n246 out.n245 0.019
R80523 out.n337 out.n336 0.019
R80524 out.n402 out.n401 0.019
R80525 out.n375 out.n374 0.019
R80526 out.n464 out.n463 0.019
R80527 out.n438 out.n437 0.019
R80528 out.n505 out.n504 0.019
R80529 out.n593 out.n592 0.019
R80530 out.n632 out.n631 0.019
R80531 out.n699 out.n698 0.019
R80532 out.n760 out.n759 0.019
R80533 out.n4935 out.n4934 0.019
R80534 out.n4047 out.n4046 0.019
R80535 out.n4020 out.n4019 0.019
R80536 out.n4086 out.n4085 0.019
R80537 out.n4177 out.n4176 0.019
R80538 out.n4148 out.n4147 0.019
R80539 out.n4240 out.n4239 0.019
R80540 out.n4213 out.n4212 0.019
R80541 out.n4370 out.n4369 0.019
R80542 out.n4344 out.n4343 0.019
R80543 out.n4435 out.n4434 0.019
R80544 out.n4407 out.n4406 0.019
R80545 out.n4472 out.n4471 0.019
R80546 out.n4630 out.n4629 0.019
R80547 out.n4603 out.n4602 0.019
R80548 out.n4692 out.n4691 0.019
R80549 out.n4667 out.n4666 0.019
R80550 out.n4755 out.n4754 0.019
R80551 out.n4731 out.n4730 0.019
R80552 out.n4794 out.n4793 0.019
R80553 out.n40 out.n39 0.019
R80554 out.n73 out.n72 0.019
R80555 out.n107 out.n106 0.019
R80556 out.n134 out.n133 0.019
R80557 out.n171 out.n170 0.019
R80558 out.n199 out.n198 0.019
R80559 out.n238 out.n237 0.019
R80560 out.n262 out.n261 0.019
R80561 out.n299 out.n298 0.019
R80562 out.n329 out.n328 0.019
R80563 out.n368 out.n367 0.019
R80564 out.n395 out.n394 0.019
R80565 out.n431 out.n430 0.019
R80566 out.n457 out.n456 0.019
R80567 out.n496 out.n495 0.019
R80568 out.n521 out.n520 0.019
R80569 out.n558 out.n557 0.019
R80570 out.n586 out.n585 0.019
R80571 out.n624 out.n623 0.019
R80572 out.n651 out.n650 0.019
R80573 out.n690 out.n689 0.019
R80574 out.n719 out.n718 0.019
R80575 out.n750 out.n749 0.019
R80576 out.n779 out.n778 0.019
R80577 out.n813 out.n812 0.019
R80578 out.n842 out.n841 0.019
R80579 out.n889 out.n888 0.019
R80580 out.n4926 out.n4925 0.019
R80581 out.n4012 out.n4011 0.019
R80582 out.n4041 out.n4040 0.019
R80583 out.n4078 out.n4077 0.019
R80584 out.n4108 out.n4107 0.019
R80585 out.n4139 out.n4138 0.019
R80586 out.n4171 out.n4170 0.019
R80587 out.n4205 out.n4204 0.019
R80588 out.n4234 out.n4233 0.019
R80589 out.n4270 out.n4269 0.019
R80590 out.n4296 out.n4295 0.019
R80591 out.n4335 out.n4334 0.019
R80592 out.n4364 out.n4363 0.019
R80593 out.n4400 out.n4399 0.019
R80594 out.n4428 out.n4427 0.019
R80595 out.n4465 out.n4464 0.019
R80596 out.n4491 out.n4490 0.019
R80597 out.n4527 out.n4526 0.019
R80598 out.n4556 out.n4555 0.019
R80599 out.n4594 out.n4593 0.019
R80600 out.n4624 out.n4623 0.019
R80601 out.n4659 out.n4658 0.019
R80602 out.n4686 out.n4685 0.019
R80603 out.n4723 out.n4722 0.019
R80604 out.n4750 out.n4749 0.019
R80605 out.n4785 out.n4784 0.019
R80606 out.n4817 out.n4816 0.019
R80607 out.n82 out.n81 0.019
R80608 out.n268 out.n267 0.019
R80609 out.n507 out.n506 0.019
R80610 out.n701 out.n700 0.019
R80611 out.n762 out.n761 0.019
R80612 out.n850 out.n849 0.019
R80613 out.n4150 out.n4149 0.019
R80614 out.n4305 out.n4304 0.019
R80615 out.n4409 out.n4408 0.019
R80616 out.n4498 out.n4497 0.019
R80617 out.n4757 out.n4756 0.019
R80618 out.n36 out.n33 0.019
R80619 out.n104 out.n103 0.019
R80620 out.n71 out.n70 0.019
R80621 out.n32 out.n31 0.019
R80622 out.n168 out.n167 0.019
R80623 out.n131 out.n130 0.019
R80624 out.n260 out.n259 0.019
R80625 out.n236 out.n235 0.019
R80626 out.n196 out.n195 0.019
R80627 out.n326 out.n325 0.019
R80628 out.n296 out.n295 0.019
R80629 out.n392 out.n391 0.019
R80630 out.n365 out.n364 0.019
R80631 out.n454 out.n453 0.019
R80632 out.n428 out.n427 0.019
R80633 out.n519 out.n518 0.019
R80634 out.n494 out.n493 0.019
R80635 out.n583 out.n582 0.019
R80636 out.n556 out.n555 0.019
R80637 out.n648 out.n647 0.019
R80638 out.n621 out.n620 0.019
R80639 out.n717 out.n716 0.019
R80640 out.n687 out.n686 0.019
R80641 out.n777 out.n776 0.019
R80642 out.n748 out.n747 0.019
R80643 out.n839 out.n838 0.019
R80644 out.n811 out.n810 0.019
R80645 out.n4923 out.n4922 0.019
R80646 out.n4941 out.n4940 0.019
R80647 out.n4038 out.n4037 0.019
R80648 out.n4009 out.n4008 0.019
R80649 out.n4105 out.n4104 0.019
R80650 out.n4075 out.n4074 0.019
R80651 out.n4168 out.n4167 0.019
R80652 out.n4136 out.n4135 0.019
R80653 out.n4231 out.n4230 0.019
R80654 out.n4202 out.n4201 0.019
R80655 out.n4294 out.n4293 0.019
R80656 out.n4268 out.n4267 0.019
R80657 out.n4361 out.n4360 0.019
R80658 out.n4333 out.n4332 0.019
R80659 out.n4425 out.n4424 0.019
R80660 out.n4397 out.n4396 0.019
R80661 out.n4489 out.n4488 0.019
R80662 out.n4463 out.n4462 0.019
R80663 out.n4553 out.n4552 0.019
R80664 out.n4525 out.n4524 0.019
R80665 out.n4621 out.n4620 0.019
R80666 out.n4591 out.n4590 0.019
R80667 out.n4683 out.n4682 0.019
R80668 out.n4656 out.n4655 0.019
R80669 out.n4748 out.n4747 0.019
R80670 out.n4720 out.n4719 0.019
R80671 out.n4783 out.n4782 0.019
R80672 out.n18 out.n17 0.019
R80673 out.n118 out.n117 0.019
R80674 out.n87 out.n86 0.019
R80675 out.n147 out.n146 0.019
R80676 out.n145 out.n144 0.019
R80677 out.n212 out.n211 0.019
R80678 out.n210 out.n209 0.019
R80679 out.n312 out.n311 0.019
R80680 out.n273 out.n272 0.019
R80681 out.n380 out.n379 0.019
R80682 out.n343 out.n342 0.019
R80683 out.n443 out.n442 0.019
R80684 out.n408 out.n407 0.019
R80685 out.n471 out.n470 0.019
R80686 out.n469 out.n468 0.019
R80687 out.n532 out.n531 0.019
R80688 out.n530 out.n529 0.019
R80689 out.n637 out.n636 0.019
R80690 out.n600 out.n599 0.019
R80691 out.n663 out.n662 0.019
R80692 out.n661 out.n660 0.019
R80693 out.n767 out.n766 0.019
R80694 out.n728 out.n727 0.019
R80695 out.n827 out.n826 0.019
R80696 out.n790 out.n789 0.019
R80697 out.n857 out.n856 0.019
R80698 out.n855 out.n854 0.019
R80699 out.n4053 out.n4052 0.019
R80700 out.n4025 out.n4024 0.019
R80701 out.n4119 out.n4118 0.019
R80702 out.n4091 out.n4090 0.019
R80703 out.n4182 out.n4181 0.019
R80704 out.n4154 out.n4153 0.019
R80705 out.n4246 out.n4245 0.019
R80706 out.n4218 out.n4217 0.019
R80707 out.n4312 out.n4311 0.019
R80708 out.n4281 out.n4280 0.019
R80709 out.n4310 out.n4309 0.019
R80710 out.n4377 out.n4376 0.019
R80711 out.n4440 out.n4439 0.019
R80712 out.n4413 out.n4412 0.019
R80713 out.n4505 out.n4504 0.019
R80714 out.n4477 out.n4476 0.019
R80715 out.n4503 out.n4502 0.019
R80716 out.n4569 out.n4568 0.019
R80717 out.n4636 out.n4635 0.019
R80718 out.n4608 out.n4607 0.019
R80719 out.n4698 out.n4697 0.019
R80720 out.n4672 out.n4671 0.019
R80721 out.n4762 out.n4761 0.019
R80722 out.n4736 out.n4735 0.019
R80723 out.n4833 out.n4832 0.019
R80724 out.n4799 out.n4798 0.019
R80725 out.n61 out.n60 0.019
R80726 out.n63 out.n62 0.019
R80727 out.n22 out.n21 0.019
R80728 out.n124 out.n123 0.019
R80729 out.n126 out.n125 0.019
R80730 out.n190 out.n189 0.019
R80731 out.n192 out.n191 0.019
R80732 out.n256 out.n255 0.019
R80733 out.n318 out.n317 0.019
R80734 out.n320 out.n319 0.019
R80735 out.n284 out.n283 0.019
R80736 out.n386 out.n385 0.019
R80737 out.n448 out.n447 0.019
R80738 out.n450 out.n449 0.019
R80739 out.n417 out.n416 0.019
R80740 out.n488 out.n486 0.019
R80741 out.n576 out.n575 0.019
R80742 out.n544 out.n543 0.019
R80743 out.n550 out.n548 0.019
R80744 out.n642 out.n641 0.019
R80745 out.n644 out.n643 0.019
R80746 out.n709 out.n708 0.019
R80747 out.n711 out.n710 0.019
R80748 out.n772 out.n771 0.019
R80749 out.n742 out.n740 0.019
R80750 out.n805 out.n804 0.019
R80751 out.n4915 out.n4914 0.019
R80752 out.n4913 out.n4912 0.019
R80753 out.n869 out.n868 0.019
R80754 out.n4031 out.n4030 0.019
R80755 out.n4033 out.n4032 0.019
R80756 out.n4097 out.n4096 0.019
R80757 out.n4099 out.n4098 0.019
R80758 out.n4160 out.n4159 0.019
R80759 out.n4162 out.n4161 0.019
R80760 out.n4224 out.n4223 0.019
R80761 out.n4226 out.n4225 0.019
R80762 out.n4287 out.n4286 0.019
R80763 out.n4289 out.n4288 0.019
R80764 out.n4353 out.n4352 0.019
R80765 out.n4355 out.n4354 0.019
R80766 out.n4391 out.n4390 0.019
R80767 out.n4483 out.n4482 0.019
R80768 out.n4452 out.n4451 0.019
R80769 out.n4457 out.n4456 0.019
R80770 out.n4546 out.n4545 0.019
R80771 out.n4613 out.n4612 0.019
R80772 out.n4615 out.n4614 0.019
R80773 out.n4580 out.n4579 0.019
R80774 out.n4678 out.n4677 0.019
R80775 out.n4741 out.n4740 0.019
R80776 out.n4743 out.n4742 0.019
R80777 out.n4708 out.n4707 0.019
R80778 out.n4806 out.n4805 0.019
R80779 out.n6757 out.n6752 0.018
R80780 out.n12277 out.n12276 0.018
R80781 out.n12275 out.n12273 0.018
R80782 out.n12162 out.n12161 0.018
R80783 out.n12037 out.n12036 0.018
R80784 out.n13557 out.n13556 0.018
R80785 out.n13555 out.n13553 0.018
R80786 out.n13436 out.n13435 0.018
R80787 out.n13311 out.n13310 0.018
R80788 out.n14012 out.n14011 0.018
R80789 out.n14010 out.n14008 0.018
R80790 out.n13891 out.n13890 0.018
R80791 out.n13766 out.n13765 0.018
R80792 out.n12176 out.n12175 0.018
R80793 out.n13325 out.n13324 0.018
R80794 out.n13780 out.n13779 0.018
R80795 out.n12284 out.n12283 0.018
R80796 out.n13549 out.n13547 0.018
R80797 out.n14004 out.n14002 0.018
R80798 out.n2118 out.n2117 0.018
R80799 out.n1506 out.n1376 0.018
R80800 out.n2353 out.n2220 0.018
R80801 out.n6555 out.n6553 0.018
R80802 out.n6590 out.n6589 0.018
R80803 out.n1582 out.n1580 0.018
R80804 out.n7637 out.n7636 0.018
R80805 out.n7171 out.n7170 0.018
R80806 out.n5772 out.n5770 0.018
R80807 out.n6906 out.n6904 0.018
R80808 out.n12269 out.n12267 0.018
R80809 out.n13564 out.n13563 0.018
R80810 out.n10916 out.n10915 0.018
R80811 out.n10791 out.n10790 0.018
R80812 out.n14019 out.n14018 0.018
R80813 out.n7751 out.n7750 0.018
R80814 out.n11019 out.n11018 0.018
R80815 out.n10909 out.n10908 0.018
R80816 out.n10784 out.n10783 0.018
R80817 out.n7166 out.n7164 0.018
R80818 out.n12051 out.n12050 0.018
R80819 out.n11026 out.n11025 0.018
R80820 out.n2893 out.n2892 0.018
R80821 out.n1797 out.n1796 0.018
R80822 out.n1604 out.n1603 0.018
R80823 out.n13050 out.n13049 0.018
R80824 out.n12923 out.n12922 0.018
R80825 out.n11765 out.n11764 0.018
R80826 out.n11638 out.n11637 0.018
R80827 out.n10498 out.n10497 0.018
R80828 out.n10371 out.n10370 0.018
R80829 out.n6695 out.n6694 0.018
R80830 out.n6020 out.n6019 0.018
R80831 out.n6142 out.n6141 0.018
R80832 out.n2678 out.n2676 0.018
R80833 out.n13450 out.n13449 0.018
R80834 out.n13905 out.n13904 0.018
R80835 out.n5204 out.n5203 0.018
R80836 out.n12730 out.n12729 0.018
R80837 out.n12485 out.n12484 0.018
R80838 out.n11438 out.n11436 0.018
R80839 out.n11343 out.n11342 0.018
R80840 out.n11221 out.n11220 0.018
R80841 out.n11011 out.n11009 0.018
R80842 out.n5321 out.n5320 0.018
R80843 out.n6352 out.n6351 0.018
R80844 out.n5492 out.n5490 0.018
R80845 out.n7350 out.n7348 0.018
R80846 out.n10181 out.n10180 0.018
R80847 out.n13102 out.n13101 0.018
R80848 out.n13166 out.n13161 0.018
R80849 out.n12882 out.n12878 0.018
R80850 out.n13002 out.n13001 0.018
R80851 out.n13067 out.n13062 0.018
R80852 out.n12929 out.n12927 0.018
R80853 out.n12409 out.n12408 0.018
R80854 out.n12413 out.n12412 0.018
R80855 out.n12701 out.n12700 0.018
R80856 out.n12763 out.n12760 0.018
R80857 out.n12445 out.n12441 0.018
R80858 out.n12237 out.n12236 0.018
R80859 out.n12301 out.n12296 0.018
R80860 out.n12015 out.n12011 0.018
R80861 out.n12137 out.n12136 0.018
R80862 out.n12202 out.n12197 0.018
R80863 out.n12064 out.n12062 0.018
R80864 out.n13254 out.n13253 0.018
R80865 out.n13258 out.n13257 0.018
R80866 out.n13535 out.n13534 0.018
R80867 out.n13597 out.n13594 0.018
R80868 out.n13289 out.n13285 0.018
R80869 out.n11411 out.n11410 0.018
R80870 out.n11470 out.n11465 0.018
R80871 out.n11183 out.n11179 0.018
R80872 out.n11311 out.n11310 0.018
R80873 out.n11376 out.n11371 0.018
R80874 out.n11241 out.n11239 0.018
R80875 out.n10984 out.n10983 0.018
R80876 out.n11043 out.n11038 0.018
R80877 out.n10757 out.n10753 0.018
R80878 out.n10884 out.n10883 0.018
R80879 out.n10949 out.n10944 0.018
R80880 out.n10811 out.n10809 0.018
R80881 out.n11817 out.n11816 0.018
R80882 out.n11881 out.n11876 0.018
R80883 out.n11597 out.n11593 0.018
R80884 out.n11717 out.n11716 0.018
R80885 out.n11782 out.n11777 0.018
R80886 out.n11644 out.n11642 0.018
R80887 out.n13709 out.n13708 0.018
R80888 out.n13713 out.n13712 0.018
R80889 out.n13990 out.n13989 0.018
R80890 out.n14052 out.n14049 0.018
R80891 out.n13744 out.n13740 0.018
R80892 out.n10550 out.n10549 0.018
R80893 out.n10614 out.n10609 0.018
R80894 out.n10330 out.n10326 0.018
R80895 out.n10450 out.n10449 0.018
R80896 out.n10515 out.n10510 0.018
R80897 out.n10377 out.n10375 0.018
R80898 out.n14204 out.n14203 0.018
R80899 out.n14342 out.n14341 0.018
R80900 out.n14321 out.n14316 0.018
R80901 out.n14379 out.n14374 0.018
R80902 out.n15564 out.n15383 0.018
R80903 out.n15905 out.n15376 0.018
R80904 out.n5029 out.n5028 0.018
R80905 out.n5008 out.n5003 0.018
R80906 out.n992 out.n991 0.018
R80907 out.n1014 out.n1013 0.018
R80908 out.n5068 out.n5063 0.018
R80909 out.n955 out.n952 0.018
R80910 out.n5856 out.n5855 0.018
R80911 out.n5763 out.n5762 0.018
R80912 out.n5648 out.n5647 0.018
R80913 out.n5739 out.n5738 0.018
R80914 out.n5727 out.n5726 0.018
R80915 out.n5726 out.n5721 0.018
R80916 out.n5653 out.n5649 0.018
R80917 out.n2863 out.n2861 0.018
R80918 out.n2838 out.n2837 0.018
R80919 out.n2846 out.n2845 0.018
R80920 out.n2822 out.n2821 0.018
R80921 out.n2755 out.n2753 0.018
R80922 out.n1413 out.n1412 0.018
R80923 out.n5485 out.n5480 0.018
R80924 out.n5621 out.n5620 0.018
R80925 out.n5347 out.n5342 0.018
R80926 out.n5210 out.n5208 0.018
R80927 out.n1199 out.n1198 0.018
R80928 out.n1176 out.n1173 0.018
R80929 out.n6529 out.n6525 0.018
R80930 out.n6649 out.n6644 0.018
R80931 out.n6763 out.n6762 0.018
R80932 out.n6428 out.n6427 0.018
R80933 out.n6340 out.n6339 0.018
R80934 out.n6225 out.n6224 0.018
R80935 out.n6316 out.n6315 0.018
R80936 out.n6304 out.n6303 0.018
R80937 out.n6303 out.n6298 0.018
R80938 out.n6230 out.n6226 0.018
R80939 out.n1987 out.n1985 0.018
R80940 out.n1962 out.n1961 0.018
R80941 out.n1970 out.n1969 0.018
R80942 out.n1946 out.n1945 0.018
R80943 out.n1884 out.n1882 0.018
R80944 out.n6159 out.n6154 0.018
R80945 out.n6099 out.n6096 0.018
R80946 out.n5899 out.n5895 0.018
R80947 out.n6026 out.n6024 0.018
R80948 out.n5970 out.n5966 0.018
R80949 out.n2979 out.n2978 0.018
R80950 out.n2982 out.n2980 0.018
R80951 out.n6990 out.n6989 0.018
R80952 out.n6897 out.n6896 0.018
R80953 out.n6782 out.n6781 0.018
R80954 out.n6873 out.n6872 0.018
R80955 out.n6861 out.n6860 0.018
R80956 out.n6860 out.n6855 0.018
R80957 out.n6787 out.n6783 0.018
R80958 out.n1767 out.n1765 0.018
R80959 out.n1742 out.n1741 0.018
R80960 out.n1750 out.n1749 0.018
R80961 out.n1726 out.n1725 0.018
R80962 out.n1659 out.n1657 0.018
R80963 out.n2257 out.n2256 0.018
R80964 out.n7343 out.n7338 0.018
R80965 out.n7016 out.n7015 0.018
R80966 out.n2394 out.n2393 0.018
R80967 out.n7177 out.n7175 0.018
R80968 out.n7051 out.n7047 0.018
R80969 out.n7069 out.n7067 0.018
R80970 out.n2486 out.n2485 0.018
R80971 out.n2469 out.n2468 0.018
R80972 out.n2460 out.n2459 0.018
R80973 out.n7723 out.n7722 0.018
R80974 out.n7498 out.n7497 0.018
R80975 out.n7507 out.n7506 0.018
R80976 out.n7517 out.n7516 0.018
R80977 out.n7516 out.n7511 0.018
R80978 out.n7523 out.n7519 0.018
R80979 out.n7627 out.n7626 0.018
R80980 out.n7560 out.n7559 0.018
R80981 out.n7557 out.n7551 0.018
R80982 out.n7601 out.n7597 0.018
R80983 out.n2633 out.n2631 0.018
R80984 out.n9438 out.n9426 0.018
R80985 out.n2917 out.n2782 0.018
R80986 out.n1297 out.n1178 0.018
R80987 out.n1821 out.n1686 0.018
R80988 out.n1111 out.n1110 0.018
R80989 out.n12603 out.n12602 0.018
R80990 out.n12478 out.n12477 0.018
R80991 out.n11336 out.n11335 0.018
R80992 out.n11214 out.n11213 0.018
R80993 out.n11017 out.n11015 0.018
R80994 out.n1248 out.n1247 0.018
R80995 out.n5315 out.n5314 0.018
R80996 out.n5313 out.n5311 0.018
R80997 out.n12492 out.n12491 0.018
R80998 out.n10923 out.n10922 0.018
R80999 out.n10798 out.n10797 0.018
R81000 out.n5534 out.n5533 0.018
R81001 out.n5330 out.n5329 0.018
R81002 out.n6359 out.n6358 0.018
R81003 out.n7392 out.n7391 0.018
R81004 out.n12715 out.n12713 0.018
R81005 out.n12610 out.n12609 0.018
R81006 out.n11453 out.n11452 0.018
R81007 out.n12058 out.n12057 0.018
R81008 out.n13332 out.n13331 0.018
R81009 out.n13787 out.n13786 0.018
R81010 out.n7054 out.n7053 0.018
R81011 out.n1048 out.n1047 0.018
R81012 out.n1102 out.n1101 0.018
R81013 out.n6683 out.n6681 0.018
R81014 out.n5780 out.n5779 0.018
R81015 out.n6914 out.n6913 0.018
R81016 out.n1082 out.n961 0.018
R81017 out.n2041 out.n1906 0.018
R81018 out.n12723 out.n12722 0.018
R81019 out.n12721 out.n12719 0.018
R81020 out.n11446 out.n11445 0.018
R81021 out.n11444 out.n11442 0.018
R81022 out.n11350 out.n11349 0.018
R81023 out.n11228 out.n11227 0.018
R81024 out.n5787 out.n5786 0.018
R81025 out.n6921 out.n6920 0.018
R81026 out.n14565 out.n14564 0.018
R81027 out.n12185 out.n12184 0.017
R81028 out.n13459 out.n13458 0.017
R81029 out.n13914 out.n13913 0.017
R81030 out.n6233 out.n6232 0.017
R81031 out.n7180 out.n7179 0.017
R81032 out.n13434 out.n13432 0.017
R81033 out.n13310 out.n13308 0.017
R81034 out.n13889 out.n13887 0.017
R81035 out.n13765 out.n13763 0.017
R81036 out.n8879 out.n8877 0.017
R81037 out.n12617 out.n12616 0.017
R81038 out.n14436 out.n14330 0.017
R81039 out.n5110 out.n5017 0.017
R81040 out.n2557 out.n2555 0.017
R81041 out.n1494 out.n1398 0.017
R81042 out.n2341 out.n2242 0.017
R81043 out.n13158 out.n13157 0.017
R81044 out.n11873 out.n11872 0.017
R81045 out.n10606 out.n10605 0.017
R81046 out.n2140 out.n2138 0.017
R81047 out.n1575 out.n1573 0.017
R81048 out.n8879 out.n8873 0.017
R81049 out.n8879 out.n8874 0.017
R81050 out.n8879 out.n8876 0.017
R81051 out.n7630 out.n7628 0.017
R81052 out.n7726 out.n7724 0.017
R81053 out.n10932 out.n10931 0.017
R81054 out.n10805 out.n10804 0.017
R81055 out.n5213 out.n5212 0.017
R81056 out.n6597 out.n6596 0.017
R81057 out.n6548 out.n6546 0.017
R81058 out.n7646 out.n7645 0.017
R81059 out.n7607 out.n7605 0.017
R81060 out.n5796 out.n5795 0.017
R81061 out.n6368 out.n6367 0.017
R81062 out.n6930 out.n6929 0.017
R81063 out.n12293 out.n12292 0.017
R81064 out.n13540 out.n13538 0.017
R81065 out.n13995 out.n13993 0.017
R81066 out.n5418 out.n5414 0.017
R81067 out.n2947 out.n2946 0.017
R81068 out.n3190 out.n3188 0.017
R81069 out.n2949 out.n2945 0.017
R81070 out.n6487 out.n6483 0.017
R81071 out.n7279 out.n7275 0.017
R81072 out.n2596 out.n2595 0.017
R81073 out.n2598 out.n2594 0.017
R81074 out.n3253 out.n3243 0.017
R81075 out.n13025 out.n13023 0.017
R81076 out.n12901 out.n12899 0.017
R81077 out.n11740 out.n11738 0.017
R81078 out.n11616 out.n11614 0.017
R81079 out.n10473 out.n10471 0.017
R81080 out.n10349 out.n10347 0.017
R81081 out.n6008 out.n6006 0.017
R81082 out.n6122 out.n6120 0.017
R81083 out.n12601 out.n12599 0.017
R81084 out.n12477 out.n12475 0.017
R81085 out.n5519 out.n5517 0.017
R81086 out.n7377 out.n7375 0.017
R81087 out.n12626 out.n12625 0.017
R81088 out.n12499 out.n12498 0.017
R81089 out.n11359 out.n11358 0.017
R81090 out.n11235 out.n11234 0.017
R81091 out.n5656 out.n5655 0.017
R81092 out.n5541 out.n5540 0.017
R81093 out.n6790 out.n6789 0.017
R81094 out.n7399 out.n7398 0.017
R81095 out.n12932 out.n12931 0.017
R81096 out.n11647 out.n11646 0.017
R81097 out.n10380 out.n10379 0.017
R81098 out.n6704 out.n6703 0.017
R81099 out.n6642 out.n6640 0.017
R81100 out.n6029 out.n6028 0.017
R81101 out.n7760 out.n7759 0.017
R81102 out.n2671 out.n2669 0.017
R81103 out.n15421 out.n15419 0.017
R81104 out.n2971 out.n2970 0.017
R81105 out.n5976 out.n5974 0.017
R81106 out.n11035 out.n11034 0.017
R81107 out.n2541 out.n2540 0.017
R81108 out.n8879 out.n8878 0.017
R81109 out.n7063 out.n7062 0.017
R81110 out.n8879 out.n8875 0.017
R81111 out.n12706 out.n12704 0.016
R81112 out.n11462 out.n11461 0.016
R81113 out.n12160 out.n12158 0.016
R81114 out.n12036 out.n12034 0.016
R81115 out.n13426 out.n13424 0.016
R81116 out.n13304 out.n13302 0.016
R81117 out.n13881 out.n13879 0.016
R81118 out.n13759 out.n13757 0.016
R81119 out.n6677 out.n6675 0.016
R81120 out.n13127 out.n13125 0.016
R81121 out.n13017 out.n13015 0.016
R81122 out.n12895 out.n12894 0.016
R81123 out.n11842 out.n11840 0.016
R81124 out.n11732 out.n11730 0.016
R81125 out.n11610 out.n11609 0.016
R81126 out.n10575 out.n10573 0.016
R81127 out.n10465 out.n10463 0.016
R81128 out.n10343 out.n10342 0.016
R81129 out.n6002 out.n6000 0.016
R81130 out.n6114 out.n6112 0.016
R81131 out.n12067 out.n12066 0.016
R81132 out.n13341 out.n13340 0.016
R81133 out.n13796 out.n13795 0.016
R81134 out.n5222 out.n5221 0.016
R81135 out.n2026 out.n2025 0.016
R81136 out.n7189 out.n7188 0.016
R81137 out.n1251 out.n1250 0.016
R81138 out.n5306 out.n5304 0.016
R81139 out.n2526 out.n2525 0.016
R81140 out.n7160 out.n7158 0.016
R81141 out.n15413 out.n15410 0.016
R81142 out.n2887 out.n2886 0.016
R81143 out.n5766 out.n5764 0.016
R81144 out.n2011 out.n2010 0.016
R81145 out.n6343 out.n6341 0.016
R81146 out.n1791 out.n1790 0.016
R81147 out.n6900 out.n6898 0.016
R81148 out.n11334 out.n11332 0.016
R81149 out.n11213 out.n11211 0.016
R81150 out.n10907 out.n10905 0.016
R81151 out.n10783 out.n10781 0.016
R81152 out.n7717 out.n7715 0.016
R81153 out.n11244 out.n11243 0.016
R81154 out.n10814 out.n10813 0.016
R81155 out.n2902 out.n2901 0.016
R81156 out.n5478 out.n5476 0.016
R81157 out.n6242 out.n6241 0.016
R81158 out.n6377 out.n6376 0.016
R81159 out.n1806 out.n1805 0.016
R81160 out.n7336 out.n7334 0.016
R81161 out.n2915 out.n2791 0.016
R81162 out.n1504 out.n1383 0.016
R81163 out.n1819 out.n1695 0.016
R81164 out.n2351 out.n2227 0.016
R81165 out.n15421 out.n15420 0.016
R81166 out.n9674 out.n9673 0.016
R81167 out.n9473 out.n9472 0.016
R81168 out.n5339 out.n5338 0.016
R81169 out.n10101 out.n10100 0.016
R81170 out.n12593 out.n12591 0.016
R81171 out.n12471 out.n12469 0.016
R81172 out.n5513 out.n5511 0.016
R81173 out.n7371 out.n7369 0.016
R81174 out.n12262 out.n12260 0.016
R81175 out.n12152 out.n12150 0.016
R81176 out.n12030 out.n12028 0.016
R81177 out.n13571 out.n13570 0.016
R81178 out.n11004 out.n11002 0.016
R81179 out.n10899 out.n10897 0.016
R81180 out.n10777 out.n10775 0.016
R81181 out.n14026 out.n14025 0.016
R81182 out.n1080 out.n965 0.016
R81183 out.n1295 out.n1183 0.016
R81184 out.n2039 out.n1915 0.016
R81185 out.n12508 out.n12507 0.016
R81186 out.n5665 out.n5664 0.016
R81187 out.n5805 out.n5804 0.016
R81188 out.n5550 out.n5549 0.016
R81189 out.n6799 out.n6798 0.016
R81190 out.n6939 out.n6938 0.016
R81191 out.n7408 out.n7407 0.016
R81192 out.n10121 out.n10120 0.016
R81193 out.n2544 out.n2543 0.016
R81194 out.n2726 out.n2724 0.015
R81195 out.n2554 out.n2552 0.015
R81196 out.n1589 out.n1587 0.015
R81197 out.n6436 out.n6435 0.015
R81198 out.n12737 out.n12736 0.015
R81199 out.n11431 out.n11429 0.015
R81200 out.n11326 out.n11324 0.015
R81201 out.n11207 out.n11205 0.015
R81202 out.n6606 out.n6605 0.015
R81203 out.n6545 out.n6543 0.015
R81204 out.n5973 out.n5972 0.015
R81205 out.n11559 out.n11558 0.015
R81206 out.n13059 out.n13058 0.015
R81207 out.n11774 out.n11773 0.015
R81208 out.n10507 out.n10506 0.015
R81209 out.n6151 out.n6150 0.015
R81210 out.n5757 out.n5755 0.015
R81211 out.n6334 out.n6332 0.015
R81212 out.n6891 out.n6889 0.015
R81213 out.n2131 out.n2129 0.015
R81214 out.n1572 out.n1570 0.015
R81215 out.n7699 out.n7697 0.015
R81216 out.n2685 out.n2683 0.015
R81217 out.n9672 out.n9671 0.015
R81218 out.n3194 out.n3191 0.015
R81219 out.n3247 out.n3245 0.015
R81220 out.n7604 out.n7603 0.015
R81221 out.n12975 out.n12973 0.015
R81222 out.n12943 out.n12942 0.015
R81223 out.n11690 out.n11688 0.015
R81224 out.n11658 out.n11657 0.015
R81225 out.n10423 out.n10421 0.015
R81226 out.n10391 out.n10390 0.015
R81227 out.n6713 out.n6712 0.015
R81228 out.n6639 out.n6637 0.015
R81229 out.n6040 out.n6039 0.015
R81230 out.n6078 out.n6076 0.015
R81231 out.n7655 out.n7654 0.015
R81232 out.n2668 out.n2666 0.015
R81233 out.n12194 out.n12193 0.015
R81234 out.n7151 out.n7149 0.015
R81235 out.n1616 out.n1614 0.015
R81236 out.n12110 out.n12108 0.015
R81237 out.n13381 out.n13379 0.015
R81238 out.n13836 out.n13834 0.015
R81239 out.n7115 out.n7113 0.015
R81240 out.n10941 out.n10940 0.015
R81241 out.n1254 out.n1253 0.015
R81242 out.n5297 out.n5295 0.015
R81243 out.n14104 out.n10288 0.014
R81244 out.n12078 out.n12077 0.014
R81245 out.n13350 out.n13349 0.014
R81246 out.n10857 out.n10855 0.014
R81247 out.n13805 out.n13804 0.014
R81248 out.n1266 out.n1265 0.014
R81249 out.n6251 out.n6250 0.014
R81250 out.n6296 out.n6294 0.014
R81251 out.n7072 out.n7071 0.014
R81252 out.n11368 out.n11367 0.014
R81253 out.n12397 out.n12396 0.014
R81254 out.n10709 out.n10290 0.014
R81255 out.n11136 out.n11135 0.014
R81256 out.n13169 out.n13168 0.014
R81257 out.n12304 out.n12303 0.014
R81258 out.n13529 out.n13527 0.014
R81259 out.n13415 out.n13413 0.014
R81260 out.n11884 out.n11883 0.014
R81261 out.n13984 out.n13982 0.014
R81262 out.n13870 out.n13868 0.014
R81263 out.n10617 out.n10616 0.014
R81264 out.n1508 out.n1369 0.014
R81265 out.n2355 out.n2213 0.014
R81266 out.n14494 out.n14270 0.014
R81267 out.n14434 out.n14339 0.014
R81268 out.n5108 out.n5026 0.014
R81269 out.n12548 out.n12546 0.014
R81270 out.n12517 out.n12516 0.014
R81271 out.n11287 out.n11285 0.014
R81272 out.n10825 out.n10824 0.014
R81273 out.n5719 out.n5717 0.014
R81274 out.n5559 out.n5558 0.014
R81275 out.n5475 out.n5473 0.014
R81276 out.n6853 out.n6851 0.014
R81277 out.n7417 out.n7416 0.014
R81278 out.n7333 out.n7331 0.014
R81279 out.n9446 ldomc_0.vdm_0.vout 0.014
R81280 out.n10067 out.n10066 0.014
R81281 out.n10186 out.n10181 0.014
R81282 out.n10105 out.n10102 0.014
R81283 out.n13123 out.n13122 0.014
R81284 out.n13122 out.n13121 0.014
R81285 out.n13131 out.n13130 0.014
R81286 out.n13153 out.n13150 0.014
R81287 out.n12982 out.n12977 0.014
R81288 out.n13022 out.n13021 0.014
R81289 out.n13038 out.n13035 0.014
R81290 out.n12898 out.n12897 0.014
R81291 out.n12913 out.n12910 0.014
R81292 out.n12946 out.n12945 0.014
R81293 out.n12712 out.n12711 0.014
R81294 out.n12734 out.n12731 0.014
R81295 out.n12745 out.n12740 0.014
R81296 out.n12740 out.n12739 0.014
R81297 out.n12589 out.n12588 0.014
R81298 out.n12614 out.n12611 0.014
R81299 out.n12645 out.n12640 0.014
R81300 out.n12489 out.n12486 0.014
R81301 out.n12505 out.n12503 0.014
R81302 out.n11983 out.n11982 0.014
R81303 out.n12258 out.n12257 0.014
R81304 out.n12257 out.n12256 0.014
R81305 out.n12266 out.n12265 0.014
R81306 out.n12288 out.n12285 0.014
R81307 out.n12117 out.n12112 0.014
R81308 out.n12157 out.n12156 0.014
R81309 out.n12173 out.n12170 0.014
R81310 out.n12033 out.n12032 0.014
R81311 out.n12048 out.n12045 0.014
R81312 out.n12081 out.n12080 0.014
R81313 out.n13546 out.n13545 0.014
R81314 out.n13568 out.n13565 0.014
R81315 out.n13579 out.n13574 0.014
R81316 out.n13574 out.n13573 0.014
R81317 out.n13422 out.n13421 0.014
R81318 out.n13447 out.n13444 0.014
R81319 out.n13478 out.n13473 0.014
R81320 out.n13322 out.n13319 0.014
R81321 out.n13338 out.n13336 0.014
R81322 out.n11143 out.n11142 0.014
R81323 out.n11427 out.n11426 0.014
R81324 out.n11426 out.n11425 0.014
R81325 out.n11435 out.n11434 0.014
R81326 out.n11457 out.n11454 0.014
R81327 out.n11294 out.n11289 0.014
R81328 out.n11331 out.n11330 0.014
R81329 out.n11347 out.n11344 0.014
R81330 out.n11210 out.n11209 0.014
R81331 out.n11225 out.n11222 0.014
R81332 out.n11258 out.n11257 0.014
R81333 out.n10720 out.n10719 0.014
R81334 out.n11000 out.n10999 0.014
R81335 out.n10999 out.n10998 0.014
R81336 out.n11008 out.n11007 0.014
R81337 out.n11030 out.n11027 0.014
R81338 out.n10864 out.n10859 0.014
R81339 out.n10904 out.n10903 0.014
R81340 out.n10920 out.n10917 0.014
R81341 out.n10780 out.n10779 0.014
R81342 out.n10795 out.n10792 0.014
R81343 out.n10828 out.n10827 0.014
R81344 out.n11566 out.n11565 0.014
R81345 out.n11838 out.n11837 0.014
R81346 out.n11837 out.n11836 0.014
R81347 out.n11846 out.n11845 0.014
R81348 out.n11868 out.n11865 0.014
R81349 out.n11697 out.n11692 0.014
R81350 out.n11737 out.n11736 0.014
R81351 out.n11753 out.n11750 0.014
R81352 out.n11613 out.n11612 0.014
R81353 out.n11628 out.n11625 0.014
R81354 out.n11661 out.n11660 0.014
R81355 out.n14001 out.n14000 0.014
R81356 out.n14023 out.n14020 0.014
R81357 out.n14034 out.n14029 0.014
R81358 out.n14029 out.n14028 0.014
R81359 out.n13877 out.n13876 0.014
R81360 out.n13902 out.n13899 0.014
R81361 out.n13933 out.n13928 0.014
R81362 out.n13777 out.n13774 0.014
R81363 out.n13793 out.n13791 0.014
R81364 out.n10299 out.n10298 0.014
R81365 out.n10571 out.n10570 0.014
R81366 out.n10570 out.n10569 0.014
R81367 out.n10579 out.n10578 0.014
R81368 out.n10601 out.n10598 0.014
R81369 out.n10430 out.n10425 0.014
R81370 out.n10470 out.n10469 0.014
R81371 out.n10486 out.n10483 0.014
R81372 out.n10346 out.n10345 0.014
R81373 out.n10361 out.n10358 0.014
R81374 out.n10394 out.n10393 0.014
R81375 out.n14267 out.n14266 0.014
R81376 out.n14502 out.n14501 0.014
R81377 out.n14236 out.n14235 0.014
R81378 out.n14328 out.n14327 0.014
R81379 out.n14327 out.n14326 0.014
R81380 out.n14440 out.n14439 0.014
R81381 out.n14462 out.n14459 0.014
R81382 out.n14169 out.n14167 0.014
R81383 out.n14407 out.n14404 0.014
R81384 out.n15383 out.n15382 0.014
R81385 out.n15564 out.n15384 0.014
R81386 out.n15366 out.n15365 0.014
R81387 out.n16202 out.n15367 0.014
R81388 out.n14147 out.n14124 0.014
R81389 out.n14634 out.n14612 0.014
R81390 out.n14705 out.n14683 0.014
R81391 out.n14776 out.n14754 0.014
R81392 out.n14847 out.n14825 0.014
R81393 out.n14918 out.n14896 0.014
R81394 out.n14989 out.n14967 0.014
R81395 out.n15054 out.n15032 0.014
R81396 out.n15119 out.n15097 0.014
R81397 out.n15157 out.n15135 0.014
R81398 out.n15198 out.n15175 0.014
R81399 out.n15263 out.n15241 0.014
R81400 out.n15328 out.n15306 0.014
R81401 out.n9015 out.n8992 0.014
R81402 out.n15492 out.n15488 0.014
R81403 out.n16263 out.n16260 0.014
R81404 out.n17277 out.n17274 0.014
R81405 out.n16166 out.n16163 0.014
R81406 out.n16105 out.n16102 0.014
R81407 out.n15978 out.n15975 0.014
R81408 out.n16014 out.n16011 0.014
R81409 out.n15869 out.n15866 0.014
R81410 out.n15808 out.n15805 0.014
R81411 out.n15747 out.n15744 0.014
R81412 out.n15676 out.n15673 0.014
R81413 out.n15605 out.n15602 0.014
R81414 out.n15528 out.n15525 0.014
R81415 out.n15455 out.n15453 0.014
R81416 out.n5015 out.n5014 0.014
R81417 out.n5014 out.n5013 0.014
R81418 out.n5114 out.n5113 0.014
R81419 out.n5136 out.n5133 0.014
R81420 out.n1001 out.n1000 0.014
R81421 out.n1030 out.n1028 0.014
R81422 out.n1036 out.n1035 0.014
R81423 out.n946 out.n944 0.014
R81424 out.n1091 out.n1090 0.014
R81425 out.n963 out.n962 0.014
R81426 out.n2738 out.n2736 0.014
R81427 out.n5808 out.n5807 0.014
R81428 out.n5793 out.n5791 0.014
R81429 out.n5784 out.n5781 0.014
R81430 out.n5671 out.n5669 0.014
R81431 out.n2873 out.n2872 0.014
R81432 out.n2813 out.n2812 0.014
R81433 out.n2759 out.n2758 0.014
R81434 out.n1344 out.n1343 0.014
R81435 out.n1346 out.n1344 0.014
R81436 out.n1440 out.n1439 0.014
R81437 out.n1431 out.n1430 0.014
R81438 out.n1458 out.n1457 0.014
R81439 out.n5448 out.n5447 0.014
R81440 out.n5547 out.n5545 0.014
R81441 out.n5531 out.n5528 0.014
R81442 out.n5487 out.n5486 0.014
R81443 out.n1360 out.n1359 0.014
R81444 out.n5389 out.n5388 0.014
R81445 out.n5607 out.n5390 0.014
R81446 out.n1533 out.n1532 0.014
R81447 out.n1147 out.n1146 0.014
R81448 out.n5342 out.n5341 0.014
R81449 out.n5325 out.n5322 0.014
R81450 out.n5260 out.n5255 0.014
R81451 out.n5201 out.n5198 0.014
R81452 out.n1236 out.n1234 0.014
R81453 out.n1223 out.n1220 0.014
R81454 out.n1209 out.n1208 0.014
R81455 out.n1216 out.n1210 0.014
R81456 out.n1217 out.n1216 0.014
R81457 out.n1206 out.n1201 0.014
R81458 out.n1310 out.n1309 0.014
R81459 out.n1334 out.n1139 0.014
R81460 out.n2080 out.n2079 0.014
R81461 out.n2082 out.n2080 0.014
R81462 out.n6510 out.n6505 0.014
R81463 out.n6518 out.n6514 0.014
R81464 out.n6580 out.n6577 0.014
R81465 out.n6493 out.n6492 0.014
R81466 out.n6701 out.n6699 0.014
R81467 out.n6463 out.n6460 0.014
R81468 out.n6651 out.n6650 0.014
R81469 out.n2094 out.n2093 0.014
R81470 out.n2106 out.n2105 0.014
R81471 out.n1867 out.n1865 0.014
R81472 out.n6380 out.n6379 0.014
R81473 out.n6365 out.n6363 0.014
R81474 out.n6356 out.n6353 0.014
R81475 out.n6248 out.n6246 0.014
R81476 out.n1997 out.n1996 0.014
R81477 out.n1937 out.n1936 0.014
R81478 out.n1888 out.n1887 0.014
R81479 out.n1544 out.n1542 0.014
R81480 out.n6130 out.n6127 0.014
R81481 out.n6119 out.n6118 0.014
R81482 out.n6085 out.n6080 0.014
R81483 out.n6043 out.n6042 0.014
R81484 out.n5909 out.n5906 0.014
R81485 out.n6005 out.n6004 0.014
R81486 out.n5928 out.n5925 0.014
R81487 out.n1550 out.n1547 0.014
R81488 out.n1560 out.n1559 0.014
R81489 out.n1611 out.n1610 0.014
R81490 out.n1850 out.n1846 0.014
R81491 out.n1642 out.n1640 0.014
R81492 out.n6942 out.n6941 0.014
R81493 out.n6927 out.n6925 0.014
R81494 out.n6918 out.n6915 0.014
R81495 out.n6805 out.n6803 0.014
R81496 out.n1777 out.n1776 0.014
R81497 out.n1717 out.n1716 0.014
R81498 out.n1663 out.n1662 0.014
R81499 out.n2188 out.n2187 0.014
R81500 out.n2190 out.n2188 0.014
R81501 out.n2284 out.n2283 0.014
R81502 out.n2275 out.n2274 0.014
R81503 out.n2302 out.n2301 0.014
R81504 out.n7306 out.n7305 0.014
R81505 out.n7405 out.n7403 0.014
R81506 out.n7389 out.n7386 0.014
R81507 out.n7345 out.n7344 0.014
R81508 out.n2204 out.n2203 0.014
R81509 out.n2380 out.n2379 0.014
R81510 out.n7250 out.n7249 0.014
R81511 out.n7464 out.n7251 0.014
R81512 out.n2396 out.n2394 0.014
R81513 out.n7236 out.n7235 0.014
R81514 out.n7229 out.n7224 0.014
R81515 out.n7034 out.n7031 0.014
R81516 out.n7156 out.n7153 0.014
R81517 out.n7046 out.n7045 0.014
R81518 out.n7137 out.n7136 0.014
R81519 out.n7135 out.n7134 0.014
R81520 out.n7134 out.n7128 0.014
R81521 out.n7123 out.n7122 0.014
R81522 out.n2519 out.n2518 0.014
R81523 out.n2494 out.n2493 0.014
R81524 out.n2416 out.n2415 0.014
R81525 out.n2628 out.n2626 0.014
R81526 out.n7763 out.n7762 0.014
R81527 out.n7748 out.n7746 0.014
R81528 out.n7739 out.n7736 0.014
R81529 out.n7652 out.n7650 0.014
R81530 out.n7535 out.n7532 0.014
R81531 out.n7581 out.n7577 0.014
R81532 out.n7248 out.n7244 0.014
R81533 out.n3984 out.n3980 0.014
R81534 out.n3923 out.n3919 0.014
R81535 out.n3846 out.n3842 0.014
R81536 out.n3769 out.n3765 0.014
R81537 out.n3692 out.n3688 0.014
R81538 out.n3615 out.n3611 0.014
R81539 out.n3538 out.n3534 0.014
R81540 out.n3461 out.n3457 0.014
R81541 out.n3384 out.n3380 0.014
R81542 out.n3307 out.n3303 0.014
R81543 out.n3150 out.n3142 0.014
R81544 out.n3023 out.n3016 0.014
R81545 out.n1128 out.n936 0.014
R81546 out.n15406 out.n15405 0.014
R81547 out.n15400 out.n15399 0.014
R81548 out.n12827 out.n12826 0.014
R81549 out.n13674 out.n13673 0.014
R81550 out.n14101 out.n14100 0.014
R81551 out.n11046 out.n11045 0.014
R81552 out.n5860 out.n5859 0.014
R81553 out.n11255 out.n11254 0.014
R81554 out.n5674 out.n5673 0.014
R81555 out.n6808 out.n6807 0.014
R81556 out.n15432 out.n15430 0.014
R81557 out.n15430 out.n15429 0.014
R81558 out.n1609 out.n1607 0.014
R81559 out.n15402 out.n15401 0.014
R81560 out.n13116 out.n13114 0.013
R81561 out.n13006 out.n13004 0.013
R81562 out.n11831 out.n11829 0.013
R81563 out.n11721 out.n11719 0.013
R81564 out.n10564 out.n10562 0.013
R81565 out.n10454 out.n10452 0.013
R81566 out.n6103 out.n6101 0.013
R81567 out.n12695 out.n12693 0.013
R81568 out.n12582 out.n12580 0.013
R81569 out.n11473 out.n11472 0.013
R81570 out.n2147 out.n2145 0.013
R81571 out.n10271 out.n10270 0.013
R81572 out.n12805 out.n12411 0.013
R81573 out.n14103 out.n13248 0.013
R81574 out.n14598 out.n14589 0.013
R81575 out.n14634 out.n14624 0.013
R81576 out.n14669 out.n14660 0.013
R81577 out.n14705 out.n14695 0.013
R81578 out.n14740 out.n14731 0.013
R81579 out.n14776 out.n14766 0.013
R81580 out.n14811 out.n14802 0.013
R81581 out.n14847 out.n14837 0.013
R81582 out.n14882 out.n14873 0.013
R81583 out.n14918 out.n14908 0.013
R81584 out.n14953 out.n14944 0.013
R81585 out.n14989 out.n14979 0.013
R81586 out.n15021 out.n15012 0.013
R81587 out.n15054 out.n15044 0.013
R81588 out.n15086 out.n15077 0.013
R81589 out.n15119 out.n15109 0.013
R81590 out.n15157 out.n15147 0.013
R81591 out.n15198 out.n15188 0.013
R81592 out.n15229 out.n15220 0.013
R81593 out.n15263 out.n15253 0.013
R81594 out.n15294 out.n15285 0.013
R81595 out.n15328 out.n15318 0.013
R81596 out.n15359 out.n15350 0.013
R81597 out.n9015 out.n9005 0.013
R81598 out.n16266 out.n16265 0.013
R81599 out.n16235 out.n16234 0.013
R81600 out.n16199 out.n16198 0.013
R81601 out.n16169 out.n16168 0.013
R81602 out.n16138 out.n16137 0.013
R81603 out.n16108 out.n16107 0.013
R81604 out.n16077 out.n16076 0.013
R81605 out.n15938 out.n15937 0.013
R81606 out.n15902 out.n15901 0.013
R81607 out.n15872 out.n15871 0.013
R81608 out.n15841 out.n15840 0.013
R81609 out.n15811 out.n15810 0.013
R81610 out.n15780 out.n15779 0.013
R81611 out.n15750 out.n15749 0.013
R81612 out.n15714 out.n15713 0.013
R81613 out.n15679 out.n15678 0.013
R81614 out.n15643 out.n15642 0.013
R81615 out.n15561 out.n15560 0.013
R81616 out.n15531 out.n15530 0.013
R81617 out.n15495 out.n15494 0.013
R81618 out.n15459 out.n15458 0.013
R81619 out.n14103 out.n12401 0.013
R81620 out.n16263 out.n16254 0.013
R81621 out.n16231 out.n16224 0.013
R81622 out.n17277 out.n17268 0.013
R81623 out.n16196 out.n16189 0.013
R81624 out.n16166 out.n16157 0.013
R81625 out.n16135 out.n16128 0.013
R81626 out.n16105 out.n16096 0.013
R81627 out.n16073 out.n16066 0.013
R81628 out.n15978 out.n15969 0.013
R81629 out.n15935 out.n15928 0.013
R81630 out.n16014 out.n16005 0.013
R81631 out.n15899 out.n15892 0.013
R81632 out.n15869 out.n15860 0.013
R81633 out.n15838 out.n15831 0.013
R81634 out.n15808 out.n15799 0.013
R81635 out.n15777 out.n15770 0.013
R81636 out.n15747 out.n15738 0.013
R81637 out.n15711 out.n15704 0.013
R81638 out.n15676 out.n15667 0.013
R81639 out.n15639 out.n15632 0.013
R81640 out.n15605 out.n15596 0.013
R81641 out.n15558 out.n15551 0.013
R81642 out.n15528 out.n15519 0.013
R81643 out.n15492 out.n15483 0.013
R81644 out.n2939 out.n2934 0.013
R81645 out.n3162 out.n3161 0.013
R81646 out.n6447 out.n6205 0.013
R81647 out.n2068 out.n2063 0.013
R81648 out.n1843 out.n1838 0.013
R81649 out.n2591 out.n2586 0.013
R81650 out.n2619 out.n2615 0.013
R81651 out.n7820 out.n7012 0.013
R81652 out.n7859 out.n7847 0.013
R81653 out.n7897 out.n7887 0.013
R81654 out.n7936 out.n7924 0.013
R81655 out.n7974 out.n7964 0.013
R81656 out.n8013 out.n8001 0.013
R81657 out.n8051 out.n8041 0.013
R81658 out.n8090 out.n8078 0.013
R81659 out.n8128 out.n8118 0.013
R81660 out.n8167 out.n8155 0.013
R81661 out.n8205 out.n8195 0.013
R81662 out.n8244 out.n8232 0.013
R81663 out.n8282 out.n8272 0.013
R81664 out.n8321 out.n8309 0.013
R81665 out.n8359 out.n8349 0.013
R81666 out.n8398 out.n8386 0.013
R81667 out.n8436 out.n8426 0.013
R81668 out.n8475 out.n8463 0.013
R81669 out.n8513 out.n8503 0.013
R81670 out.n8552 out.n8540 0.013
R81671 out.n8590 out.n8580 0.013
R81672 out.n8629 out.n8617 0.013
R81673 out.n8667 out.n8657 0.013
R81674 out.n8706 out.n8694 0.013
R81675 out.n8744 out.n8734 0.013
R81676 out.n8792 out.n8777 0.013
R81677 out.n907 out.n899 0.013
R81678 out.n3948 out.n3937 0.013
R81679 out.n3910 out.n3899 0.013
R81680 out.n3871 out.n3860 0.013
R81681 out.n3833 out.n3822 0.013
R81682 out.n3794 out.n3783 0.013
R81683 out.n3756 out.n3745 0.013
R81684 out.n3717 out.n3706 0.013
R81685 out.n3679 out.n3668 0.013
R81686 out.n3640 out.n3629 0.013
R81687 out.n3602 out.n3591 0.013
R81688 out.n3563 out.n3552 0.013
R81689 out.n3525 out.n3514 0.013
R81690 out.n3486 out.n3475 0.013
R81691 out.n3448 out.n3437 0.013
R81692 out.n3409 out.n3398 0.013
R81693 out.n3371 out.n3360 0.013
R81694 out.n3332 out.n3321 0.013
R81695 out.n3294 out.n3283 0.013
R81696 out.n3238 out.n3207 0.013
R81697 out.n3150 out.n3123 0.013
R81698 out.n3121 out.n3091 0.013
R81699 out.n3057 out.n3046 0.013
R81700 out.n2996 out.n2976 0.013
R81701 out.n2943 out.n2184 0.013
R81702 out.n2180 out.n1633 0.013
R81703 out.n6766 out.n6449 0.013
R81704 out.n7844 out.n7843 0.013
R81705 out.n7884 out.n7881 0.013
R81706 out.n7921 out.n7920 0.013
R81707 out.n7961 out.n7958 0.013
R81708 out.n7998 out.n7997 0.013
R81709 out.n8038 out.n8035 0.013
R81710 out.n8075 out.n8074 0.013
R81711 out.n8115 out.n8112 0.013
R81712 out.n8152 out.n8151 0.013
R81713 out.n8192 out.n8189 0.013
R81714 out.n8229 out.n8228 0.013
R81715 out.n8269 out.n8266 0.013
R81716 out.n8306 out.n8305 0.013
R81717 out.n8346 out.n8343 0.013
R81718 out.n8383 out.n8382 0.013
R81719 out.n8423 out.n8420 0.013
R81720 out.n8460 out.n8459 0.013
R81721 out.n8500 out.n8497 0.013
R81722 out.n8537 out.n8536 0.013
R81723 out.n8577 out.n8574 0.013
R81724 out.n8614 out.n8613 0.013
R81725 out.n8654 out.n8651 0.013
R81726 out.n8691 out.n8690 0.013
R81727 out.n8731 out.n8728 0.013
R81728 out.n8774 out.n8771 0.013
R81729 out.n907 out.n906 0.013
R81730 out.n3948 out.n3947 0.013
R81731 out.n3910 out.n3909 0.013
R81732 out.n3871 out.n3870 0.013
R81733 out.n3833 out.n3832 0.013
R81734 out.n3794 out.n3793 0.013
R81735 out.n3756 out.n3755 0.013
R81736 out.n3717 out.n3716 0.013
R81737 out.n3679 out.n3678 0.013
R81738 out.n3640 out.n3639 0.013
R81739 out.n3602 out.n3601 0.013
R81740 out.n3563 out.n3562 0.013
R81741 out.n3525 out.n3524 0.013
R81742 out.n3486 out.n3485 0.013
R81743 out.n3448 out.n3447 0.013
R81744 out.n3409 out.n3408 0.013
R81745 out.n3371 out.n3370 0.013
R81746 out.n3332 out.n3331 0.013
R81747 out.n3294 out.n3293 0.013
R81748 out.n3238 out.n3237 0.013
R81749 out.n3113 out.n3111 0.013
R81750 out.n3118 out.n3104 0.013
R81751 out.n3121 out.n3120 0.013
R81752 out.n3057 out.n3056 0.013
R81753 out.n2996 out.n2995 0.013
R81754 out.n2172 out.n2072 0.013
R81755 out.n2180 out.n2179 0.013
R81756 out.n7823 out.n5617 0.013
R81757 out.n7862 out.n7828 0.013
R81758 out.n7900 out.n7868 0.013
R81759 out.n7939 out.n7905 0.013
R81760 out.n7977 out.n7945 0.013
R81761 out.n8016 out.n7982 0.013
R81762 out.n8054 out.n8022 0.013
R81763 out.n8093 out.n8059 0.013
R81764 out.n8131 out.n8099 0.013
R81765 out.n8170 out.n8136 0.013
R81766 out.n8208 out.n8176 0.013
R81767 out.n8247 out.n8213 0.013
R81768 out.n8285 out.n8253 0.013
R81769 out.n8324 out.n8290 0.013
R81770 out.n8362 out.n8330 0.013
R81771 out.n8401 out.n8367 0.013
R81772 out.n8439 out.n8407 0.013
R81773 out.n8478 out.n8444 0.013
R81774 out.n8516 out.n8484 0.013
R81775 out.n8555 out.n8521 0.013
R81776 out.n8593 out.n8561 0.013
R81777 out.n8632 out.n8598 0.013
R81778 out.n8670 out.n8638 0.013
R81779 out.n8709 out.n8675 0.013
R81780 out.n8747 out.n8715 0.013
R81781 out.n8794 out.n8752 0.013
R81782 out.n3991 out.n3990 0.013
R81783 out.n3968 out.n3967 0.013
R81784 out.n3930 out.n3929 0.013
R81785 out.n3891 out.n3890 0.013
R81786 out.n3853 out.n3852 0.013
R81787 out.n3814 out.n3813 0.013
R81788 out.n3776 out.n3775 0.013
R81789 out.n3737 out.n3736 0.013
R81790 out.n3699 out.n3698 0.013
R81791 out.n3660 out.n3659 0.013
R81792 out.n3622 out.n3621 0.013
R81793 out.n3583 out.n3582 0.013
R81794 out.n3545 out.n3544 0.013
R81795 out.n3506 out.n3505 0.013
R81796 out.n3468 out.n3467 0.013
R81797 out.n3429 out.n3428 0.013
R81798 out.n3391 out.n3390 0.013
R81799 out.n3352 out.n3351 0.013
R81800 out.n3314 out.n3313 0.013
R81801 out.n3275 out.n3274 0.013
R81802 out.n3198 out.n3197 0.013
R81803 out.n3183 out.n3182 0.013
R81804 out.n3157 out.n3156 0.013
R81805 out.n3077 out.n3076 0.013
R81806 out.n3039 out.n3038 0.013
R81807 out.n2952 out.n1138 0.013
R81808 out.n2957 out.n2956 0.013
R81809 out.n7821 out.n5865 0.013
R81810 out.n7860 out.n7832 0.013
R81811 out.n7898 out.n7872 0.013
R81812 out.n7937 out.n7909 0.013
R81813 out.n7975 out.n7949 0.013
R81814 out.n8014 out.n7986 0.013
R81815 out.n8052 out.n8026 0.013
R81816 out.n8091 out.n8063 0.013
R81817 out.n8129 out.n8103 0.013
R81818 out.n8168 out.n8140 0.013
R81819 out.n8206 out.n8180 0.013
R81820 out.n8245 out.n8217 0.013
R81821 out.n8283 out.n8257 0.013
R81822 out.n8322 out.n8294 0.013
R81823 out.n8360 out.n8334 0.013
R81824 out.n8399 out.n8371 0.013
R81825 out.n8437 out.n8411 0.013
R81826 out.n8476 out.n8448 0.013
R81827 out.n8514 out.n8488 0.013
R81828 out.n8553 out.n8525 0.013
R81829 out.n8591 out.n8565 0.013
R81830 out.n8630 out.n8602 0.013
R81831 out.n8668 out.n8642 0.013
R81832 out.n8707 out.n8679 0.013
R81833 out.n8745 out.n8719 0.013
R81834 out.n8793 out.n8758 0.013
R81835 out.n3984 out.n3978 0.013
R81836 out.n3961 out.n3955 0.013
R81837 out.n3923 out.n3917 0.013
R81838 out.n3884 out.n3878 0.013
R81839 out.n3846 out.n3840 0.013
R81840 out.n3807 out.n3801 0.013
R81841 out.n3769 out.n3763 0.013
R81842 out.n3730 out.n3724 0.013
R81843 out.n3692 out.n3686 0.013
R81844 out.n3653 out.n3647 0.013
R81845 out.n3615 out.n3609 0.013
R81846 out.n3576 out.n3570 0.013
R81847 out.n3538 out.n3532 0.013
R81848 out.n3499 out.n3493 0.013
R81849 out.n3461 out.n3455 0.013
R81850 out.n3422 out.n3416 0.013
R81851 out.n3384 out.n3378 0.013
R81852 out.n3345 out.n3339 0.013
R81853 out.n3307 out.n3301 0.013
R81854 out.n3268 out.n3260 0.013
R81855 out.n3177 out.n3167 0.013
R81856 out.n3176 out.n3170 0.013
R81857 out.n3150 out.n3140 0.013
R81858 out.n3070 out.n3064 0.013
R81859 out.n3023 out.n3012 0.013
R81860 out.n2944 out.n1537 0.013
R81861 out.n2943 out.n2614 0.013
R81862 out.n12251 out.n12249 0.013
R81863 out.n12141 out.n12139 0.013
R81864 out.n13582 out.n13581 0.013
R81865 out.n13470 out.n13469 0.013
R81866 out.n14037 out.n14036 0.013
R81867 out.n13925 out.n13924 0.013
R81868 out.n15487 out.n15486 0.013
R81869 out.n14141 out.n14140 0.013
R81870 out.n16258 out.n16257 0.013
R81871 out.n17272 out.n17271 0.013
R81872 out.n16161 out.n16160 0.013
R81873 out.n16100 out.n16099 0.013
R81874 out.n15973 out.n15972 0.013
R81875 out.n16009 out.n16008 0.013
R81876 out.n15864 out.n15863 0.013
R81877 out.n15803 out.n15802 0.013
R81878 out.n15742 out.n15741 0.013
R81879 out.n15671 out.n15670 0.013
R81880 out.n15600 out.n15599 0.013
R81881 out.n15523 out.n15522 0.013
R81882 out.n14145 out.n14144 0.013
R81883 out.n14632 out.n14631 0.013
R81884 out.n14703 out.n14702 0.013
R81885 out.n14774 out.n14773 0.013
R81886 out.n14845 out.n14844 0.013
R81887 out.n14916 out.n14915 0.013
R81888 out.n14987 out.n14986 0.013
R81889 out.n15052 out.n15051 0.013
R81890 out.n15117 out.n15116 0.013
R81891 out.n15155 out.n15154 0.013
R81892 out.n15196 out.n15195 0.013
R81893 out.n15261 out.n15260 0.013
R81894 out.n15326 out.n15325 0.013
R81895 out.n9013 out.n9012 0.013
R81896 out.n15396 out.n15395 0.013
R81897 out.n3022 out.n3020 0.013
R81898 out.n2942 out.n2729 0.013
R81899 out.n1620 out.n1619 0.013
R81900 out.n2606 out.n2604 0.013
R81901 out.n3006 out.n3005 0.013
R81902 out.n3138 out.n3136 0.013
R81903 out.n3255 out.n3254 0.013
R81904 out.n8785 out.n8783 0.013
R81905 out.n8700 out.n8698 0.013
R81906 out.n8623 out.n8621 0.013
R81907 out.n8546 out.n8544 0.013
R81908 out.n8469 out.n8467 0.013
R81909 out.n8392 out.n8390 0.013
R81910 out.n8315 out.n8313 0.013
R81911 out.n8238 out.n8236 0.013
R81912 out.n8161 out.n8159 0.013
R81913 out.n8084 out.n8082 0.013
R81914 out.n8007 out.n8005 0.013
R81915 out.n7930 out.n7928 0.013
R81916 out.n7853 out.n7851 0.013
R81917 out.n7474 out.n7472 0.013
R81918 out.n2600 out.n2599 0.013
R81919 out.n2723 out.n2718 0.013
R81920 out.n7818 out.n7477 0.013
R81921 out.n3250 out.n3248 0.013
R81922 out.n7468 out.n7467 0.013
R81923 out.n2387 out.n2386 0.013
R81924 out.n6197 out.n6196 0.013
R81925 out.n3089 out.n3088 0.013
R81926 out.n1626 out.n1625 0.013
R81927 out.n2715 out.n2620 0.013
R81928 out.n15404 out.n15403 0.013
R81929 out.n15424 out.n15423 0.013
R81930 out.n12748 out.n12747 0.013
R81931 out.n12637 out.n12636 0.013
R81932 out.n11420 out.n11418 0.013
R81933 out.n11315 out.n11313 0.013
R81934 out.n10993 out.n10991 0.013
R81935 out.n10888 out.n10886 0.013
R81936 out.n14110 out.n14109 0.013
R81937 out.n15408 out.n15407 0.012
R81938 out.n5716 out.n5715 0.012
R81939 out.n2913 out.n2798 0.012
R81940 out.n5472 out.n5471 0.012
R81941 out.n1502 out.n1390 0.012
R81942 out.n6850 out.n6849 0.012
R81943 out.n1817 out.n1702 0.012
R81944 out.n7330 out.n7329 0.012
R81945 out.n2349 out.n2234 0.012
R81946 out.n2993 out.n2992 0.012
R81947 out.n2720 out.n2719 0.012
R81948 out.n1349 out.n1348 0.012
R81949 out.n6749 out.n6748 0.012
R81950 out.n2193 out.n2192 0.012
R81951 out.n2399 out.n2398 0.012
R81952 out.n6293 out.n6292 0.012
R81953 out.n2037 out.n1922 0.012
R81954 out.n14428 out.n14362 0.012
R81955 out.n5102 out.n5051 0.012
R81956 out.n7112 out.n7111 0.012
R81957 out.n13639 out.n13256 0.012
R81958 out.n14094 out.n13711 0.012
R81959 out.n15426 out.n15416 0.012
R81960 out.n2941 out.n2940 0.012
R81961 out.n1333 out.n1325 0.012
R81962 out.n2070 out.n2069 0.012
R81963 out.n1845 out.n1844 0.012
R81964 out.n2712 out.n2711 0.012
R81965 out.n9457 out.n9456 0.012
R81966 out.n9000 out.n8999 0.012
R81967 out.n15346 out.n15345 0.012
R81968 out.n15314 out.n15313 0.012
R81969 out.n15281 out.n15280 0.012
R81970 out.n15249 out.n15248 0.012
R81971 out.n15216 out.n15215 0.012
R81972 out.n15183 out.n15182 0.012
R81973 out.n8950 out.n8949 0.012
R81974 out.n15143 out.n15142 0.012
R81975 out.n8913 out.n8912 0.012
R81976 out.n15105 out.n15104 0.012
R81977 out.n15073 out.n15072 0.012
R81978 out.n15040 out.n15039 0.012
R81979 out.n15008 out.n15007 0.012
R81980 out.n14975 out.n14974 0.012
R81981 out.n14940 out.n14939 0.012
R81982 out.n14904 out.n14903 0.012
R81983 out.n14869 out.n14868 0.012
R81984 out.n14833 out.n14832 0.012
R81985 out.n14798 out.n14797 0.012
R81986 out.n14762 out.n14761 0.012
R81987 out.n14727 out.n14726 0.012
R81988 out.n14691 out.n14690 0.012
R81989 out.n14656 out.n14655 0.012
R81990 out.n14620 out.n14619 0.012
R81991 out.n14583 out.n14582 0.012
R81992 out.n1857 out.n1856 0.012
R81993 out.n3100 out.n3099 0.012
R81994 out.n6203 out.n6202 0.012
R81995 out.n3218 out.n3217 0.012
R81996 out.n2984 out.n2983 0.012
R81997 out.n1852 out.n1851 0.012
R81998 out.n7247 out.n7245 0.012
R81999 out.n2551 out.n2443 0.012
R82000 out.n15459 out.n15390 0.012
R82001 out.n8872 out.n5 0.012
R82002 out.n6542 out.n6540 0.012
R82003 out.n6636 out.n6635 0.012
R82004 out.n2128 out.n2124 0.012
R82005 out.n5965 out.n5964 0.012
R82006 out.n7596 out.n7594 0.012
R82007 out.n2710 out.n2708 0.012
R82008 out.n6075 out.n6074 0.012
R82009 out.n17181 out.n17179 0.011
R82010 out.n13206 out.n13205 0.011
R82011 out.n11921 out.n11920 0.011
R82012 out.n10654 out.n10653 0.011
R82013 out.n6618 out.n6617 0.011
R82014 out.n1569 out.n1564 0.011
R82015 out.n7696 out.n7695 0.011
R82016 out.n2665 out.n2663 0.011
R82017 out.n17150 out.n17148 0.011
R82018 out.n13085 out.n13083 0.011
R82019 out.n12972 out.n12970 0.011
R82020 out.n11800 out.n11798 0.011
R82021 out.n11687 out.n11685 0.011
R82022 out.n10533 out.n10531 0.011
R82023 out.n10420 out.n10418 0.011
R82024 out.n3993 out.n3992 0.011
R82025 out.n14110 out.n14106 0.011
R82026 out.n12341 out.n12340 0.011
R82027 out.n13499 out.n13497 0.011
R82028 out.n13954 out.n13952 0.011
R82029 out.n2546 out.n2545 0.011
R82030 out.n7222 out.n7220 0.011
R82031 out.n12220 out.n12218 0.011
R82032 out.n12107 out.n12105 0.011
R82033 out.n13617 out.n13616 0.011
R82034 out.n13378 out.n13376 0.011
R82035 out.n14072 out.n14071 0.011
R82036 out.n13833 out.n13831 0.011
R82037 out.n2702 out.n2701 0.011
R82038 out.n17173 out.n17172 0.011
R82039 out.n15909 out.n15908 0.011
R82040 out.n3232 out.n3228 0.011
R82041 out.n3040 out.n933 0.011
R82042 out.n3158 out.n932 0.011
R82043 out.n3079 out.n3078 0.011
R82044 out.n3199 out.n931 0.011
R82045 out.n3185 out.n3184 0.011
R82046 out.n3315 out.n930 0.011
R82047 out.n3277 out.n3276 0.011
R82048 out.n3392 out.n929 0.011
R82049 out.n3354 out.n3353 0.011
R82050 out.n3469 out.n928 0.011
R82051 out.n3431 out.n3430 0.011
R82052 out.n3546 out.n927 0.011
R82053 out.n3508 out.n3507 0.011
R82054 out.n3623 out.n926 0.011
R82055 out.n3585 out.n3584 0.011
R82056 out.n3700 out.n925 0.011
R82057 out.n3662 out.n3661 0.011
R82058 out.n3777 out.n924 0.011
R82059 out.n3739 out.n3738 0.011
R82060 out.n3854 out.n923 0.011
R82061 out.n3816 out.n3815 0.011
R82062 out.n3931 out.n922 0.011
R82063 out.n3893 out.n3892 0.011
R82064 out.n3970 out.n3969 0.011
R82065 out.n8712 out.n8711 0.011
R82066 out.n8749 out.n4943 0.011
R82067 out.n8635 out.n8634 0.011
R82068 out.n8672 out.n4944 0.011
R82069 out.n8558 out.n8557 0.011
R82070 out.n8595 out.n4945 0.011
R82071 out.n8481 out.n8480 0.011
R82072 out.n8518 out.n4946 0.011
R82073 out.n8404 out.n8403 0.011
R82074 out.n8441 out.n4947 0.011
R82075 out.n8327 out.n8326 0.011
R82076 out.n8364 out.n4948 0.011
R82077 out.n8250 out.n8249 0.011
R82078 out.n8287 out.n4949 0.011
R82079 out.n8173 out.n8172 0.011
R82080 out.n8210 out.n4950 0.011
R82081 out.n8096 out.n8095 0.011
R82082 out.n8133 out.n4951 0.011
R82083 out.n8019 out.n8018 0.011
R82084 out.n8056 out.n4952 0.011
R82085 out.n7942 out.n7941 0.011
R82086 out.n7979 out.n4953 0.011
R82087 out.n7865 out.n7864 0.011
R82088 out.n7902 out.n4954 0.011
R82089 out.n5614 out.n5613 0.011
R82090 out.n7825 out.n4955 0.011
R82091 out.n1134 out.n1133 0.011
R82092 out.n11083 out.n11082 0.011
R82093 out.n5253 out.n5251 0.011
R82094 out.n2032 out.n2031 0.011
R82095 out.n10115 out.n10114 0.011
R82096 out.n10123 out.n10122 0.011
R82097 out.n12868 out.n12864 0.011
R82098 out.n13177 out.n13172 0.011
R82099 out.n13199 out.n13198 0.011
R82100 out.n13186 out.n13184 0.011
R82101 out.n13184 out.n13181 0.011
R82102 out.n13212 out.n13211 0.011
R82103 out.n12888 out.n12884 0.011
R82104 out.n12984 out.n12983 0.011
R82105 out.n13047 out.n13045 0.011
R82106 out.n12805 out.n12804 0.011
R82107 out.n12434 out.n12430 0.011
R82108 out.n12681 out.n12680 0.011
R82109 out.n12680 out.n12677 0.011
R82110 out.n12670 out.n12668 0.011
R82111 out.n12690 out.n12689 0.011
R82112 out.n12789 out.n12788 0.011
R82113 out.n12556 out.n12550 0.011
R82114 out.n12559 out.n12558 0.011
R82115 out.n12588 out.n12587 0.011
R82116 out.n12598 out.n12597 0.011
R82117 out.n12474 out.n12473 0.011
R82118 out.n12001 out.n11997 0.011
R82119 out.n12312 out.n12307 0.011
R82120 out.n12334 out.n12333 0.011
R82121 out.n12321 out.n12319 0.011
R82122 out.n12319 out.n12316 0.011
R82123 out.n12347 out.n12346 0.011
R82124 out.n12021 out.n12017 0.011
R82125 out.n12119 out.n12118 0.011
R82126 out.n12182 out.n12180 0.011
R82127 out.n13639 out.n13638 0.011
R82128 out.n13278 out.n13274 0.011
R82129 out.n13515 out.n13514 0.011
R82130 out.n13514 out.n13511 0.011
R82131 out.n13503 out.n13501 0.011
R82132 out.n13524 out.n13523 0.011
R82133 out.n13623 out.n13622 0.011
R82134 out.n13389 out.n13383 0.011
R82135 out.n13392 out.n13391 0.011
R82136 out.n13421 out.n13420 0.011
R82137 out.n13431 out.n13430 0.011
R82138 out.n13654 out.n13651 0.011
R82139 out.n13307 out.n13306 0.011
R82140 out.n11536 out.n11145 0.011
R82141 out.n11166 out.n11162 0.011
R82142 out.n11481 out.n11476 0.011
R82143 out.n11503 out.n11502 0.011
R82144 out.n11490 out.n11488 0.011
R82145 out.n11488 out.n11485 0.011
R82146 out.n11516 out.n11515 0.011
R82147 out.n11189 out.n11185 0.011
R82148 out.n11296 out.n11295 0.011
R82149 out.n11356 out.n11354 0.011
R82150 out.n11109 out.n10722 0.011
R82151 out.n10743 out.n10739 0.011
R82152 out.n11054 out.n11049 0.011
R82153 out.n11076 out.n11075 0.011
R82154 out.n11063 out.n11061 0.011
R82155 out.n11061 out.n11058 0.011
R82156 out.n11089 out.n11088 0.011
R82157 out.n10763 out.n10759 0.011
R82158 out.n10866 out.n10865 0.011
R82159 out.n10929 out.n10927 0.011
R82160 out.n11583 out.n11579 0.011
R82161 out.n11892 out.n11887 0.011
R82162 out.n11914 out.n11913 0.011
R82163 out.n11901 out.n11899 0.011
R82164 out.n11899 out.n11896 0.011
R82165 out.n11927 out.n11926 0.011
R82166 out.n11603 out.n11599 0.011
R82167 out.n11699 out.n11698 0.011
R82168 out.n11762 out.n11760 0.011
R82169 out.n14094 out.n14093 0.011
R82170 out.n13733 out.n13729 0.011
R82171 out.n13970 out.n13969 0.011
R82172 out.n13969 out.n13966 0.011
R82173 out.n13958 out.n13956 0.011
R82174 out.n13979 out.n13978 0.011
R82175 out.n14078 out.n14077 0.011
R82176 out.n13844 out.n13838 0.011
R82177 out.n13847 out.n13846 0.011
R82178 out.n13876 out.n13875 0.011
R82179 out.n13886 out.n13885 0.011
R82180 out.n13687 out.n13684 0.011
R82181 out.n13762 out.n13761 0.011
R82182 out.n10316 out.n10312 0.011
R82183 out.n10625 out.n10620 0.011
R82184 out.n10647 out.n10646 0.011
R82185 out.n10634 out.n10632 0.011
R82186 out.n10632 out.n10629 0.011
R82187 out.n10660 out.n10659 0.011
R82188 out.n10336 out.n10332 0.011
R82189 out.n10432 out.n10431 0.011
R82190 out.n10495 out.n10493 0.011
R82191 out.n14513 out.n14511 0.011
R82192 out.n14241 out.n14236 0.011
R82193 out.n14207 out.n14206 0.011
R82194 out.n14215 out.n14214 0.011
R82195 out.n14360 out.n14356 0.011
R82196 out.n14312 out.n14307 0.011
R82197 out.n14289 out.n14288 0.011
R82198 out.n14299 out.n14297 0.011
R82199 out.n14297 out.n14295 0.011
R82200 out.n14282 out.n14281 0.011
R82201 out.n14393 out.n14391 0.011
R82202 out.n14555 out.n14553 0.011
R82203 out.n15904 out.n15377 0.011
R82204 out.n15161 out.n10041 0.011
R82205 out.n14103 out.n10713 0.011
R82206 out.n14147 out.n14119 0.011
R82207 out.n14598 out.n14114 0.011
R82208 out.n14634 out.n14604 0.011
R82209 out.n14669 out.n14641 0.011
R82210 out.n14705 out.n14675 0.011
R82211 out.n14740 out.n14712 0.011
R82212 out.n14776 out.n14746 0.011
R82213 out.n14811 out.n14783 0.011
R82214 out.n14847 out.n14817 0.011
R82215 out.n14882 out.n14854 0.011
R82216 out.n14918 out.n14888 0.011
R82217 out.n14953 out.n14925 0.011
R82218 out.n14989 out.n14959 0.011
R82219 out.n15021 out.n14996 0.011
R82220 out.n15054 out.n15027 0.011
R82221 out.n15086 out.n15061 0.011
R82222 out.n15119 out.n15092 0.011
R82223 out.n8929 out.n8901 0.011
R82224 out.n15157 out.n15130 0.011
R82225 out.n8964 out.n8938 0.011
R82226 out.n15198 out.n15170 0.011
R82227 out.n15229 out.n15204 0.011
R82228 out.n15263 out.n15236 0.011
R82229 out.n15294 out.n15269 0.011
R82230 out.n15328 out.n15301 0.011
R82231 out.n15359 out.n15334 0.011
R82232 out.n9015 out.n8987 0.011
R82233 out.n17305 out.n17241 0.011
R82234 out.n17303 out.n17244 0.011
R82235 out.n17300 out.n17246 0.011
R82236 out.n17298 out.n17280 0.011
R82237 out.n17295 out.n17282 0.011
R82238 out.n17293 out.n17285 0.011
R82239 out.n17290 out.n17287 0.011
R82240 out.n16050 out.n15945 0.011
R82241 out.n16047 out.n15947 0.011
R82242 out.n16045 out.n15981 0.011
R82243 out.n16042 out.n15983 0.011
R82244 out.n16040 out.n16017 0.011
R82245 out.n16037 out.n16019 0.011
R82246 out.n16035 out.n16022 0.011
R82247 out.n16032 out.n16024 0.011
R82248 out.n16030 out.n16027 0.011
R82249 out.n15722 out.n15719 0.011
R82250 out.n15688 out.n15685 0.011
R82251 out.n15651 out.n15648 0.011
R82252 out.n15616 out.n15572 0.011
R82253 out.n15613 out.n15574 0.011
R82254 out.n15611 out.n15608 0.011
R82255 out.n15503 out.n15500 0.011
R82256 out.n15468 out.n15465 0.011
R82257 out.n15433 out.n15398 0.011
R82258 out.n5049 out.n5045 0.011
R82259 out.n4999 out.n4994 0.011
R82260 out.n4975 out.n4974 0.011
R82261 out.n4986 out.n4984 0.011
R82262 out.n4984 out.n4981 0.011
R82263 out.n4968 out.n4967 0.011
R82264 out.n985 out.n984 0.011
R82265 out.n995 out.n994 0.011
R82266 out.n5082 out.n5080 0.011
R82267 out.n5849 out.n5844 0.011
R82268 out.n5762 out.n5759 0.011
R82269 out.n5741 out.n5740 0.011
R82270 out.n5740 out.n5739 0.011
R82271 out.n5738 out.n5732 0.011
R82272 out.n2853 out.n2852 0.011
R82273 out.n2827 out.n2823 0.011
R82274 out.n5713 out.n5709 0.011
R82275 out.n5638 out.n5634 0.011
R82276 out.n5596 out.n5595 0.011
R82277 out.n5600 out.n5597 0.011
R82278 out.n1419 out.n1415 0.011
R82279 out.n1453 out.n1450 0.011
R82280 out.n5516 out.n5515 0.011
R82281 out.n5499 out.n5498 0.011
R82282 out.n5407 out.n5406 0.011
R82283 out.n5406 out.n5403 0.011
R82284 out.n5486 out.n5485 0.011
R82285 out.n5413 out.n5412 0.011
R82286 out.n5469 out.n5465 0.011
R82287 out.n1363 out.n1360 0.011
R82288 out.n1375 out.n1374 0.011
R82289 out.n1382 out.n1381 0.011
R82290 out.n1389 out.n1388 0.011
R82291 out.n3035 out.n3034 0.011
R82292 out.n5327 out.n5325 0.011
R82293 out.n5283 out.n5282 0.011
R82294 out.n5282 out.n5280 0.011
R82295 out.n5271 out.n5270 0.011
R82296 out.n5219 out.n5217 0.011
R82297 out.n1192 out.n1191 0.011
R82298 out.n5189 out.n5185 0.011
R82299 out.n6756 out.n6753 0.011
R82300 out.n6524 out.n6523 0.011
R82301 out.n6502 out.n6501 0.011
R82302 out.n6680 out.n6679 0.011
R82303 out.n6663 out.n6662 0.011
R82304 out.n6476 out.n6475 0.011
R82305 out.n6475 out.n6472 0.011
R82306 out.n6650 out.n6649 0.011
R82307 out.n6482 out.n6481 0.011
R82308 out.n6633 out.n6629 0.011
R82309 out.n2097 out.n2094 0.011
R82310 out.n2137 out.n2136 0.011
R82311 out.n2104 out.n2103 0.011
R82312 out.n2111 out.n2110 0.011
R82313 out.n6421 out.n6416 0.011
R82314 out.n6339 out.n6336 0.011
R82315 out.n6318 out.n6317 0.011
R82316 out.n6317 out.n6316 0.011
R82317 out.n6315 out.n6309 0.011
R82318 out.n1977 out.n1976 0.011
R82319 out.n1951 out.n1947 0.011
R82320 out.n6290 out.n6286 0.011
R82321 out.n6210 out.n6206 0.011
R82322 out.n6139 out.n6137 0.011
R82323 out.n6087 out.n6086 0.011
R82324 out.n5985 out.n5984 0.011
R82325 out.n5935 out.n5934 0.011
R82326 out.n5962 out.n5958 0.011
R82327 out.n6072 out.n6068 0.011
R82328 out.n5877 out.n5874 0.011
R82329 out.n6983 out.n6978 0.011
R82330 out.n6896 out.n6893 0.011
R82331 out.n6875 out.n6874 0.011
R82332 out.n6874 out.n6873 0.011
R82333 out.n6872 out.n6866 0.011
R82334 out.n1757 out.n1756 0.011
R82335 out.n1731 out.n1727 0.011
R82336 out.n6847 out.n6843 0.011
R82337 out.n6772 out.n6768 0.011
R82338 out.n7454 out.n7453 0.011
R82339 out.n7458 out.n7455 0.011
R82340 out.n2263 out.n2259 0.011
R82341 out.n2297 out.n2294 0.011
R82342 out.n7374 out.n7373 0.011
R82343 out.n7357 out.n7356 0.011
R82344 out.n7268 out.n7267 0.011
R82345 out.n7267 out.n7264 0.011
R82346 out.n7344 out.n7343 0.011
R82347 out.n7274 out.n7273 0.011
R82348 out.n7327 out.n7323 0.011
R82349 out.n2207 out.n2204 0.011
R82350 out.n2219 out.n2218 0.011
R82351 out.n2226 out.n2225 0.011
R82352 out.n2233 out.n2232 0.011
R82353 out.n2385 out.n2384 0.011
R82354 out.n7186 out.n7184 0.011
R82355 out.n2475 out.n2471 0.011
R82356 out.n7109 out.n7105 0.011
R82357 out.n7022 out.n7018 0.011
R82358 out.n7722 out.n7719 0.011
R82359 out.n7509 out.n7508 0.011
R82360 out.n7508 out.n7507 0.011
R82361 out.n7506 out.n7500 0.011
R82362 out.n7548 out.n7545 0.011
R82363 out.n7575 out.n7574 0.011
R82364 out.n7693 out.n7689 0.011
R82365 out.n7483 out.n7479 0.011
R82366 out.n2604 out.n2603 0.011
R82367 out.n2386 out.n2385 0.011
R82368 out.n1856 out.n1855 0.011
R82369 out.n1625 out.n1624 0.011
R82370 out.n1132 out.n1131 0.011
R82371 out.n2718 out.n2717 0.011
R82372 ldomc_0.out out.n17312 0.011
R82373 out.n10967 out.n10965 0.011
R82374 out.n10854 out.n10852 0.011
R82375 out.n6414 out.n6412 0.011
R82376 out.n15126 out.n15125 0.011
R82377 out.n15939 out.n15373 0.011
R82378 out.n46 out.n45 0.011
R82379 out.n2160 out.n2086 0.011
R82380 out.n15563 out.n15562 0.011
R82381 out.n16201 out.n16200 0.011
R82382 out.n3173 out.n3172 0.011
R82383 out.n9510 out.n9392 0.011
R82384 out.n9546 out.n9358 0.011
R82385 out.n9544 out.n9391 0.011
R82386 out.n9582 out.n9324 0.011
R82387 out.n9580 out.n9357 0.011
R82388 out.n9616 out.n9323 0.011
R82389 out.n9677 out.n9257 0.011
R82390 out.n9675 out.n9290 0.011
R82391 out.n9619 out.n9618 0.011
R82392 out.n9713 out.n9223 0.011
R82393 out.n9711 out.n9256 0.011
R82394 out.n9749 out.n9189 0.011
R82395 out.n9747 out.n9222 0.011
R82396 out.n9785 out.n9155 0.011
R82397 out.n9783 out.n9188 0.011
R82398 out.n9821 out.n9121 0.011
R82399 out.n9819 out.n9154 0.011
R82400 out.n9855 out.n9120 0.011
R82401 out.n9926 out.n9086 0.011
R82402 out.n9892 out.n9087 0.011
R82403 out.n9858 out.n9857 0.011
R82404 out.n9964 out.n9054 0.011
R82405 out.n9962 out.n9085 0.011
R82406 out.n9998 out.n9053 0.011
R82407 out.n17237 out.n16319 0.011
R82408 out.n17239 out.n16286 0.011
R82409 out.n10001 out.n10000 0.011
R82410 out.n17233 out.n16385 0.011
R82411 out.n17235 out.n16352 0.011
R82412 out.n17229 out.n16451 0.011
R82413 out.n17231 out.n16420 0.011
R82414 out.n17225 out.n16517 0.011
R82415 out.n17227 out.n16486 0.011
R82416 out.n17221 out.n16585 0.011
R82417 out.n17223 out.n16550 0.011
R82418 out.n17217 out.n16649 0.011
R82419 out.n17219 out.n16616 0.011
R82420 out.n17213 out.n16715 0.011
R82421 out.n17215 out.n16682 0.011
R82422 out.n17209 out.n16783 0.011
R82423 out.n17211 out.n16748 0.011
R82424 out.n17205 out.n16849 0.011
R82425 out.n17207 out.n16814 0.011
R82426 out.n17201 out.n16913 0.011
R82427 out.n17203 out.n16880 0.011
R82428 out.n17197 out.n16981 0.011
R82429 out.n17199 out.n16946 0.011
R82430 out.n17193 out.n17045 0.011
R82431 out.n17195 out.n17012 0.011
R82432 out.n17189 out.n17111 0.011
R82433 out.n17191 out.n17078 0.011
R82434 out.n17187 out.n17145 0.011
R82435 out.n12666 out.n12664 0.011
R82436 out.n11510 out.n11509 0.011
R82437 out.n2908 out.n2907 0.011
R82438 out.n1812 out.n1811 0.011
R82439 out.n2576 out.n2407 0.011
R82440 out.n15940 out.n15939 0.011
R82441 out.n15126 out.n15122 0.011
R82442 out.n12783 out.n12782 0.011
R82443 out.n12545 out.n12543 0.011
R82444 out.n11394 out.n11392 0.011
R82445 out.n11284 out.n11282 0.011
R82446 out.n5842 out.n5840 0.011
R82447 out.n6976 out.n6974 0.011
R82448 out.n6571 out.n6570 0.011
R82449 out.n9481 out.n9479 0.011
R82450 out.n10179 out.n10178 0.011
R82451 out.n2171 out.n2076 0.011
R82452 out.n4802 out.n4801 0.01
R82453 out.n1108 out.n1107 0.01
R82454 out.n111 out.n110 0.01
R82455 out.n176 out.n175 0.01
R82456 out.n243 out.n242 0.01
R82457 out.n303 out.n302 0.01
R82458 out.n372 out.n371 0.01
R82459 out.n435 out.n434 0.01
R82460 out.n501 out.n500 0.01
R82461 out.n561 out.n560 0.01
R82462 out.n629 out.n628 0.01
R82463 out.n695 out.n694 0.01
R82464 out.n754 out.n753 0.01
R82465 out.n817 out.n816 0.01
R82466 out.n895 out.n894 0.01
R82467 out.n4017 out.n4016 0.01
R82468 out.n4083 out.n4082 0.01
R82469 out.n4144 out.n4143 0.01
R82470 out.n4210 out.n4209 0.01
R82471 out.n4274 out.n4273 0.01
R82472 out.n4338 out.n4337 0.01
R82473 out.n4404 out.n4403 0.01
R82474 out.n4469 out.n4468 0.01
R82475 out.n4531 out.n4530 0.01
R82476 out.n4599 out.n4598 0.01
R82477 out.n4664 out.n4663 0.01
R82478 out.n4728 out.n4727 0.01
R82479 out.n4789 out.n4788 0.01
R82480 out.n1521 out.n1352 0.01
R82481 out.n2368 out.n2196 0.01
R82482 out.n7816 out.n7478 0.01
R82483 out.n17181 out.n17180 0.01
R82484 out.n6765 out.n6761 0.01
R82485 out.n17150 out.n17149 0.01
R82486 out.n9493 out.n9492 0.01
R82487 out.n9498 out.n9495 0.01
R82488 out.n4835 out.n4834 0.01
R82489 out.n1477 out.n1476 0.01
R82490 out.n2324 out.n2323 0.01
R82491 out.n17173 out.n17171 0.01
R82492 out.n3212 out.n3211 0.01
R82493 out.n2157 out.n2156 0.01
R82494 out.n10254 out.n10251 0.01
R82495 out.n10194 out.n10191 0.01
R82496 out.n10170 out.n10169 0.01
R82497 out.n10168 out.n10167 0.01
R82498 out.n10166 out.n10165 0.01
R82499 out.n10146 out.n10145 0.01
R82500 out.n10277 out.n10276 0.01
R82501 out.n13237 out.n13236 0.01
R82502 out.n13237 out.n13235 0.01
R82503 out.n13220 out.n13217 0.01
R82504 out.n13080 out.n13079 0.01
R82505 out.n13243 out.n13242 0.01
R82506 out.n12794 out.n12793 0.01
R82507 out.n12451 out.n12447 0.01
R82508 out.n12661 out.n12659 0.01
R82509 out.n12367 out.n12366 0.01
R82510 out.n12367 out.n11985 0.01
R82511 out.n12355 out.n12352 0.01
R82512 out.n12215 out.n12214 0.01
R82513 out.n12369 out.n12368 0.01
R82514 out.n13628 out.n13627 0.01
R82515 out.n13295 out.n13291 0.01
R82516 out.n13494 out.n13492 0.01
R82517 out.n11524 out.n11521 0.01
R82518 out.n11389 out.n11388 0.01
R82519 out.n11538 out.n11537 0.01
R82520 out.n11097 out.n11094 0.01
R82521 out.n10962 out.n10961 0.01
R82522 out.n11111 out.n11110 0.01
R82523 out.n11947 out.n11946 0.01
R82524 out.n11947 out.n11568 0.01
R82525 out.n11935 out.n11932 0.01
R82526 out.n11795 out.n11794 0.01
R82527 out.n11949 out.n11948 0.01
R82528 out.n14083 out.n14082 0.01
R82529 out.n13750 out.n13746 0.01
R82530 out.n13949 out.n13947 0.01
R82531 out.n10680 out.n10679 0.01
R82532 out.n10680 out.n10301 0.01
R82533 out.n10668 out.n10665 0.01
R82534 out.n10528 out.n10527 0.01
R82535 out.n10682 out.n10681 0.01
R82536 out.n14197 out.n14196 0.01
R82537 out.n14482 out.n14479 0.01
R82538 out.n14424 out.n14423 0.01
R82539 out.n14551 out.n14550 0.01
R82540 out.n15392 out.n15391 0.01
R82541 out.n15568 out.n15567 0.01
R82542 out.n15910 out.n15909 0.01
R82543 out.n16206 out.n16205 0.01
R82544 out.n15164 out.n15163 0.01
R82545 out.n15124 out.n15123 0.01
R82546 out.n14108 out.n14107 0.01
R82547 out.n17265 out.n17264 0.01
R82548 out.n15428 out.n15427 0.01
R82549 out.n5156 out.n5153 0.01
R82550 out.n5098 out.n5097 0.01
R82551 out.n5837 out.n5834 0.01
R82552 out.n5395 out.n5391 0.01
R82553 out.n5248 out.n5247 0.01
R82554 out.n5358 out.n5357 0.01
R82555 out.n5381 out.n5378 0.01
R82556 out.n6454 out.n6450 0.01
R82557 out.n2177 out.n2173 0.01
R82558 out.n6409 out.n6406 0.01
R82559 out.n6172 out.n6171 0.01
R82560 out.n6193 out.n6192 0.01
R82561 out.n6971 out.n6968 0.01
R82562 out.n7256 out.n7252 0.01
R82563 out.n7217 out.n7216 0.01
R82564 out.n7792 out.n7789 0.01
R82565 out.n7471 out.n7470 0.01
R82566 out.n7816 out.n7815 0.01
R82567 out.n7248 out.n7247 0.01
R82568 out.n7464 out.n7463 0.01
R82569 out.n2183 out.n2182 0.01
R82570 out.n7821 out.n5622 0.01
R82571 out.n7823 out.n7822 0.01
R82572 out.n7860 out.n7830 0.01
R82573 out.n7862 out.n7861 0.01
R82574 out.n7898 out.n7870 0.01
R82575 out.n7900 out.n7899 0.01
R82576 out.n7937 out.n7907 0.01
R82577 out.n7939 out.n7938 0.01
R82578 out.n7975 out.n7947 0.01
R82579 out.n7977 out.n7976 0.01
R82580 out.n8014 out.n7984 0.01
R82581 out.n8016 out.n8015 0.01
R82582 out.n8052 out.n8024 0.01
R82583 out.n8054 out.n8053 0.01
R82584 out.n8091 out.n8061 0.01
R82585 out.n8093 out.n8092 0.01
R82586 out.n8129 out.n8101 0.01
R82587 out.n8131 out.n8130 0.01
R82588 out.n8168 out.n8138 0.01
R82589 out.n8170 out.n8169 0.01
R82590 out.n8206 out.n8178 0.01
R82591 out.n8208 out.n8207 0.01
R82592 out.n8245 out.n8215 0.01
R82593 out.n8247 out.n8246 0.01
R82594 out.n8283 out.n8255 0.01
R82595 out.n8285 out.n8284 0.01
R82596 out.n8322 out.n8292 0.01
R82597 out.n8324 out.n8323 0.01
R82598 out.n8360 out.n8332 0.01
R82599 out.n8362 out.n8361 0.01
R82600 out.n8399 out.n8369 0.01
R82601 out.n8401 out.n8400 0.01
R82602 out.n8437 out.n8409 0.01
R82603 out.n8439 out.n8438 0.01
R82604 out.n8476 out.n8446 0.01
R82605 out.n8478 out.n8477 0.01
R82606 out.n8514 out.n8486 0.01
R82607 out.n8516 out.n8515 0.01
R82608 out.n8553 out.n8523 0.01
R82609 out.n8555 out.n8554 0.01
R82610 out.n8591 out.n8563 0.01
R82611 out.n8593 out.n8592 0.01
R82612 out.n8630 out.n8600 0.01
R82613 out.n8632 out.n8631 0.01
R82614 out.n8668 out.n8640 0.01
R82615 out.n8670 out.n8669 0.01
R82616 out.n8707 out.n8677 0.01
R82617 out.n8709 out.n8708 0.01
R82618 out.n8745 out.n8717 0.01
R82619 out.n8747 out.n8746 0.01
R82620 out.n8793 out.n8755 0.01
R82621 out.n3988 out.n3987 0.01
R82622 out.n3965 out.n3964 0.01
R82623 out.n3927 out.n3926 0.01
R82624 out.n3888 out.n3887 0.01
R82625 out.n3850 out.n3849 0.01
R82626 out.n3811 out.n3810 0.01
R82627 out.n3773 out.n3772 0.01
R82628 out.n3734 out.n3733 0.01
R82629 out.n3696 out.n3695 0.01
R82630 out.n3657 out.n3656 0.01
R82631 out.n3619 out.n3618 0.01
R82632 out.n3580 out.n3579 0.01
R82633 out.n3542 out.n3541 0.01
R82634 out.n3503 out.n3502 0.01
R82635 out.n3465 out.n3464 0.01
R82636 out.n3426 out.n3425 0.01
R82637 out.n3388 out.n3387 0.01
R82638 out.n3349 out.n3348 0.01
R82639 out.n3311 out.n3310 0.01
R82640 out.n3272 out.n3271 0.01
R82641 out.n3195 out.n3190 0.01
R82642 out.n3180 out.n3179 0.01
R82643 out.n3154 out.n3153 0.01
R82644 out.n3074 out.n3073 0.01
R82645 out.n3031 out.n3030 0.01
R82646 out.n2944 out.n1340 0.01
R82647 out.n2952 out.n2951 0.01
R82648 out.n1536 out.n1535 0.01
R82649 out.n17312 out 0.01
R82650 out.n7007 out.n7005 0.01
R82651 out.n9481 out.n9480 0.01
R82652 out.n9527 out.n9526 0.01
R82653 out.n9563 out.n9562 0.01
R82654 out.n9380 out.n9379 0.01
R82655 out.n9599 out.n9598 0.01
R82656 out.n9346 out.n9345 0.01
R82657 out.n9638 out.n9637 0.01
R82658 out.n9312 out.n9311 0.01
R82659 out.n9694 out.n9693 0.01
R82660 out.n9279 out.n9278 0.01
R82661 out.n9730 out.n9729 0.01
R82662 out.n9245 out.n9244 0.01
R82663 out.n9766 out.n9765 0.01
R82664 out.n9211 out.n9210 0.01
R82665 out.n9802 out.n9801 0.01
R82666 out.n9177 out.n9176 0.01
R82667 out.n9838 out.n9837 0.01
R82668 out.n9143 out.n9142 0.01
R82669 out.n9877 out.n9876 0.01
R82670 out.n9109 out.n9108 0.01
R82671 out.n9945 out.n9944 0.01
R82672 out.n9912 out.n9911 0.01
R82673 out.n9981 out.n9980 0.01
R82674 out.n9943 out.n9942 0.01
R82675 out.n9042 out.n9041 0.01
R82676 out.n16336 out.n16335 0.01
R82677 out.n16308 out.n16307 0.01
R82678 out.n16404 out.n16403 0.01
R82679 out.n16374 out.n16373 0.01
R82680 out.n16470 out.n16469 0.01
R82681 out.n16402 out.n16401 0.01
R82682 out.n16534 out.n16533 0.01
R82683 out.n16468 out.n16467 0.01
R82684 out.n16638 out.n16637 0.01
R82685 out.n16572 out.n16571 0.01
R82686 out.n16574 out.n16573 0.01
R82687 out.n16704 out.n16703 0.01
R82688 out.n16666 out.n16665 0.01
R82689 out.n16772 out.n16771 0.01
R82690 out.n16732 out.n16731 0.01
R82691 out.n16838 out.n16837 0.01
R82692 out.n16770 out.n16769 0.01
R82693 out.n16902 out.n16901 0.01
R82694 out.n16836 out.n16835 0.01
R82695 out.n16970 out.n16969 0.01
R82696 out.n16930 out.n16929 0.01
R82697 out.n17034 out.n17033 0.01
R82698 out.n16968 out.n16967 0.01
R82699 out.n17100 out.n17099 0.01
R82700 out.n17062 out.n17061 0.01
R82701 out.n17126 out.n17125 0.01
R82702 out.n17128 out.n17127 0.01
R82703 out.n2990 out.n2987 0.01
R82704 out.n1601 out.n1600 0.01
R82705 out.n6193 out.n5867 0.01
R82706 out.n9485 out.n9482 0.01
R82707 out.n4812 out.n4810 0.01
R82708 out.n5286 out.n5284 0.01
R82709 out.n4820 out.n4819 0.01
R82710 out.n9485 out.n9484 0.01
R82711 out.n1518 out.n1517 0.01
R82712 out.n2365 out.n2364 0.01
R82713 out.n14106 out.n14105 0.01
R82714 out.n3053 out.n3052 0.01
R82715 out.n3115 out.n3114 0.01
R82716 out.n3117 out.n3116 0.01
R82717 out.n3328 out.n3327 0.01
R82718 out.n3290 out.n3289 0.01
R82719 out.n3405 out.n3404 0.01
R82720 out.n3367 out.n3366 0.01
R82721 out.n3482 out.n3481 0.01
R82722 out.n3444 out.n3443 0.01
R82723 out.n3559 out.n3558 0.01
R82724 out.n3521 out.n3520 0.01
R82725 out.n3636 out.n3635 0.01
R82726 out.n3598 out.n3597 0.01
R82727 out.n3713 out.n3712 0.01
R82728 out.n3675 out.n3674 0.01
R82729 out.n3790 out.n3789 0.01
R82730 out.n3752 out.n3751 0.01
R82731 out.n3867 out.n3866 0.01
R82732 out.n3829 out.n3828 0.01
R82733 out.n3944 out.n3943 0.01
R82734 out.n3906 out.n3905 0.01
R82735 out.n909 out.n908 0.01
R82736 out.n8730 out.n8729 0.01
R82737 out.n8769 out.n8768 0.01
R82738 out.n8653 out.n8652 0.01
R82739 out.n8688 out.n8687 0.01
R82740 out.n8576 out.n8575 0.01
R82741 out.n8611 out.n8610 0.01
R82742 out.n8499 out.n8498 0.01
R82743 out.n8534 out.n8533 0.01
R82744 out.n8422 out.n8421 0.01
R82745 out.n8457 out.n8456 0.01
R82746 out.n8345 out.n8344 0.01
R82747 out.n8380 out.n8379 0.01
R82748 out.n8268 out.n8267 0.01
R82749 out.n8303 out.n8302 0.01
R82750 out.n8191 out.n8190 0.01
R82751 out.n8226 out.n8225 0.01
R82752 out.n8114 out.n8113 0.01
R82753 out.n8149 out.n8148 0.01
R82754 out.n8037 out.n8036 0.01
R82755 out.n8072 out.n8071 0.01
R82756 out.n7960 out.n7959 0.01
R82757 out.n7995 out.n7994 0.01
R82758 out.n7883 out.n7882 0.01
R82759 out.n7918 out.n7917 0.01
R82760 out.n7841 out.n7840 0.01
R82761 out.n12822 out.n12807 0.009
R82762 out.n15122 out.n15121 0.009
R82763 out.n15941 out.n15940 0.009
R82764 out.n9475 out.n9474 0.009
R82765 out.n16236 out.n15364 0.009
R82766 out.n16078 out.n15370 0.009
R82767 out.n15644 out.n15381 0.009
R82768 out.n15496 out.n15386 0.009
R82769 out.n15461 out.n15460 0.009
R82770 out.n15533 out.n15532 0.009
R82771 out.n15715 out.n15380 0.009
R82772 out.n15681 out.n15680 0.009
R82773 out.n15781 out.n15379 0.009
R82774 out.n15752 out.n15751 0.009
R82775 out.n15842 out.n15378 0.009
R82776 out.n15813 out.n15812 0.009
R82777 out.n15874 out.n15873 0.009
R82778 out.n16139 out.n15369 0.009
R82779 out.n16110 out.n16109 0.009
R82780 out.n16171 out.n16170 0.009
R82781 out.n15362 out.n15361 0.009
R82782 out.n15297 out.n15296 0.009
R82783 out.n15330 out.n10038 0.009
R82784 out.n15232 out.n15231 0.009
R82785 out.n15265 out.n10039 0.009
R82786 out.n15200 out.n10040 0.009
R82787 out.n15057 out.n15056 0.009
R82788 out.n15088 out.n10045 0.009
R82789 out.n14992 out.n14991 0.009
R82790 out.n15023 out.n10046 0.009
R82791 out.n14921 out.n14920 0.009
R82792 out.n14955 out.n10047 0.009
R82793 out.n14850 out.n14849 0.009
R82794 out.n14884 out.n10048 0.009
R82795 out.n14779 out.n14778 0.009
R82796 out.n14813 out.n10049 0.009
R82797 out.n14708 out.n14707 0.009
R82798 out.n14742 out.n10050 0.009
R82799 out.n14637 out.n14636 0.009
R82800 out.n14671 out.n10051 0.009
R82801 out.n14600 out.n10052 0.009
R82802 out.n15164 out.n15162 0.009
R82803 out.n7463 out.n7462 0.009
R82804 out.n9489 out.n9488 0.009
R82805 out.n5611 out.n5387 0.009
R82806 out.n3106 out.n3105 0.009
R82807 ldomc_0.vdm_0.vout out.n9445 0.009
R82808 out.n10248 out.n10247 0.009
R82809 out.n10204 out.n10201 0.009
R82810 out.n12537 out.n12536 0.009
R82811 out.n13370 out.n13369 0.009
R82812 out.n11536 out.n11535 0.009
R82813 out.n11109 out.n11108 0.009
R82814 out.n13825 out.n13824 0.009
R82815 out.n14536 out.n14534 0.009
R82816 out.n14562 out.n14561 0.009
R82817 out.n14560 out.n14557 0.009
R82818 out.n16202 out.n15366 0.009
R82819 out.n15160 out.n10043 0.009
R82820 out.n15966 out.n15965 0.009
R82821 out.n16014 out.n16002 0.009
R82822 out.n15593 out.n15592 0.009
R82823 out.n17311 out.n17310 0.009
R82824 out.n1127 out.n1116 0.009
R82825 out.n5702 out.n5701 0.009
R82826 out.n5828 out.n5827 0.009
R82827 out.n5584 out.n5583 0.009
R82828 out.n1338 out.n1337 0.009
R82829 out.n6738 out.n6737 0.009
R82830 out.n3221 out.n3220 0.009
R82831 out.n6279 out.n6278 0.009
R82832 out.n6400 out.n6399 0.009
R82833 out.n2982 out.n2979 0.009
R82834 out.n3098 out.n3095 0.009
R82835 out.n6201 out.n6200 0.009
R82836 out.n7008 out.n7004 0.009
R82837 out.n6836 out.n6835 0.009
R82838 out.n6962 out.n6961 0.009
R82839 out.n7442 out.n7441 0.009
R82840 out.n2383 out.n2382 0.009
R82841 out.n2593 out.n2592 0.009
R82842 out.n7683 out.n7682 0.009
R82843 out.n7783 out.n7782 0.009
R82844 out.n3015 out.n3014 0.009
R82845 out.n2602 out.n2601 0.009
R82846 out.n3004 out.n3003 0.009
R82847 out.n6999 out.n6998 0.009
R82848 out.n7008 out.n7007 0.009
R82849 out.n6443 out.n6442 0.009
R82850 out.n1129 out.n1128 0.009
R82851 out.n3036 out.n3035 0.009
R82852 out.n5611 out.n5607 0.009
R82853 out.n5625 out.n5624 0.009
R82854 out.n17157 out.n17156 0.009
R82855 out.n9498 out.n9497 0.009
R82856 out.n3175 out.n3174 0.009
R82857 out.n15904 out.n15903 0.009
R82858 out.n15166 out.n15161 0.009
R82859 out.n15502 out.n15501 0.009
R82860 out.n15467 out.n15466 0.009
R82861 out.n15612 out.n15606 0.009
R82862 out.n15610 out.n15609 0.009
R82863 out.n15650 out.n15649 0.009
R82864 out.n15615 out.n15614 0.009
R82865 out.n15721 out.n15720 0.009
R82866 out.n15687 out.n15686 0.009
R82867 out.n16031 out.n16025 0.009
R82868 out.n16029 out.n16028 0.009
R82869 out.n16036 out.n16020 0.009
R82870 out.n16034 out.n16033 0.009
R82871 out.n16041 out.n16015 0.009
R82872 out.n16039 out.n16038 0.009
R82873 out.n16046 out.n15979 0.009
R82874 out.n16044 out.n16043 0.009
R82875 out.n17289 out.n17288 0.009
R82876 out.n16049 out.n16048 0.009
R82877 out.n17294 out.n17283 0.009
R82878 out.n17292 out.n17291 0.009
R82879 out.n17299 out.n17278 0.009
R82880 out.n17297 out.n17296 0.009
R82881 out.n17304 out.n17242 0.009
R82882 out.n17302 out.n17301 0.009
R82883 out.n8977 out.n8976 0.009
R82884 out.n8979 out.n8880 0.009
R82885 out.n8972 out.n8971 0.009
R82886 out.n8974 out.n8881 0.009
R82887 out.n8967 out.n8966 0.009
R82888 out.n8969 out.n8882 0.009
R82889 out.n8932 out.n8931 0.009
R82890 out.n8934 out.n8883 0.009
R82891 out.n8895 out.n8894 0.009
R82892 out.n8897 out.n8884 0.009
R82893 out.n8890 out.n8889 0.009
R82894 out.n8892 out.n8885 0.009
R82895 out.n14961 out.n14960 0.009
R82896 out.n8887 out.n8886 0.009
R82897 out.n14890 out.n14889 0.009
R82898 out.n14927 out.n14926 0.009
R82899 out.n14819 out.n14818 0.009
R82900 out.n14856 out.n14855 0.009
R82901 out.n14748 out.n14747 0.009
R82902 out.n14785 out.n14784 0.009
R82903 out.n14677 out.n14676 0.009
R82904 out.n14714 out.n14713 0.009
R82905 out.n14606 out.n14605 0.009
R82906 out.n14643 out.n14642 0.009
R82907 out.n14568 out.n14567 0.009
R82908 out.n14570 out.n14115 0.009
R82909 out.n3136 out.n3135 0.009
R82910 out.n4812 out.n4811 0.009
R82911 out.n17307 out.n17306 0.009
R82912 out.n17310 out.n8981 0.009
R82913 out.n17153 out.n17152 0.009
R82914 out.n17161 out.n17160 0.009
R82915 out.n9465 out.n9464 0.009
R82916 out.n4820 out.n4818 0.009
R82917 out.n10283 out.n10282 0.008
R82918 out.n15593 out.n15590 0.008
R82919 out.n14136 out.n14135 0.008
R82920 out.n4835 out.n4809 0.008
R82921 out.n5628 out.n5627 0.008
R82922 out.n7002 out.n7001 0.008
R82923 out.n15412 out.n15411 0.008
R82924 out.n10245 out.n10242 0.008
R82925 out.n10238 out.n10235 0.008
R82926 out.n10230 out.n10229 0.008
R82927 out.n13226 out.n13224 0.008
R82928 out.n12964 out.n12963 0.008
R82929 out.n12653 out.n12652 0.008
R82930 out.n12807 out.n12806 0.008
R82931 out.n12361 out.n12359 0.008
R82932 out.n12099 out.n12098 0.008
R82933 out.n13486 out.n13485 0.008
R82934 out.n13641 out.n13640 0.008
R82935 out.n11530 out.n11528 0.008
R82936 out.n11276 out.n11275 0.008
R82937 out.n11103 out.n11101 0.008
R82938 out.n10846 out.n10845 0.008
R82939 out.n11941 out.n11939 0.008
R82940 out.n11679 out.n11678 0.008
R82941 out.n13941 out.n13940 0.008
R82942 out.n14096 out.n14095 0.008
R82943 out.n10674 out.n10672 0.008
R82944 out.n10412 out.n10411 0.008
R82945 out.n14488 out.n14486 0.008
R82946 out.n5162 out.n5160 0.008
R82947 out.n1069 out.n1067 0.008
R82948 out.n5695 out.n5694 0.008
R82949 out.n5243 out.n5242 0.008
R82950 out.n1277 out.n1275 0.008
R82951 out.n6272 out.n6271 0.008
R82952 out.n6062 out.n6061 0.008
R82953 out.n6829 out.n6828 0.008
R82954 out.n7098 out.n7097 0.008
R82955 out.n7212 out.n7211 0.008
R82956 out.n7676 out.n7675 0.008
R82957 out.n3254 out.n3253 0.008
R82958 out.n3247 out.n3246 0.008
R82959 out.n3215 out.n3214 0.008
R82960 out.n2982 out.n2981 0.008
R82961 out.n2969 out.n2968 0.008
R82962 out.n6445 out.n6444 0.008
R82963 out.n5605 out.n5604 0.008
R82964 out.n3194 out.n3193 0.008
R82965 out.n2949 out.n2948 0.008
R82966 out.n3166 out.n3165 0.008
R82967 out.n12392 out.n12369 0.008
R82968 out.n36 out.n35 0.008
R82969 out.n9504 out.n9503 0.008
R82970 out.n40 out.n38 0.008
R82971 out.n22 out.n20 0.008
R82972 out.n18 out.n16 0.008
R82973 out.n43 out.n41 0.008
R82974 out.n13180 out.n13179 0.008
R82975 out.n11895 out.n11894 0.008
R82976 out.n10628 out.n10627 0.008
R82977 out.n12315 out.n12314 0.008
R82978 out.n13518 out.n13516 0.008
R82979 out.n11057 out.n11056 0.008
R82980 out.n13973 out.n13971 0.008
R82981 out.n1325 out.n1323 0.008
R82982 out.n17185 out.n17162 0.008
R82983 out.n17185 out.n17178 0.008
R82984 out.n12684 out.n12682 0.008
R82985 out.n11484 out.n11483 0.008
R82986 out.n7814 out.n7813 0.007
R82987 out.n6757 out.n6756 0.007
R82988 out.n4815 out.n4814 0.007
R82989 out.n30 out.n28 0.007
R82990 out.n55 out.n53 0.007
R82991 out.n5387 out.n5386 0.007
R82992 out.n4831 out.n4830 0.007
R82993 out.n4826 out.n4825 0.007
R82994 out.n4808 out.n4807 0.007
R82995 out.n10228 out.n10227 0.007
R82996 out.n10113 out.n10109 0.007
R82997 out.n10118 out.n10115 0.007
R82998 out.n10089 out.n10088 0.007
R82999 out.n13095 out.n13092 0.007
R83000 out.n13111 out.n13110 0.007
R83001 out.n13137 out.n13136 0.007
R83002 out.n13146 out.n13143 0.007
R83003 out.n13161 out.n13160 0.007
R83004 out.n12990 out.n12987 0.007
R83005 out.n13012 out.n13011 0.007
R83006 out.n13021 out.n13019 0.007
R83007 out.n13031 out.n13028 0.007
R83008 out.n13075 out.n13074 0.007
R83009 out.n12838 out.n12835 0.007
R83010 out.n12839 out.n12838 0.007
R83011 out.n12906 out.n12903 0.007
R83012 out.n12935 out.n12934 0.007
R83013 out.n12800 out.n12798 0.007
R83014 out.n12702 out.n12701 0.007
R83015 out.n12718 out.n12717 0.007
R83016 out.n12727 out.n12724 0.007
R83017 out.n12756 out.n12751 0.007
R83018 out.n12774 out.n12773 0.007
R83019 out.n12780 out.n12779 0.007
R83020 out.n12607 out.n12604 0.007
R83021 out.n12623 out.n12621 0.007
R83022 out.n12629 out.n12628 0.007
R83023 out.n12482 out.n12479 0.007
R83024 out.n12531 out.n12530 0.007
R83025 out.n12230 out.n12227 0.007
R83026 out.n12246 out.n12245 0.007
R83027 out.n12272 out.n12271 0.007
R83028 out.n12281 out.n12278 0.007
R83029 out.n12296 out.n12295 0.007
R83030 out.n12125 out.n12122 0.007
R83031 out.n12147 out.n12146 0.007
R83032 out.n12156 out.n12154 0.007
R83033 out.n12166 out.n12163 0.007
R83034 out.n12210 out.n12209 0.007
R83035 out.n12379 out.n12376 0.007
R83036 out.n12380 out.n12379 0.007
R83037 out.n12041 out.n12038 0.007
R83038 out.n12070 out.n12069 0.007
R83039 out.n13634 out.n13632 0.007
R83040 out.n13536 out.n13535 0.007
R83041 out.n13552 out.n13551 0.007
R83042 out.n13561 out.n13558 0.007
R83043 out.n13590 out.n13585 0.007
R83044 out.n13608 out.n13607 0.007
R83045 out.n13614 out.n13613 0.007
R83046 out.n13440 out.n13437 0.007
R83047 out.n13456 out.n13454 0.007
R83048 out.n13462 out.n13461 0.007
R83049 out.n13315 out.n13312 0.007
R83050 out.n13364 out.n13363 0.007
R83051 out.n11404 out.n11401 0.007
R83052 out.n11441 out.n11440 0.007
R83053 out.n11450 out.n11447 0.007
R83054 out.n11465 out.n11464 0.007
R83055 out.n11302 out.n11299 0.007
R83056 out.n11321 out.n11320 0.007
R83057 out.n11330 out.n11328 0.007
R83058 out.n11340 out.n11337 0.007
R83059 out.n11384 out.n11383 0.007
R83060 out.n11548 out.n11547 0.007
R83061 out.n11218 out.n11215 0.007
R83062 out.n11247 out.n11246 0.007
R83063 out.n10977 out.n10974 0.007
R83064 out.n11014 out.n11013 0.007
R83065 out.n11023 out.n11020 0.007
R83066 out.n11038 out.n11037 0.007
R83067 out.n10872 out.n10869 0.007
R83068 out.n10894 out.n10893 0.007
R83069 out.n10903 out.n10901 0.007
R83070 out.n10913 out.n10910 0.007
R83071 out.n10957 out.n10956 0.007
R83072 out.n11123 out.n11120 0.007
R83073 out.n11124 out.n11123 0.007
R83074 out.n10788 out.n10785 0.007
R83075 out.n10817 out.n10816 0.007
R83076 out.n11810 out.n11807 0.007
R83077 out.n11826 out.n11825 0.007
R83078 out.n11852 out.n11851 0.007
R83079 out.n11861 out.n11858 0.007
R83080 out.n11876 out.n11875 0.007
R83081 out.n11705 out.n11702 0.007
R83082 out.n11727 out.n11726 0.007
R83083 out.n11736 out.n11734 0.007
R83084 out.n11746 out.n11743 0.007
R83085 out.n11790 out.n11789 0.007
R83086 out.n11959 out.n11956 0.007
R83087 out.n11960 out.n11959 0.007
R83088 out.n11621 out.n11618 0.007
R83089 out.n11650 out.n11649 0.007
R83090 out.n14089 out.n14087 0.007
R83091 out.n13991 out.n13990 0.007
R83092 out.n14007 out.n14006 0.007
R83093 out.n14016 out.n14013 0.007
R83094 out.n14045 out.n14040 0.007
R83095 out.n14063 out.n14062 0.007
R83096 out.n14069 out.n14068 0.007
R83097 out.n13895 out.n13892 0.007
R83098 out.n13911 out.n13909 0.007
R83099 out.n13917 out.n13916 0.007
R83100 out.n13770 out.n13767 0.007
R83101 out.n13819 out.n13818 0.007
R83102 out.n10543 out.n10540 0.007
R83103 out.n10559 out.n10558 0.007
R83104 out.n10585 out.n10584 0.007
R83105 out.n10594 out.n10591 0.007
R83106 out.n10609 out.n10608 0.007
R83107 out.n10438 out.n10435 0.007
R83108 out.n10460 out.n10459 0.007
R83109 out.n10469 out.n10467 0.007
R83110 out.n10479 out.n10476 0.007
R83111 out.n10523 out.n10522 0.007
R83112 out.n10692 out.n10689 0.007
R83113 out.n10693 out.n10692 0.007
R83114 out.n10354 out.n10351 0.007
R83115 out.n10383 out.n10382 0.007
R83116 out.n14259 out.n14258 0.007
R83117 out.n14250 out.n14247 0.007
R83118 out.n14245 out.n14244 0.007
R83119 out.n14545 out.n14543 0.007
R83120 out.n14354 out.n14351 0.007
R83121 out.n14336 out.n14335 0.007
R83122 out.n14446 out.n14445 0.007
R83123 out.n14455 out.n14452 0.007
R83124 out.n14316 out.n14315 0.007
R83125 out.n14165 out.n14160 0.007
R83126 out.n14171 out.n14169 0.007
R83127 out.n14400 out.n14397 0.007
R83128 out.n14419 out.n14418 0.007
R83129 out.n14588 out.n14587 0.007
R83130 out.n13245 out.n12854 0.007
R83131 out.n11975 out.n11560 0.007
R83132 out.n11975 out.n11561 0.007
R83133 out.n5043 out.n5040 0.007
R83134 out.n5023 out.n5022 0.007
R83135 out.n5120 out.n5119 0.007
R83136 out.n5129 out.n5126 0.007
R83137 out.n5003 out.n5002 0.007
R83138 out.n1010 out.n1009 0.007
R83139 out.n1026 out.n1021 0.007
R83140 out.n1032 out.n1030 0.007
R83141 out.n1043 out.n1042 0.007
R83142 out.n5093 out.n5092 0.007
R83143 out.n942 out.n939 0.007
R83144 out.n943 out.n942 0.007
R83145 out.n1098 out.n1097 0.007
R83146 out.n959 out.n958 0.007
R83147 out.n2745 out.n2744 0.007
R83148 out.n5851 out.n5850 0.007
R83149 out.n5802 out.n5800 0.007
R83150 out.n5777 out.n5774 0.007
R83151 out.n5728 out.n5727 0.007
R83152 out.n5677 out.n5676 0.007
R83153 out.n2866 out.n2865 0.007
R83154 out.n2830 out.n2829 0.007
R83155 out.n2753 out.n2752 0.007
R83156 out.n1446 out.n1445 0.007
R83157 out.n1450 out.n1449 0.007
R83158 out.n5423 out.n5422 0.007
R83159 out.n5524 out.n5521 0.007
R83160 out.n5575 out.n5574 0.007
R83161 out.n1357 out.n1355 0.007
R83162 out.n1530 out.n1529 0.007
R83163 out.n1153 out.n1152 0.007
R83164 out.n5318 out.n5316 0.007
R83165 out.n5310 out.n5309 0.007
R83166 out.n5302 out.n5299 0.007
R83167 out.n5292 out.n5291 0.007
R83168 out.n5274 out.n5271 0.007
R83169 out.n5225 out.n5224 0.007
R83170 out.n1244 out.n1243 0.007
R83171 out.n1239 out.n1237 0.007
R83172 out.n1224 out.n1223 0.007
R83173 out.n5177 out.n5174 0.007
R83174 out.n1163 out.n1160 0.007
R83175 out.n1160 out.n1159 0.007
R83176 out.n1284 out.n1282 0.007
R83177 out.n6565 out.n6561 0.007
R83178 out.n6504 out.n6502 0.007
R83179 out.n6609 out.n6608 0.007
R83180 out.n6468 out.n6465 0.007
R83181 out.n6729 out.n6728 0.007
R83182 out.n2091 out.n2089 0.007
R83183 out.n2168 out.n2167 0.007
R83184 out.n1874 out.n1873 0.007
R83185 out.n6423 out.n6422 0.007
R83186 out.n6374 out.n6372 0.007
R83187 out.n6218 out.n6215 0.007
R83188 out.n6305 out.n6304 0.007
R83189 out.n6254 out.n6253 0.007
R83190 out.n1990 out.n1989 0.007
R83191 out.n1954 out.n1953 0.007
R83192 out.n1882 out.n1881 0.007
R83193 out.n5886 out.n5883 0.007
R83194 out.n6118 out.n6116 0.007
R83195 out.n6109 out.n6108 0.007
R83196 out.n5893 out.n5890 0.007
R83197 out.n6032 out.n6031 0.007
R83198 out.n5914 out.n5911 0.007
R83199 out.n5921 out.n5920 0.007
R83200 out.n5920 out.n5917 0.007
R83201 out.n5929 out.n5928 0.007
R83202 out.n5984 out.n5983 0.007
R83203 out.n6167 out.n6166 0.007
R83204 out.n1547 out.n1546 0.007
R83205 out.n5943 out.n5942 0.007
R83206 out.n1649 out.n1648 0.007
R83207 out.n6985 out.n6984 0.007
R83208 out.n6936 out.n6934 0.007
R83209 out.n6911 out.n6908 0.007
R83210 out.n6862 out.n6861 0.007
R83211 out.n6811 out.n6810 0.007
R83212 out.n1770 out.n1769 0.007
R83213 out.n1734 out.n1733 0.007
R83214 out.n1657 out.n1656 0.007
R83215 out.n2290 out.n2289 0.007
R83216 out.n2294 out.n2293 0.007
R83217 out.n7284 out.n7283 0.007
R83218 out.n7382 out.n7379 0.007
R83219 out.n7433 out.n7432 0.007
R83220 out.n2201 out.n2199 0.007
R83221 out.n2377 out.n2376 0.007
R83222 out.n2404 out.n2402 0.007
R83223 out.n7240 out.n7237 0.007
R83224 out.n7192 out.n7191 0.007
R83225 out.n7039 out.n7036 0.007
R83226 out.n7163 out.n7162 0.007
R83227 out.n7045 out.n7042 0.007
R83228 out.n2505 out.n2504 0.007
R83229 out.n2508 out.n2505 0.007
R83230 out.n2499 out.n2498 0.007
R83231 out.n7091 out.n7090 0.007
R83232 out.n2419 out.n2416 0.007
R83233 out.n2410 out.n2409 0.007
R83234 out.n2428 out.n2427 0.007
R83235 out.n2436 out.n2435 0.007
R83236 out.n2438 out.n2437 0.007
R83237 out.n2442 out.n2441 0.007
R83238 out.n7757 out.n7755 0.007
R83239 out.n7491 out.n7488 0.007
R83240 out.n7518 out.n7517 0.007
R83241 out.n7658 out.n7657 0.007
R83242 out.n7542 out.n7540 0.007
R83243 out.n7569 out.n7568 0.007
R83244 out.n2631 out.n2630 0.007
R83245 out.n7472 out.n7471 0.007
R83246 out.n2620 out.n2619 0.007
R83247 out.n7466 out.n7465 0.007
R83248 out.n7467 out.n7466 0.007
R83249 out.n2599 out.n2598 0.007
R83250 out.n7011 out.n7010 0.007
R83251 out.n6202 out.n6201 0.007
R83252 out.n3099 out.n3098 0.007
R83253 out.n6196 out.n6195 0.007
R83254 out.n5610 out.n5609 0.007
R83255 out.n5864 out.n5863 0.007
R83256 out.n7477 out.n7476 0.007
R83257 out.n10708 out.n10292 0.007
R83258 out.n10708 out.n10294 0.007
R83259 out.n16269 out.n16268 0.007
R83260 out.n14569 out.n14568 0.007
R83261 out.n14570 out.n14569 0.007
R83262 out.n14607 out.n14606 0.007
R83263 out.n14678 out.n14677 0.007
R83264 out.n14749 out.n14748 0.007
R83265 out.n14820 out.n14819 0.007
R83266 out.n14891 out.n14890 0.007
R83267 out.n14962 out.n14961 0.007
R83268 out.n8891 out.n8890 0.007
R83269 out.n8892 out.n8891 0.007
R83270 out.n8896 out.n8895 0.007
R83271 out.n8897 out.n8896 0.007
R83272 out.n8933 out.n8932 0.007
R83273 out.n8934 out.n8933 0.007
R83274 out.n8968 out.n8967 0.007
R83275 out.n8969 out.n8968 0.007
R83276 out.n8973 out.n8972 0.007
R83277 out.n8974 out.n8973 0.007
R83278 out.n8978 out.n8977 0.007
R83279 out.n8979 out.n8978 0.007
R83280 out.n17304 out.n17303 0.007
R83281 out.n17303 out.n17302 0.007
R83282 out.n17299 out.n17298 0.007
R83283 out.n17298 out.n17297 0.007
R83284 out.n17294 out.n17293 0.007
R83285 out.n17293 out.n17292 0.007
R83286 out.n16050 out.n16049 0.007
R83287 out.n16046 out.n16045 0.007
R83288 out.n16045 out.n16044 0.007
R83289 out.n16041 out.n16040 0.007
R83290 out.n16040 out.n16039 0.007
R83291 out.n16036 out.n16035 0.007
R83292 out.n16035 out.n16034 0.007
R83293 out.n16031 out.n16030 0.007
R83294 out.n16030 out.n16029 0.007
R83295 out.n15688 out.n15687 0.007
R83296 out.n15616 out.n15615 0.007
R83297 out.n15612 out.n15611 0.007
R83298 out.n15611 out.n15610 0.007
R83299 out.n15468 out.n15467 0.007
R83300 out.n8917 out.n8916 0.007
R83301 out.n16076 out.n16075 0.007
R83302 out.n8955 out.n8954 0.007
R83303 out.n3135 out.n3134 0.006
R83304 out.n3020 out.n3019 0.006
R83305 out.n9 out.n7 0.006
R83306 out.n3236 out.n3235 0.006
R83307 out.n3258 out.n3257 0.006
R83308 out.n3205 out.n3204 0.006
R83309 out.n10707 out.n10682 0.006
R83310 out.n11974 out.n11949 0.006
R83311 out.n4835 out.n4808 0.006
R83312 out.n4835 out.n4826 0.006
R83313 out.n2955 out.n2954 0.006
R83314 out.n12394 out.n11977 0.006
R83315 out.n10264 out.n10263 0.006
R83316 out.n10161 out.n10160 0.006
R83317 out.n12957 out.n12956 0.006
R83318 out.n12092 out.n12091 0.006
R83319 out.n11269 out.n11268 0.006
R83320 out.n10839 out.n10838 0.006
R83321 out.n11672 out.n11671 0.006
R83322 out.n10405 out.n10404 0.006
R83323 out.n15563 out.n15385 0.006
R83324 out.n14587 out.n14586 0.006
R83325 out.n15159 out.n15158 0.006
R83326 out.n16235 out.n16203 0.006
R83327 out.n15938 out.n15906 0.006
R83328 out.n15643 out.n15565 0.006
R83329 out.n8929 out.n8918 0.006
R83330 out.n12823 out.n12404 0.006
R83331 out.n12393 out.n11978 0.006
R83332 out.n13670 out.n13643 0.006
R83333 out.n11555 out.n11540 0.006
R83334 out.n11132 out.n11113 0.006
R83335 out.n13703 out.n13676 0.006
R83336 out.n14149 out.n14148 0.006
R83337 out.n1077 out.n1075 0.006
R83338 out.n5819 out.n5818 0.006
R83339 out.n5353 out.n5352 0.006
R83340 out.n6391 out.n6390 0.006
R83341 out.n6054 out.n6053 0.006
R83342 out.n6953 out.n6952 0.006
R83343 out.n7774 out.n7773 0.006
R83344 out.n2603 out.n2602 0.006
R83345 out.n3133 out.n3130 0.006
R83346 out.n3016 out.n3015 0.006
R83347 out.n3253 out.n3252 0.006
R83348 out.n3005 out.n3004 0.006
R83349 out.n2598 out.n2597 0.006
R83350 out.n7010 out.n7009 0.006
R83351 out.n1632 out.n1631 0.006
R83352 out.n1631 out.n1630 0.006
R83353 out.n3098 out.n3097 0.006
R83354 out.n1851 out.n1850 0.006
R83355 out.n1619 out.n1618 0.006
R83356 out.n6446 out.n6445 0.006
R83357 out.n6447 out.n6446 0.006
R83358 out.n6448 out.n6447 0.006
R83359 out.n2178 out.n2177 0.006
R83360 out.n2177 out.n2176 0.006
R83361 out.n5607 out.n5606 0.006
R83362 out.n5863 out.n5862 0.006
R83363 out.n3009 out.n3008 0.006
R83364 out.n2613 out.n2612 0.006
R83365 out.n2612 out.n2611 0.006
R83366 out.n2729 out.n2728 0.006
R83367 out.n35 out.n34 0.006
R83368 out.n14600 out.n14599 0.006
R83369 out.n14670 out.n14637 0.006
R83370 out.n14671 out.n14670 0.006
R83371 out.n14741 out.n14708 0.006
R83372 out.n14742 out.n14741 0.006
R83373 out.n14812 out.n14779 0.006
R83374 out.n14813 out.n14812 0.006
R83375 out.n14883 out.n14850 0.006
R83376 out.n14884 out.n14883 0.006
R83377 out.n14954 out.n14921 0.006
R83378 out.n14955 out.n14954 0.006
R83379 out.n15022 out.n14992 0.006
R83380 out.n15023 out.n15022 0.006
R83381 out.n15087 out.n15057 0.006
R83382 out.n15088 out.n15087 0.006
R83383 out.n15200 out.n15199 0.006
R83384 out.n15264 out.n15232 0.006
R83385 out.n15265 out.n15264 0.006
R83386 out.n15329 out.n15297 0.006
R83387 out.n15330 out.n15329 0.006
R83388 out.n15363 out.n15362 0.006
R83389 out.n16236 out.n16235 0.006
R83390 out.n16199 out.n16171 0.006
R83391 out.n16139 out.n16138 0.006
R83392 out.n16138 out.n16110 0.006
R83393 out.n16078 out.n16077 0.006
R83394 out.n15902 out.n15874 0.006
R83395 out.n15842 out.n15841 0.006
R83396 out.n15841 out.n15813 0.006
R83397 out.n15781 out.n15780 0.006
R83398 out.n15780 out.n15752 0.006
R83399 out.n15715 out.n15714 0.006
R83400 out.n15714 out.n15681 0.006
R83401 out.n15644 out.n15643 0.006
R83402 out.n15561 out.n15533 0.006
R83403 out.n15496 out.n15495 0.006
R83404 out.n15495 out.n15461 0.006
R83405 out.n15503 out.n15502 0.006
R83406 out.n15615 out.n15613 0.006
R83407 out.n15613 out.n15612 0.006
R83408 out.n15651 out.n15650 0.006
R83409 out.n15722 out.n15721 0.006
R83410 out.n16034 out.n16032 0.006
R83411 out.n16032 out.n16031 0.006
R83412 out.n16039 out.n16037 0.006
R83413 out.n16037 out.n16036 0.006
R83414 out.n16044 out.n16042 0.006
R83415 out.n16042 out.n16041 0.006
R83416 out.n16049 out.n16047 0.006
R83417 out.n16047 out.n16046 0.006
R83418 out.n17292 out.n17290 0.006
R83419 out.n17290 out.n17289 0.006
R83420 out.n17297 out.n17295 0.006
R83421 out.n17295 out.n17294 0.006
R83422 out.n17302 out.n17300 0.006
R83423 out.n17300 out.n17299 0.006
R83424 out.n17305 out.n17304 0.006
R83425 out.n8980 out.n8979 0.006
R83426 out.n8975 out.n8974 0.006
R83427 out.n8977 out.n8975 0.006
R83428 out.n8970 out.n8969 0.006
R83429 out.n8972 out.n8970 0.006
R83430 out.n8965 out.n8934 0.006
R83431 out.n8967 out.n8965 0.006
R83432 out.n8930 out.n8897 0.006
R83433 out.n8932 out.n8930 0.006
R83434 out.n8893 out.n8892 0.006
R83435 out.n8895 out.n8893 0.006
R83436 out.n8888 out.n8887 0.006
R83437 out.n8890 out.n8888 0.006
R83438 out.n14928 out.n14927 0.006
R83439 out.n14857 out.n14856 0.006
R83440 out.n14786 out.n14785 0.006
R83441 out.n14715 out.n14714 0.006
R83442 out.n14644 out.n14643 0.006
R83443 out.n14571 out.n14570 0.006
R83444 out.n14568 out.n14566 0.006
R83445 out.n48 out.n47 0.006
R83446 out.n4835 out.n4831 0.006
R83447 out.n17185 out.n17151 0.006
R83448 out.n1535 out.n1534 0.006
R83449 out.n2182 out.n2181 0.006
R83450 out.n6437 out.n6436 0.006
R83451 out.n2961 out.n934 0.006
R83452 out.n1624 out.n1623 0.006
R83453 out.n12824 out.n12403 0.006
R83454 out.n17265 out.n17262 0.006
R83455 out.n5861 out.n5860 0.006
R83456 out.n7797 out.n7795 0.005
R83457 out.n10283 out.n10271 0.005
R83458 out.n15937 out.n15936 0.005
R83459 out.n13 out.n12 0.005
R83460 out.n15461 out.n15459 0.005
R83461 out.n15533 out.n15531 0.005
R83462 out.n15531 out.n15496 0.005
R83463 out.n15681 out.n15679 0.005
R83464 out.n15679 out.n15644 0.005
R83465 out.n15752 out.n15750 0.005
R83466 out.n15750 out.n15715 0.005
R83467 out.n15813 out.n15811 0.005
R83468 out.n15811 out.n15781 0.005
R83469 out.n15874 out.n15872 0.005
R83470 out.n15872 out.n15842 0.005
R83471 out.n16110 out.n16108 0.005
R83472 out.n16108 out.n16078 0.005
R83473 out.n16171 out.n16169 0.005
R83474 out.n16169 out.n16139 0.005
R83475 out.n16266 out.n16236 0.005
R83476 out.n15360 out.n15330 0.005
R83477 out.n15362 out.n15360 0.005
R83478 out.n15295 out.n15265 0.005
R83479 out.n15297 out.n15295 0.005
R83480 out.n15230 out.n15200 0.005
R83481 out.n15232 out.n15230 0.005
R83482 out.n15120 out.n15088 0.005
R83483 out.n15055 out.n15023 0.005
R83484 out.n15057 out.n15055 0.005
R83485 out.n14990 out.n14955 0.005
R83486 out.n14992 out.n14990 0.005
R83487 out.n14919 out.n14884 0.005
R83488 out.n14921 out.n14919 0.005
R83489 out.n14848 out.n14813 0.005
R83490 out.n14850 out.n14848 0.005
R83491 out.n14777 out.n14742 0.005
R83492 out.n14779 out.n14777 0.005
R83493 out.n14706 out.n14671 0.005
R83494 out.n14708 out.n14706 0.005
R83495 out.n14635 out.n14600 0.005
R83496 out.n14637 out.n14635 0.005
R83497 out.n15158 out.n15126 0.005
R83498 out.n15939 out.n15938 0.005
R83499 out.n4835 out.n4815 0.005
R83500 out.n6746 out.n6744 0.005
R83501 out.n6182 out.n6180 0.005
R83502 out.n7884 out.n7883 0.005
R83503 out.n7961 out.n7960 0.005
R83504 out.n8038 out.n8037 0.005
R83505 out.n8115 out.n8114 0.005
R83506 out.n8192 out.n8191 0.005
R83507 out.n8269 out.n8268 0.005
R83508 out.n8346 out.n8345 0.005
R83509 out.n8423 out.n8422 0.005
R83510 out.n8500 out.n8499 0.005
R83511 out.n8577 out.n8576 0.005
R83512 out.n8654 out.n8653 0.005
R83513 out.n8731 out.n8730 0.005
R83514 out.n910 out.n909 0.005
R83515 out.n3907 out.n3906 0.005
R83516 out.n3830 out.n3829 0.005
R83517 out.n3753 out.n3752 0.005
R83518 out.n3676 out.n3675 0.005
R83519 out.n3599 out.n3598 0.005
R83520 out.n3522 out.n3521 0.005
R83521 out.n3445 out.n3444 0.005
R83522 out.n3368 out.n3367 0.005
R83523 out.n3291 out.n3290 0.005
R83524 out.n3118 out.n3115 0.005
R83525 out.n3118 out.n3117 0.005
R83526 out.n2994 out.n2993 0.005
R83527 out.n2610 out.n2609 0.005
R83528 out.n1629 out.n1628 0.005
R83529 out.n6759 out.n6758 0.005
R83530 out.n5604 out.n5603 0.005
R83531 out.n14432 out.n14343 0.005
R83532 out.n5106 out.n5030 0.005
R83533 out.n9447 out.n9446 0.005
R83534 out.n5592 out.n5590 0.005
R83535 out.n7450 out.n7448 0.005
R83536 out.n10288 out.n10287 0.005
R83537 out.n15642 out.n15641 0.005
R83538 out.n3135 out.n3133 0.005
R83539 out.n14562 out.n14180 0.005
R83540 out.n14557 out.n14555 0.005
R83541 out.n15966 out.n15963 0.005
R83542 out.n16201 out.n15368 0.005
R83543 out.n8920 out.n8919 0.005
R83544 out.n15161 out.n15160 0.005
R83545 out.n16269 out.n15363 0.005
R83546 out.n16202 out.n16201 0.005
R83547 out.n15905 out.n15904 0.005
R83548 out.n15564 out.n15563 0.005
R83549 out.n8929 out.n8920 0.005
R83550 out.n15187 out.n15186 0.005
R83551 out.n15978 out.n15966 0.005
R83552 out.n16002 out.n16001 0.005
R83553 out.n15605 out.n15593 0.005
R83554 out.n17142 out.n17141 0.005
R83555 out.n17075 out.n17074 0.005
R83556 out.n17009 out.n17008 0.005
R83557 out.n16943 out.n16942 0.005
R83558 out.n16877 out.n16876 0.005
R83559 out.n16811 out.n16810 0.005
R83560 out.n16745 out.n16744 0.005
R83561 out.n16679 out.n16678 0.005
R83562 out.n16613 out.n16612 0.005
R83563 out.n16547 out.n16546 0.005
R83564 out.n16483 out.n16482 0.005
R83565 out.n16417 out.n16416 0.005
R83566 out.n16349 out.n16348 0.005
R83567 out.n9994 out.n9993 0.005
R83568 out.n9958 out.n9957 0.005
R83569 out.n9890 out.n9889 0.005
R83570 out.n9851 out.n9850 0.005
R83571 out.n9815 out.n9814 0.005
R83572 out.n9779 out.n9778 0.005
R83573 out.n9743 out.n9742 0.005
R83574 out.n9707 out.n9706 0.005
R83575 out.n9651 out.n9650 0.005
R83576 out.n9612 out.n9611 0.005
R83577 out.n9576 out.n9575 0.005
R83578 out.n9540 out.n9539 0.005
R83579 out.n9423 out.n9422 0.005
R83580 out.n5688 out.n5687 0.005
R83581 out.n3028 out.n3026 0.005
R83582 out.n5236 out.n5235 0.005
R83583 out.n6265 out.n6264 0.005
R83584 out.n1855 out.n1854 0.005
R83585 out.n4800 out.n4786 0.005
R83586 out.n4763 out.n4751 0.005
R83587 out.n4737 out.n4724 0.005
R83588 out.n4699 out.n4687 0.005
R83589 out.n4673 out.n4660 0.005
R83590 out.n4637 out.n4625 0.005
R83591 out.n4609 out.n4595 0.005
R83592 out.n4541 out.n4528 0.005
R83593 out.n4506 out.n4492 0.005
R83594 out.n4478 out.n4466 0.005
R83595 out.n4441 out.n4429 0.005
R83596 out.n4414 out.n4401 0.005
R83597 out.n4313 out.n4297 0.005
R83598 out.n4282 out.n4271 0.005
R83599 out.n4247 out.n4235 0.005
R83600 out.n4219 out.n4206 0.005
R83601 out.n4183 out.n4172 0.005
R83602 out.n4155 out.n4140 0.005
R83603 out.n4120 out.n4109 0.005
R83604 out.n4092 out.n4079 0.005
R83605 out.n4054 out.n4042 0.005
R83606 out.n4026 out.n4013 0.005
R83607 out.n919 out.n890 0.005
R83608 out.n858 out.n843 0.005
R83609 out.n768 out.n751 0.005
R83610 out.n729 out.n720 0.005
R83611 out.n705 out.n691 0.005
R83612 out.n664 out.n652 0.005
R83613 out.n638 out.n625 0.005
R83614 out.n511 out.n497 0.005
R83615 out.n472 out.n458 0.005
R83616 out.n444 out.n432 0.005
R83617 out.n409 out.n396 0.005
R83618 out.n381 out.n369 0.005
R83619 out.n344 out.n330 0.005
R83620 out.n313 out.n300 0.005
R83621 out.n274 out.n263 0.005
R83622 out.n251 out.n239 0.005
R83623 out.n213 out.n200 0.005
R83624 out.n185 out.n172 0.005
R83625 out.n148 out.n135 0.005
R83626 out.n119 out.n108 0.005
R83627 out.n88 out.n74 0.005
R83628 out.n6822 out.n6821 0.005
R83629 out.n3004 out.n3001 0.005
R83630 out.n7203 out.n7202 0.005
R83631 out.n7669 out.n7668 0.005
R83632 out.n2619 out.n2618 0.005
R83633 out.n7465 out.n7464 0.005
R83634 out.n3252 out.n3247 0.005
R83635 out.n2983 out.n2982 0.005
R83636 out.n1850 out.n1849 0.005
R83637 out.n1618 out.n1617 0.005
R83638 out.n5862 out.n5861 0.005
R83639 out.n2728 out.n2727 0.005
R83640 out.n4506 out.n4481 0.005
R83641 out.n4441 out.n4417 0.005
R83642 out.n4313 out.n4285 0.005
R83643 out.n4247 out.n4222 0.005
R83644 out.n4183 out.n4158 0.005
R83645 out.n4120 out.n4095 0.005
R83646 out.n4054 out.n4029 0.005
R83647 out.n919 out.n918 0.005
R83648 out.n858 out.n831 0.005
R83649 out.n344 out.n316 0.005
R83650 out.n213 out.n188 0.005
R83651 out.n148 out.n122 0.005
R83652 out.n88 out.n59 0.005
R83653 out.n16234 out.n16233 0.005
R83654 out.n13105 out.n13103 0.005
R83655 out.n11820 out.n11818 0.005
R83656 out.n10553 out.n10551 0.005
R83657 out.n5620 out.n5618 0.005
R83658 out.n7015 out.n7013 0.005
R83659 out.n2954 out.n2953 0.005
R83660 out.n8954 out.n8953 0.005
R83661 out.n3054 out.n3053 0.005
R83662 out.n3115 out.n3113 0.005
R83663 out.n3329 out.n3328 0.005
R83664 out.n3406 out.n3405 0.005
R83665 out.n3483 out.n3482 0.005
R83666 out.n3560 out.n3559 0.005
R83667 out.n3637 out.n3636 0.005
R83668 out.n3714 out.n3713 0.005
R83669 out.n3791 out.n3790 0.005
R83670 out.n3868 out.n3867 0.005
R83671 out.n3945 out.n3944 0.005
R83672 out.n8774 out.n8769 0.005
R83673 out.n8691 out.n8688 0.005
R83674 out.n8614 out.n8611 0.005
R83675 out.n8537 out.n8534 0.005
R83676 out.n8460 out.n8457 0.005
R83677 out.n8383 out.n8380 0.005
R83678 out.n8306 out.n8303 0.005
R83679 out.n8229 out.n8226 0.005
R83680 out.n8152 out.n8149 0.005
R83681 out.n8075 out.n8072 0.005
R83682 out.n7998 out.n7995 0.005
R83683 out.n7921 out.n7918 0.005
R83684 out.n7844 out.n7841 0.005
R83685 out.n5170 out.n5169 0.005
R83686 out.n12240 out.n12238 0.005
R83687 out.n13593 out.n13592 0.005
R83688 out.n14048 out.n14047 0.005
R83689 out.n2975 out.n2974 0.005
R83690 out.n3011 out.n3010 0.005
R83691 out.n7462 out.n7461 0.005
R83692 out.n17185 out.n17153 0.005
R83693 out.n2956 out.n2955 0.005
R83694 out.n9506 out.n9491 0.005
R83695 out.n17185 out.n17157 0.005
R83696 out.n6761 out.n6760 0.005
R83697 out.n14599 out.n14110 0.005
R83698 out.n17185 out.n17161 0.005
R83699 out.n5859 out.n5858 0.005
R83700 out.n3206 out.n3205 0.005
R83701 out.n3259 out.n3258 0.005
R83702 out.n10987 out.n10985 0.005
R83703 out.n12759 out.n12758 0.004
R83704 out.n11414 out.n11412 0.004
R83705 out.n17184 out.n17182 0.004
R83706 out.n17136 out.n17135 0.004
R83707 out.n17070 out.n17069 0.004
R83708 out.n17004 out.n17003 0.004
R83709 out.n16938 out.n16937 0.004
R83710 out.n16872 out.n16871 0.004
R83711 out.n16806 out.n16805 0.004
R83712 out.n16740 out.n16739 0.004
R83713 out.n16674 out.n16673 0.004
R83714 out.n16608 out.n16607 0.004
R83715 out.n16542 out.n16541 0.004
R83716 out.n16478 out.n16477 0.004
R83717 out.n16412 out.n16411 0.004
R83718 out.n16344 out.n16343 0.004
R83719 out.n9989 out.n9988 0.004
R83720 out.n9953 out.n9952 0.004
R83721 out.n9885 out.n9884 0.004
R83722 out.n9846 out.n9845 0.004
R83723 out.n9810 out.n9809 0.004
R83724 out.n9774 out.n9773 0.004
R83725 out.n9738 out.n9737 0.004
R83726 out.n9702 out.n9701 0.004
R83727 out.n9646 out.n9645 0.004
R83728 out.n9607 out.n9606 0.004
R83729 out.n9571 out.n9570 0.004
R83730 out.n9535 out.n9534 0.004
R83731 out.n9401 out.n9399 0.004
R83732 out.n505 out.n503 0.004
R83733 out.n525 out.n524 0.004
R83734 out.n566 out.n565 0.004
R83735 out.n760 out.n758 0.004
R83736 out.n784 out.n783 0.004
R83737 out.n4928 out.n4927 0.004
R83738 out.n4303 out.n4302 0.004
R83739 out.n4344 out.n4342 0.004
R83740 out.n4536 out.n4535 0.004
R83741 out.n4794 out.n4792 0.004
R83742 out.n915 out.n914 0.004
R83743 out.n873 out.n872 0.004
R83744 out.n4777 out.n4776 0.004
R83745 out.n4714 out.n4713 0.004
R83746 out.n4649 out.n4648 0.004
R83747 out.n4584 out.n4583 0.004
R83748 out.n4519 out.n4518 0.004
R83749 out.n4327 out.n4326 0.004
R83750 out.n742 out.n741 0.004
R83751 out.n680 out.n679 0.004
R83752 out.n615 out.n614 0.004
R83753 out.n550 out.n549 0.004
R83754 out.n488 out.n487 0.004
R83755 out.n422 out.n421 0.004
R83756 out.n358 out.n357 0.004
R83757 out.n228 out.n227 0.004
R83758 out.n2063 out.n2061 0.004
R83759 out.n2934 out.n2932 0.004
R83760 out.n1838 out.n1836 0.004
R83761 out.n2586 out.n2584 0.004
R83762 out.n15426 out.n15408 0.004
R83763 out.n3176 out.n3175 0.004
R83764 out.n3097 out.n3096 0.004
R83765 out.n3109 out.n3106 0.004
R83766 out.n5612 out.n5170 0.004
R83767 out.n15390 out.n15389 0.004
R83768 out.n10265 out.n10264 0.004
R83769 out.n10160 out.n10159 0.004
R83770 out.n10276 out.n10275 0.004
R83771 out.n15160 out.n15159 0.004
R83772 out.n15906 out.n15905 0.004
R83773 out.n17185 out.n17177 0.004
R83774 out.n17142 out.n17129 0.004
R83775 out.n17110 out.n17101 0.004
R83776 out.n17075 out.n17063 0.004
R83777 out.n17044 out.n17035 0.004
R83778 out.n17009 out.n16997 0.004
R83779 out.n16980 out.n16971 0.004
R83780 out.n16943 out.n16931 0.004
R83781 out.n16912 out.n16903 0.004
R83782 out.n16877 out.n16865 0.004
R83783 out.n16848 out.n16839 0.004
R83784 out.n16811 out.n16799 0.004
R83785 out.n16782 out.n16773 0.004
R83786 out.n16745 out.n16733 0.004
R83787 out.n16714 out.n16705 0.004
R83788 out.n16679 out.n16667 0.004
R83789 out.n16648 out.n16639 0.004
R83790 out.n16613 out.n16601 0.004
R83791 out.n16584 out.n16575 0.004
R83792 out.n16547 out.n16535 0.004
R83793 out.n16516 out.n16507 0.004
R83794 out.n16483 out.n16471 0.004
R83795 out.n16450 out.n16441 0.004
R83796 out.n16417 out.n16405 0.004
R83797 out.n16384 out.n16375 0.004
R83798 out.n16349 out.n16337 0.004
R83799 out.n16318 out.n16309 0.004
R83800 out.n9052 out.n9045 0.004
R83801 out.n9994 out.n9982 0.004
R83802 out.n9084 out.n9075 0.004
R83803 out.n9958 out.n9946 0.004
R83804 out.n9922 out.n9913 0.004
R83805 out.n9890 out.n9878 0.004
R83806 out.n9119 out.n9110 0.004
R83807 out.n9851 out.n9839 0.004
R83808 out.n9153 out.n9144 0.004
R83809 out.n9815 out.n9803 0.004
R83810 out.n9187 out.n9178 0.004
R83811 out.n9779 out.n9767 0.004
R83812 out.n9221 out.n9212 0.004
R83813 out.n9743 out.n9731 0.004
R83814 out.n9255 out.n9246 0.004
R83815 out.n9707 out.n9695 0.004
R83816 out.n9289 out.n9280 0.004
R83817 out.n9651 out.n9639 0.004
R83818 out.n9322 out.n9313 0.004
R83819 out.n9612 out.n9600 0.004
R83820 out.n9356 out.n9347 0.004
R83821 out.n9576 out.n9564 0.004
R83822 out.n9390 out.n9381 0.004
R83823 out.n9540 out.n9528 0.004
R83824 out.n9423 out.n9413 0.004
R83825 out.n14147 out.n14137 0.004
R83826 out.n17277 out.n17265 0.004
R83827 out.n9506 out.n9501 0.004
R83828 out.n16285 out.n10009 0.004
R83829 out.n9506 out.n9476 0.004
R83830 out.n17186 out.n17147 0.004
R83831 out.n17188 out.n17144 0.004
R83832 out.n17190 out.n17080 0.004
R83833 out.n17192 out.n17077 0.004
R83834 out.n17194 out.n17014 0.004
R83835 out.n17196 out.n17011 0.004
R83836 out.n17198 out.n16948 0.004
R83837 out.n17200 out.n16945 0.004
R83838 out.n17202 out.n16882 0.004
R83839 out.n17204 out.n16879 0.004
R83840 out.n17206 out.n16816 0.004
R83841 out.n17208 out.n16813 0.004
R83842 out.n17210 out.n16750 0.004
R83843 out.n17212 out.n16747 0.004
R83844 out.n17214 out.n16684 0.004
R83845 out.n17216 out.n16681 0.004
R83846 out.n17218 out.n16618 0.004
R83847 out.n17220 out.n16615 0.004
R83848 out.n17222 out.n16552 0.004
R83849 out.n17224 out.n16549 0.004
R83850 out.n17226 out.n16488 0.004
R83851 out.n17228 out.n16485 0.004
R83852 out.n17230 out.n16422 0.004
R83853 out.n17232 out.n16419 0.004
R83854 out.n17234 out.n16354 0.004
R83855 out.n17236 out.n16351 0.004
R83856 out.n17238 out.n16288 0.004
R83857 out.n9999 out.n9022 0.004
R83858 out.n9997 out.n9996 0.004
R83859 out.n9963 out.n9056 0.004
R83860 out.n9961 out.n9960 0.004
R83861 out.n9925 out.n9924 0.004
R83862 out.n9891 out.n9860 0.004
R83863 out.n9856 out.n9089 0.004
R83864 out.n9854 out.n9853 0.004
R83865 out.n9820 out.n9123 0.004
R83866 out.n9818 out.n9817 0.004
R83867 out.n9784 out.n9157 0.004
R83868 out.n9782 out.n9781 0.004
R83869 out.n9748 out.n9191 0.004
R83870 out.n9746 out.n9745 0.004
R83871 out.n9712 out.n9225 0.004
R83872 out.n9710 out.n9709 0.004
R83873 out.n9676 out.n9259 0.004
R83874 out.n9674 out.n9621 0.004
R83875 out.n9617 out.n9292 0.004
R83876 out.n9615 out.n9614 0.004
R83877 out.n9581 out.n9326 0.004
R83878 out.n9579 out.n9578 0.004
R83879 out.n9545 out.n9360 0.004
R83880 out.n9543 out.n9542 0.004
R83881 out.n9509 out.n9393 0.004
R83882 out.n9506 out.n9505 0.004
R83883 out.n17310 out.n17309 0.004
R83884 out.n5620 out.n5619 0.004
R83885 out.n1290 out.n1289 0.004
R83886 out.n1335 out.n1334 0.004
R83887 out.n3235 out.n3234 0.004
R83888 out.n4699 out.n4688 0.004
R83889 out.n4637 out.n4626 0.004
R83890 out.n4570 out.n4557 0.004
R83891 out.n4441 out.n4430 0.004
R83892 out.n4378 out.n4365 0.004
R83893 out.n4247 out.n4236 0.004
R83894 out.n4183 out.n4173 0.004
R83895 out.n4120 out.n4110 0.004
R83896 out.n4054 out.n4043 0.004
R83897 out.n4942 out.n4929 0.004
R83898 out.n4942 out.n4933 0.004
R83899 out.n858 out.n844 0.004
R83900 out.n664 out.n653 0.004
R83901 out.n601 out.n587 0.004
R83902 out.n472 out.n459 0.004
R83903 out.n409 out.n397 0.004
R83904 out.n344 out.n331 0.004
R83905 out.n213 out.n201 0.004
R83906 out.n88 out.n75 0.004
R83907 out.n56 out.n49 0.004
R83908 out.n7015 out.n7014 0.004
R83909 out.n4737 out.n4721 0.004
R83910 out.n4699 out.n4684 0.004
R83911 out.n4673 out.n4657 0.004
R83912 out.n4637 out.n4622 0.004
R83913 out.n4609 out.n4592 0.004
R83914 out.n4570 out.n4554 0.004
R83915 out.n4441 out.n4426 0.004
R83916 out.n4414 out.n4398 0.004
R83917 out.n4378 out.n4362 0.004
R83918 out.n4247 out.n4232 0.004
R83919 out.n4219 out.n4203 0.004
R83920 out.n4183 out.n4169 0.004
R83921 out.n4155 out.n4137 0.004
R83922 out.n4120 out.n4106 0.004
R83923 out.n4092 out.n4076 0.004
R83924 out.n4054 out.n4039 0.004
R83925 out.n4026 out.n4010 0.004
R83926 out.n4942 out.n4924 0.004
R83927 out.n858 out.n840 0.004
R83928 out.n705 out.n688 0.004
R83929 out.n664 out.n649 0.004
R83930 out.n638 out.n622 0.004
R83931 out.n601 out.n584 0.004
R83932 out.n472 out.n455 0.004
R83933 out.n444 out.n429 0.004
R83934 out.n409 out.n393 0.004
R83935 out.n381 out.n366 0.004
R83936 out.n344 out.n327 0.004
R83937 out.n313 out.n297 0.004
R83938 out.n251 out.n234 0.004
R83939 out.n213 out.n197 0.004
R83940 out.n185 out.n169 0.004
R83941 out.n148 out.n132 0.004
R83942 out.n119 out.n105 0.004
R83943 out.n88 out.n69 0.004
R83944 out.n56 out.n37 0.004
R83945 out.n7087 out.n7084 0.004
R83946 out.n2717 out.n2716 0.004
R83947 out.n7465 out.n7248 0.004
R83948 out.n2597 out.n2596 0.004
R83949 out.n3222 out.n3215 0.004
R83950 out.n7009 out.n7008 0.004
R83951 out.n6446 out.n6437 0.004
R83952 out.n3222 out.n3221 0.004
R83953 out.n911 out.n910 0.004
R83954 out.n2959 out.n2958 0.004
R83955 out.n5606 out.n5605 0.004
R83956 out.n7823 out.n7821 0.004
R83957 out.n7862 out.n7860 0.004
R83958 out.n7900 out.n7898 0.004
R83959 out.n7939 out.n7937 0.004
R83960 out.n7977 out.n7975 0.004
R83961 out.n8016 out.n8014 0.004
R83962 out.n8054 out.n8052 0.004
R83963 out.n8093 out.n8091 0.004
R83964 out.n8131 out.n8129 0.004
R83965 out.n8170 out.n8168 0.004
R83966 out.n8208 out.n8206 0.004
R83967 out.n8247 out.n8245 0.004
R83968 out.n8285 out.n8283 0.004
R83969 out.n8324 out.n8322 0.004
R83970 out.n8362 out.n8360 0.004
R83971 out.n8401 out.n8399 0.004
R83972 out.n8439 out.n8437 0.004
R83973 out.n8478 out.n8476 0.004
R83974 out.n8516 out.n8514 0.004
R83975 out.n8555 out.n8553 0.004
R83976 out.n8593 out.n8591 0.004
R83977 out.n8632 out.n8630 0.004
R83978 out.n8670 out.n8668 0.004
R83979 out.n8709 out.n8707 0.004
R83980 out.n8747 out.n8745 0.004
R83981 out.n8794 out.n8793 0.004
R83982 out.n3988 out.n3985 0.004
R83983 out.n3987 out.n3986 0.004
R83984 out.n3965 out.n3962 0.004
R83985 out.n3964 out.n3963 0.004
R83986 out.n3927 out.n3924 0.004
R83987 out.n3926 out.n3925 0.004
R83988 out.n3888 out.n3885 0.004
R83989 out.n3887 out.n3886 0.004
R83990 out.n3850 out.n3847 0.004
R83991 out.n3849 out.n3848 0.004
R83992 out.n3811 out.n3808 0.004
R83993 out.n3810 out.n3809 0.004
R83994 out.n3773 out.n3770 0.004
R83995 out.n3772 out.n3771 0.004
R83996 out.n3734 out.n3731 0.004
R83997 out.n3733 out.n3732 0.004
R83998 out.n3696 out.n3693 0.004
R83999 out.n3695 out.n3694 0.004
R84000 out.n3657 out.n3654 0.004
R84001 out.n3656 out.n3655 0.004
R84002 out.n3619 out.n3616 0.004
R84003 out.n3618 out.n3617 0.004
R84004 out.n3580 out.n3577 0.004
R84005 out.n3579 out.n3578 0.004
R84006 out.n3542 out.n3539 0.004
R84007 out.n3541 out.n3540 0.004
R84008 out.n3503 out.n3500 0.004
R84009 out.n3502 out.n3501 0.004
R84010 out.n3465 out.n3462 0.004
R84011 out.n3464 out.n3463 0.004
R84012 out.n3426 out.n3423 0.004
R84013 out.n3425 out.n3424 0.004
R84014 out.n3388 out.n3385 0.004
R84015 out.n3387 out.n3386 0.004
R84016 out.n3349 out.n3346 0.004
R84017 out.n3348 out.n3347 0.004
R84018 out.n3311 out.n3308 0.004
R84019 out.n3310 out.n3309 0.004
R84020 out.n3272 out.n3269 0.004
R84021 out.n3271 out.n3270 0.004
R84022 out.n3193 out.n3192 0.004
R84023 out.n3180 out.n3177 0.004
R84024 out.n3179 out.n3178 0.004
R84025 out.n3154 out.n3151 0.004
R84026 out.n3153 out.n3152 0.004
R84027 out.n3074 out.n3071 0.004
R84028 out.n3073 out.n3072 0.004
R84029 out.n3031 out.n3024 0.004
R84030 out.n3030 out.n3029 0.004
R84031 out.n1340 out.n1339 0.004
R84032 out.n2952 out.n2944 0.004
R84033 out.n2951 out.n2950 0.004
R84034 out.n10285 out.n10284 0.004
R84035 out.n13244 out.n13239 0.004
R84036 out.n13245 out.n13244 0.004
R84037 out.n10286 out.n10285 0.004
R84038 out.n3010 out.n3009 0.004
R84039 out.n2974 out.n2973 0.004
R84040 out.n15426 out.n15404 0.004
R84041 out.n15426 out.n15424 0.004
R84042 out.n2721 out.n2720 0.004
R84043 out.n15458 out.n15457 0.004
R84044 out.n15426 out.n15402 0.004
R84045 out.n1616 out.n1615 0.004
R84046 out.n2726 out.n2725 0.004
R84047 out.n10036 out.n10035 0.004
R84048 out.n16274 out.n16273 0.004
R84049 out.n10030 out.n10029 0.004
R84050 out.n16279 out.n16278 0.004
R84051 out.n10020 out.n10019 0.004
R84052 out.n10025 out.n10024 0.004
R84053 out.n16284 out.n16282 0.004
R84054 out.n10007 out.n10006 0.004
R84055 out.n867 out.n865 0.004
R84056 out.n881 out.n880 0.004
R84057 out.n178 out.n177 0.004
R84058 out.n306 out.n305 0.004
R84059 out.n564 out.n563 0.004
R84060 out.n757 out.n756 0.004
R84061 out.n820 out.n819 0.004
R84062 out.n4341 out.n4340 0.004
R84063 out.n4534 out.n4533 0.004
R84064 out.n4791 out.n4790 0.004
R84065 out.n528 out.n527 0.004
R84066 out.n597 out.n595 0.004
R84067 out.n787 out.n786 0.004
R84068 out.n853 out.n851 0.004
R84069 out.n4308 out.n4306 0.004
R84070 out.n4374 out.n4372 0.004
R84071 out.n4501 out.n4499 0.004
R84072 out.n4566 out.n4564 0.004
R84073 out.n4829 out.n4827 0.004
R84074 out.n4797 out.n4796 0.004
R84075 out.n4539 out.n4538 0.004
R84076 out.n4347 out.n4346 0.004
R84077 out.n887 out.n886 0.004
R84078 out.n825 out.n823 0.004
R84079 out.n765 out.n763 0.004
R84080 out.n570 out.n568 0.004
R84081 out.n310 out.n309 0.004
R84082 out.n884 out.n883 0.004
R84083 out.n4835 out.n4820 0.004
R84084 out.n4835 out.n4821 0.004
R84085 out.n7001 out.n7000 0.004
R84086 out.n5627 out.n5626 0.004
R84087 out.n15426 out.n15400 0.004
R84088 out.n15426 out.n15406 0.004
R84089 out.n49 out.n48 0.004
R84090 out.n9463 out.n9462 0.003
R84091 out.n9462 out.n9461 0.003
R84092 out.n13642 out.n13249 0.003
R84093 out.n11539 out.n11138 0.003
R84094 out.n11112 out.n10715 0.003
R84095 out.n14097 out.n13704 0.003
R84096 out.n14564 out.n14563 0.003
R84097 out.n14098 out.n14097 0.003
R84098 out.n11133 out.n11112 0.003
R84099 out.n11556 out.n11539 0.003
R84100 out.n13671 out.n13642 0.003
R84101 out.n14563 out.n14150 0.003
R84102 out.n3109 out.n3108 0.003
R84103 out.n4835 out.n4812 0.003
R84104 out.n3033 out.n3032 0.003
R84105 out.n17186 out.n4 0.003
R84106 out.n2617 out.n2616 0.003
R84107 out.n1848 out.n1847 0.003
R84108 out.n2175 out.n2174 0.003
R84109 out.n3176 out.n3173 0.003
R84110 out.n17142 out.n17128 0.003
R84111 out.n17075 out.n17062 0.003
R84112 out.n16943 out.n16930 0.003
R84113 out.n16745 out.n16732 0.003
R84114 out.n16679 out.n16666 0.003
R84115 out.n16584 out.n16574 0.003
R84116 out.n16384 out.n16374 0.003
R84117 out.n16318 out.n16308 0.003
R84118 out.n9052 out.n9042 0.003
R84119 out.n9922 out.n9912 0.003
R84120 out.n9119 out.n9109 0.003
R84121 out.n9153 out.n9143 0.003
R84122 out.n9187 out.n9177 0.003
R84123 out.n9221 out.n9211 0.003
R84124 out.n9255 out.n9245 0.003
R84125 out.n9289 out.n9279 0.003
R84126 out.n9322 out.n9312 0.003
R84127 out.n9356 out.n9346 0.003
R84128 out.n9390 out.n9380 0.003
R84129 out.n4 out.n3 0.003
R84130 out.n9440 out.n9434 0.003
R84131 out.n10282 out.n10278 0.003
R84132 out.n10227 out.n10226 0.003
R84133 out.n10226 out.n10225 0.003
R84134 out.n10216 out.n10215 0.003
R84135 out.n10215 out.n10214 0.003
R84136 out.n10153 out.n10148 0.003
R84137 out.n13101 out.n13098 0.003
R84138 out.n13092 out.n13091 0.003
R84139 out.n13155 out.n13153 0.003
R84140 out.n13198 out.n13196 0.003
R84141 out.n13190 out.n13187 0.003
R84142 out.n13203 out.n13202 0.003
R84143 out.n13003 out.n13002 0.003
R84144 out.n13074 out.n13072 0.003
R84145 out.n12960 out.n12957 0.003
R84146 out.n12803 out.n12800 0.003
R84147 out.n12429 out.n12428 0.003
R84148 out.n12425 out.n12422 0.003
R84149 out.n12673 out.n12670 0.003
R84150 out.n12711 out.n12708 0.003
R84151 out.n12775 out.n12774 0.003
R84152 out.n12764 out.n12763 0.003
R84153 out.n12565 out.n12562 0.003
R84154 out.n12558 out.n12557 0.003
R84155 out.n12577 out.n12576 0.003
R84156 out.n12597 out.n12595 0.003
R84157 out.n12816 out.n12815 0.003
R84158 out.n12466 out.n12465 0.003
R84159 out.n12530 out.n12528 0.003
R84160 out.n12236 out.n12233 0.003
R84161 out.n12227 out.n12226 0.003
R84162 out.n12290 out.n12288 0.003
R84163 out.n12333 out.n12331 0.003
R84164 out.n12325 out.n12322 0.003
R84165 out.n12338 out.n12337 0.003
R84166 out.n12138 out.n12137 0.003
R84167 out.n12209 out.n12207 0.003
R84168 out.n12095 out.n12092 0.003
R84169 out.n13637 out.n13634 0.003
R84170 out.n13273 out.n13272 0.003
R84171 out.n13506 out.n13503 0.003
R84172 out.n13545 out.n13542 0.003
R84173 out.n13609 out.n13608 0.003
R84174 out.n13598 out.n13597 0.003
R84175 out.n13398 out.n13395 0.003
R84176 out.n13391 out.n13390 0.003
R84177 out.n13410 out.n13409 0.003
R84178 out.n13430 out.n13428 0.003
R84179 out.n13655 out.n13654 0.003
R84180 out.n13661 out.n13656 0.003
R84181 out.n13363 out.n13361 0.003
R84182 out.n11410 out.n11407 0.003
R84183 out.n11401 out.n11400 0.003
R84184 out.n11459 out.n11457 0.003
R84185 out.n11502 out.n11500 0.003
R84186 out.n11494 out.n11491 0.003
R84187 out.n11507 out.n11506 0.003
R84188 out.n11312 out.n11311 0.003
R84189 out.n11383 out.n11381 0.003
R84190 out.n11272 out.n11269 0.003
R84191 out.n10983 out.n10980 0.003
R84192 out.n10974 out.n10973 0.003
R84193 out.n11032 out.n11030 0.003
R84194 out.n11075 out.n11073 0.003
R84195 out.n11067 out.n11064 0.003
R84196 out.n11080 out.n11079 0.003
R84197 out.n10885 out.n10884 0.003
R84198 out.n10956 out.n10954 0.003
R84199 out.n10842 out.n10839 0.003
R84200 out.n11816 out.n11813 0.003
R84201 out.n11807 out.n11806 0.003
R84202 out.n11870 out.n11868 0.003
R84203 out.n11913 out.n11911 0.003
R84204 out.n11905 out.n11902 0.003
R84205 out.n11918 out.n11917 0.003
R84206 out.n11718 out.n11717 0.003
R84207 out.n11789 out.n11787 0.003
R84208 out.n11675 out.n11672 0.003
R84209 out.n14092 out.n14089 0.003
R84210 out.n13728 out.n13727 0.003
R84211 out.n13961 out.n13958 0.003
R84212 out.n14000 out.n13997 0.003
R84213 out.n14064 out.n14063 0.003
R84214 out.n14053 out.n14052 0.003
R84215 out.n13853 out.n13850 0.003
R84216 out.n13846 out.n13845 0.003
R84217 out.n13865 out.n13864 0.003
R84218 out.n13885 out.n13883 0.003
R84219 out.n13688 out.n13687 0.003
R84220 out.n13694 out.n13689 0.003
R84221 out.n13818 out.n13816 0.003
R84222 out.n10549 out.n10546 0.003
R84223 out.n10540 out.n10539 0.003
R84224 out.n10603 out.n10601 0.003
R84225 out.n10646 out.n10644 0.003
R84226 out.n10638 out.n10635 0.003
R84227 out.n10651 out.n10650 0.003
R84228 out.n10451 out.n10450 0.003
R84229 out.n10522 out.n10520 0.003
R84230 out.n10408 out.n10405 0.003
R84231 out.n14515 out.n14513 0.003
R84232 out.n14232 out.n14227 0.003
R84233 out.n14208 out.n14207 0.003
R84234 out.n14223 out.n14222 0.003
R84235 out.n14548 out.n14545 0.003
R84236 out.n14341 out.n14340 0.003
R84237 out.n14351 out.n14350 0.003
R84238 out.n14464 out.n14462 0.003
R84239 out.n14288 out.n14286 0.003
R84240 out.n14303 out.n14300 0.003
R84241 out.n14293 out.n14292 0.003
R84242 out.n14418 out.n14416 0.003
R84243 out.n9507 out.n9506 0.003
R84244 out.n10713 out.n10712 0.003
R84245 out.n14119 out.n14118 0.003
R84246 out.n14569 out.n14147 0.003
R84247 out.n14114 out.n14113 0.003
R84248 out.n14598 out.n14571 0.003
R84249 out.n14604 out.n14603 0.003
R84250 out.n14634 out.n14607 0.003
R84251 out.n14641 out.n14640 0.003
R84252 out.n14669 out.n14644 0.003
R84253 out.n14675 out.n14674 0.003
R84254 out.n14705 out.n14678 0.003
R84255 out.n14712 out.n14711 0.003
R84256 out.n14740 out.n14715 0.003
R84257 out.n14746 out.n14745 0.003
R84258 out.n14776 out.n14749 0.003
R84259 out.n14783 out.n14782 0.003
R84260 out.n14811 out.n14786 0.003
R84261 out.n14817 out.n14816 0.003
R84262 out.n14847 out.n14820 0.003
R84263 out.n14854 out.n14853 0.003
R84264 out.n14882 out.n14857 0.003
R84265 out.n14888 out.n14887 0.003
R84266 out.n14918 out.n14891 0.003
R84267 out.n14925 out.n14924 0.003
R84268 out.n14953 out.n14928 0.003
R84269 out.n14959 out.n14958 0.003
R84270 out.n14989 out.n14962 0.003
R84271 out.n14996 out.n14995 0.003
R84272 out.n15027 out.n15026 0.003
R84273 out.n15061 out.n15060 0.003
R84274 out.n15092 out.n15091 0.003
R84275 out.n8901 out.n8900 0.003
R84276 out.n8930 out.n8929 0.003
R84277 out.n15130 out.n15129 0.003
R84278 out.n8938 out.n8937 0.003
R84279 out.n8965 out.n8964 0.003
R84280 out.n15170 out.n15169 0.003
R84281 out.n15204 out.n15203 0.003
R84282 out.n15236 out.n15235 0.003
R84283 out.n15269 out.n15268 0.003
R84284 out.n15301 out.n15300 0.003
R84285 out.n15334 out.n15333 0.003
R84286 out.n8987 out.n8986 0.003
R84287 out.n17309 out.n9015 0.003
R84288 out.n9019 out.n9018 0.003
R84289 out.n17241 out.n17240 0.003
R84290 out.n17244 out.n17243 0.003
R84291 out.n17300 out.n17277 0.003
R84292 out.n17246 out.n17245 0.003
R84293 out.n17280 out.n17279 0.003
R84294 out.n17282 out.n17281 0.003
R84295 out.n17285 out.n17284 0.003
R84296 out.n17287 out.n17286 0.003
R84297 out.n16073 out.n16050 0.003
R84298 out.n15945 out.n15944 0.003
R84299 out.n16047 out.n15978 0.003
R84300 out.n15947 out.n15946 0.003
R84301 out.n15981 out.n15980 0.003
R84302 out.n16042 out.n16014 0.003
R84303 out.n15983 out.n15982 0.003
R84304 out.n16017 out.n16016 0.003
R84305 out.n16019 out.n16018 0.003
R84306 out.n16022 out.n16021 0.003
R84307 out.n16024 out.n16023 0.003
R84308 out.n16027 out.n16026 0.003
R84309 out.n15747 out.n15722 0.003
R84310 out.n15719 out.n15718 0.003
R84311 out.n15711 out.n15688 0.003
R84312 out.n15685 out.n15684 0.003
R84313 out.n15676 out.n15651 0.003
R84314 out.n15648 out.n15647 0.003
R84315 out.n15639 out.n15616 0.003
R84316 out.n15572 out.n15571 0.003
R84317 out.n15613 out.n15605 0.003
R84318 out.n15574 out.n15573 0.003
R84319 out.n15608 out.n15607 0.003
R84320 out.n15528 out.n15503 0.003
R84321 out.n15500 out.n15499 0.003
R84322 out.n15492 out.n15468 0.003
R84323 out.n15465 out.n15464 0.003
R84324 out.n15455 out.n15433 0.003
R84325 out.n15398 out.n15397 0.003
R84326 out.n15430 out.n15428 0.003
R84327 out.n5028 out.n5027 0.003
R84328 out.n5040 out.n5039 0.003
R84329 out.n5138 out.n5136 0.003
R84330 out.n4974 out.n4972 0.003
R84331 out.n4990 out.n4987 0.003
R84332 out.n4979 out.n4978 0.003
R84333 out.n1013 out.n1012 0.003
R84334 out.n5092 out.n5090 0.003
R84335 out.n1075 out.n1074 0.003
R84336 out.n1127 out.n1126 0.003
R84337 out.n5632 out.n5629 0.003
R84338 out.n5769 out.n5768 0.003
R84339 out.n5752 out.n5751 0.003
R84340 out.n5647 out.n5644 0.003
R84341 out.n2869 out.n2866 0.003
R84342 out.n2859 out.n2854 0.003
R84343 out.n2860 out.n2859 0.003
R84344 out.n2852 out.n2849 0.003
R84345 out.n2839 out.n2838 0.003
R84346 out.n2845 out.n2839 0.003
R84347 out.n2835 out.n2830 0.003
R84348 out.n5691 out.n5688 0.003
R84349 out.n2762 out.n2759 0.003
R84350 out.n2781 out.n2780 0.003
R84351 out.n2790 out.n2789 0.003
R84352 out.n2797 out.n2796 0.003
R84353 out.n5508 out.n5507 0.003
R84354 out.n5498 out.n5495 0.003
R84355 out.n5574 out.n5572 0.003
R84356 out.n1337 out.n1336 0.003
R84357 out.n5336 out.n5334 0.003
R84358 out.n5262 out.n5261 0.003
R84359 out.n1210 out.n1209 0.003
R84360 out.n1201 out.n1200 0.003
R84361 out.n5239 out.n5236 0.003
R84362 out.n5363 out.n5362 0.003
R84363 out.n1282 out.n1281 0.003
R84364 out.n1286 out.n1284 0.003
R84365 out.n1292 out.n1290 0.003
R84366 out.n1333 out.n1332 0.003
R84367 out.n4838 out.n4837 0.003
R84368 out.n4841 out.n4771 0.003
R84369 out.n4844 out.n4765 0.003
R84370 out.n4847 out.n4706 0.003
R84371 out.n4850 out.n4700 0.003
R84372 out.n4673 out.n4654 0.003
R84373 out.n4853 out.n4644 0.003
R84374 out.n4856 out.n4638 0.003
R84375 out.n4609 out.n4589 0.003
R84376 out.n4859 out.n4578 0.003
R84377 out.n4570 out.n4547 0.003
R84378 out.n4861 out.n4572 0.003
R84379 out.n4864 out.n4514 0.003
R84380 out.n4867 out.n4508 0.003
R84381 out.n4870 out.n4450 0.003
R84382 out.n4872 out.n4443 0.003
R84383 out.n4875 out.n4386 0.003
R84384 out.n4878 out.n4380 0.003
R84385 out.n4881 out.n4322 0.003
R84386 out.n4883 out.n4315 0.003
R84387 out.n4886 out.n4256 0.003
R84388 out.n4888 out.n4249 0.003
R84389 out.n4890 out.n4192 0.003
R84390 out.n4893 out.n4185 0.003
R84391 out.n4896 out.n4126 0.003
R84392 out.n4120 out.n4100 0.003
R84393 out.n4899 out.n4121 0.003
R84394 out.n4092 out.n4073 0.003
R84395 out.n4902 out.n4063 0.003
R84396 out.n4904 out.n4056 0.003
R84397 out.n4906 out.n3997 0.003
R84398 out.n4942 out.n4920 0.003
R84399 out.n8796 out.n4911 0.003
R84400 out.n919 out.n878 0.003
R84401 out.n8799 out.n920 0.003
R84402 out.n858 out.n834 0.003
R84403 out.n8802 out.n860 0.003
R84404 out.n8805 out.n799 0.003
R84405 out.n8808 out.n793 0.003
R84406 out.n8811 out.n735 0.003
R84407 out.n729 out.n712 0.003
R84408 out.n8814 out.n730 0.003
R84409 out.n705 out.n685 0.003
R84410 out.n8817 out.n673 0.003
R84411 out.n8819 out.n666 0.003
R84412 out.n8822 out.n609 0.003
R84413 out.n8825 out.n603 0.003
R84414 out.n8827 out.n542 0.003
R84415 out.n8830 out.n535 0.003
R84416 out.n8833 out.n480 0.003
R84417 out.n8836 out.n474 0.003
R84418 out.n8839 out.n415 0.003
R84419 out.n409 out.n387 0.003
R84420 out.n8842 out.n410 0.003
R84421 out.n381 out.n363 0.003
R84422 out.n8844 out.n352 0.003
R84423 out.n344 out.n321 0.003
R84424 out.n8846 out.n345 0.003
R84425 out.n313 out.n294 0.003
R84426 out.n8848 out.n282 0.003
R84427 out.n8851 out.n275 0.003
R84428 out.n251 out.n233 0.003
R84429 out.n8854 out.n221 0.003
R84430 out.n8857 out.n215 0.003
R84431 out.n8860 out.n156 0.003
R84432 out.n8863 out.n150 0.003
R84433 out.n8866 out.n94 0.003
R84434 out.n88 out.n64 0.003
R84435 out.n8869 out.n89 0.003
R84436 out.n56 out.n27 0.003
R84437 out.n8871 out.n15 0.003
R84438 out.n14 out.n13 0.003
R84439 out.n6672 out.n6671 0.003
R84440 out.n6662 out.n6659 0.003
R84441 out.n6728 out.n6726 0.003
R84442 out.n2169 out.n2168 0.003
R84443 out.n2989 out.n2988 0.003
R84444 out.n6432 out.n6429 0.003
R84445 out.n6346 out.n6345 0.003
R84446 out.n6329 out.n6328 0.003
R84447 out.n6224 out.n6221 0.003
R84448 out.n1993 out.n1990 0.003
R84449 out.n1983 out.n1978 0.003
R84450 out.n1984 out.n1983 0.003
R84451 out.n1976 out.n1973 0.003
R84452 out.n1963 out.n1962 0.003
R84453 out.n1969 out.n1963 0.003
R84454 out.n1959 out.n1954 0.003
R84455 out.n6268 out.n6265 0.003
R84456 out.n1891 out.n1888 0.003
R84457 out.n1905 out.n1904 0.003
R84458 out.n1914 out.n1913 0.003
R84459 out.n1921 out.n1920 0.003
R84460 out.n6100 out.n6099 0.003
R84461 out.n6057 out.n6054 0.003
R84462 out.n6166 out.n6164 0.003
R84463 out.n1612 out.n1611 0.003
R84464 out.n6994 out.n6991 0.003
R84465 out.n6903 out.n6902 0.003
R84466 out.n6886 out.n6885 0.003
R84467 out.n6781 out.n6778 0.003
R84468 out.n1773 out.n1770 0.003
R84469 out.n1763 out.n1758 0.003
R84470 out.n1764 out.n1763 0.003
R84471 out.n1756 out.n1753 0.003
R84472 out.n1743 out.n1742 0.003
R84473 out.n1749 out.n1743 0.003
R84474 out.n1739 out.n1734 0.003
R84475 out.n6825 out.n6822 0.003
R84476 out.n1666 out.n1663 0.003
R84477 out.n1685 out.n1684 0.003
R84478 out.n1694 out.n1693 0.003
R84479 out.n1701 out.n1700 0.003
R84480 out.n7366 out.n7365 0.003
R84481 out.n7356 out.n7353 0.003
R84482 out.n7432 out.n7430 0.003
R84483 out.n2382 out.n2381 0.003
R84484 out.n7231 out.n7230 0.003
R84485 out.n7136 out.n7135 0.003
R84486 out.n7124 out.n7123 0.003
R84487 out.n2480 out.n2479 0.003
R84488 out.n7095 out.n7091 0.003
R84489 out.n7090 out.n7088 0.003
R84490 out.n7084 out.n7083 0.003
R84491 out.n7206 out.n7203 0.003
R84492 out.n7813 out.n7810 0.003
R84493 out.n7729 out.n7728 0.003
R84494 out.n7712 out.n7711 0.003
R84495 out.n7497 out.n7494 0.003
R84496 out.n7540 out.n7539 0.003
R84497 out.n7621 out.n7620 0.003
R84498 out.n7620 out.n7615 0.003
R84499 out.n7549 out.n7548 0.003
R84500 out.n7559 out.n7558 0.003
R84501 out.n7558 out.n7557 0.003
R84502 out.n7568 out.n7567 0.003
R84503 out.n7672 out.n7669 0.003
R84504 out.n2637 out.n2634 0.003
R84505 out.n2645 out.n2644 0.003
R84506 out.n2653 out.n2652 0.003
R84507 out.n2659 out.n2658 0.003
R84508 out.n2713 out.n2712 0.003
R84509 out.n7009 out.n7002 0.003
R84510 out.n1134 out.n935 0.003
R84511 out.n5611 out.n5610 0.003
R84512 out.n2950 out.n2949 0.003
R84513 out.n5862 out.n5628 0.003
R84514 out.n9432 out.n9427 0.003
R84515 out.n9445 out.n9427 0.003
R84516 out.n9443 out.n9434 0.003
R84517 out.n6998 out.n6997 0.003
R84518 out.n5624 out.n5623 0.003
R84519 out.n9461 out.n9447 0.003
R84520 out.n6442 out.n6441 0.003
R84521 out.n3038 out.n3037 0.003
R84522 out.n1532 out.n1531 0.003
R84523 out.n2379 out.n2378 0.003
R84524 out.n9506 out.n9504 0.003
R84525 out.n14566 out.n14565 0.003
R84526 out.n17185 out.n17173 0.003
R84527 out.n17185 out.n17181 0.003
R84528 out.n17185 out.n17150 0.003
R84529 out.n9506 out.n9489 0.003
R84530 out.n17309 out.n17308 0.003
R84531 out.n11135 out.n11134 0.003
R84532 out.n11558 out.n11557 0.003
R84533 out.n9540 out.n9527 0.003
R84534 out.n9576 out.n9563 0.003
R84535 out.n9612 out.n9599 0.003
R84536 out.n9651 out.n9638 0.003
R84537 out.n9707 out.n9694 0.003
R84538 out.n9743 out.n9730 0.003
R84539 out.n9779 out.n9766 0.003
R84540 out.n9815 out.n9802 0.003
R84541 out.n9851 out.n9838 0.003
R84542 out.n9890 out.n9877 0.003
R84543 out.n9958 out.n9943 0.003
R84544 out.n9958 out.n9945 0.003
R84545 out.n9994 out.n9981 0.003
R84546 out.n16349 out.n16336 0.003
R84547 out.n16417 out.n16402 0.003
R84548 out.n16417 out.n16404 0.003
R84549 out.n16483 out.n16468 0.003
R84550 out.n16483 out.n16470 0.003
R84551 out.n16584 out.n16572 0.003
R84552 out.n16547 out.n16534 0.003
R84553 out.n16648 out.n16638 0.003
R84554 out.n16714 out.n16704 0.003
R84555 out.n16782 out.n16770 0.003
R84556 out.n16782 out.n16772 0.003
R84557 out.n16848 out.n16836 0.003
R84558 out.n16848 out.n16838 0.003
R84559 out.n16912 out.n16902 0.003
R84560 out.n16980 out.n16968 0.003
R84561 out.n16980 out.n16970 0.003
R84562 out.n17044 out.n17034 0.003
R84563 out.n17142 out.n17126 0.003
R84564 out.n17110 out.n17100 0.003
R84565 out.n15641 out.n15640 0.003
R84566 out.n3039 out.n2961 0.002
R84567 out.n10288 out.n10286 0.002
R84568 out.n7824 out.n5614 0.002
R84569 out.n7825 out.n7824 0.002
R84570 out.n7901 out.n7865 0.002
R84571 out.n7902 out.n7901 0.002
R84572 out.n7978 out.n7942 0.002
R84573 out.n7979 out.n7978 0.002
R84574 out.n8055 out.n8019 0.002
R84575 out.n8056 out.n8055 0.002
R84576 out.n8132 out.n8096 0.002
R84577 out.n8133 out.n8132 0.002
R84578 out.n8209 out.n8173 0.002
R84579 out.n8210 out.n8209 0.002
R84580 out.n8286 out.n8250 0.002
R84581 out.n8287 out.n8286 0.002
R84582 out.n8363 out.n8327 0.002
R84583 out.n8364 out.n8363 0.002
R84584 out.n8440 out.n8404 0.002
R84585 out.n8441 out.n8440 0.002
R84586 out.n8517 out.n8481 0.002
R84587 out.n8518 out.n8517 0.002
R84588 out.n8594 out.n8558 0.002
R84589 out.n8595 out.n8594 0.002
R84590 out.n8671 out.n8635 0.002
R84591 out.n8672 out.n8671 0.002
R84592 out.n8748 out.n8712 0.002
R84593 out.n8749 out.n8748 0.002
R84594 out.n3991 out.n3970 0.002
R84595 out.n3931 out.n3930 0.002
R84596 out.n3930 out.n3893 0.002
R84597 out.n3854 out.n3853 0.002
R84598 out.n3853 out.n3816 0.002
R84599 out.n3777 out.n3776 0.002
R84600 out.n3776 out.n3739 0.002
R84601 out.n3700 out.n3699 0.002
R84602 out.n3699 out.n3662 0.002
R84603 out.n3623 out.n3622 0.002
R84604 out.n3622 out.n3585 0.002
R84605 out.n3546 out.n3545 0.002
R84606 out.n3545 out.n3508 0.002
R84607 out.n3469 out.n3468 0.002
R84608 out.n3468 out.n3431 0.002
R84609 out.n3392 out.n3391 0.002
R84610 out.n3391 out.n3354 0.002
R84611 out.n3315 out.n3314 0.002
R84612 out.n3314 out.n3277 0.002
R84613 out.n3199 out.n3198 0.002
R84614 out.n3198 out.n3185 0.002
R84615 out.n3158 out.n3157 0.002
R84616 out.n3157 out.n3079 0.002
R84617 out.n3040 out.n3039 0.002
R84618 out.n8879 out.n8872 0.002
R84619 out.n9506 out.n9475 0.002
R84620 out.n13248 out.n13247 0.002
R84621 out.n17308 out.n9020 0.002
R84622 out.n9506 out.n9498 0.002
R84623 out.n1130 out.n1129 0.002
R84624 out.n9444 out.n9433 0.002
R84625 out.n9459 out.n9458 0.002
R84626 out.n9440 out.n9432 0.002
R84627 out.n10278 out.n10277 0.002
R84628 out.n10263 out.n10262 0.002
R84629 out.n10148 out.n10147 0.002
R84630 out.n12534 out.n12531 0.002
R84631 out.n13367 out.n13364 0.002
R84632 out.n13822 out.n13819 0.002
R84633 out.n14543 out.n14542 0.002
R84634 out.n15909 out.n15907 0.002
R84635 out.n15165 out.n15164 0.002
R84636 out.n16203 out.n16202 0.002
R84637 out.n15565 out.n15564 0.002
R84638 out.n8964 out.n8955 0.002
R84639 out.n10035 out.n10034 0.002
R84640 out.n16014 out.n15999 0.002
R84641 out.n16273 out.n16272 0.002
R84642 out.n10029 out.n10028 0.002
R84643 out.n16278 out.n16277 0.002
R84644 out.n10024 out.n10023 0.002
R84645 out.n10015 out.n10014 0.002
R84646 out.n10019 out.n10018 0.002
R84647 out.n9020 out.n9019 0.002
R84648 out.n12824 out.n12823 0.002
R84649 out.n11556 out.n11555 0.002
R84650 out.n16282 out.n16281 0.002
R84651 out.n10006 out.n10005 0.002
R84652 out.n5168 out.n5167 0.002
R84653 out.n5699 out.n5695 0.002
R84654 out.n5694 out.n5692 0.002
R84655 out.n5822 out.n5819 0.002
R84656 out.n5578 out.n5575 0.002
R84657 out.n3161 out.n3160 0.002
R84658 out.n6732 out.n6729 0.002
R84659 out.n2170 out.n2169 0.002
R84660 out.n3231 out.n3230 0.002
R84661 out.n6764 out.n6763 0.002
R84662 out.n6276 out.n6272 0.002
R84663 out.n6271 out.n6269 0.002
R84664 out.n6394 out.n6391 0.002
R84665 out.n1613 out.n1612 0.002
R84666 out.n6833 out.n6829 0.002
R84667 out.n6828 out.n6826 0.002
R84668 out.n6956 out.n6953 0.002
R84669 out.n7436 out.n7433 0.002
R84670 out.n3211 out.n3210 0.002
R84671 out.n7680 out.n7676 0.002
R84672 out.n7675 out.n7673 0.002
R84673 out.n7777 out.n7774 0.002
R84674 out.n2714 out.n2713 0.002
R84675 out.n3144 out.n3143 0.002
R84676 out.n7817 out.n7816 0.002
R84677 out.n2968 out.n2967 0.002
R84678 out.n6434 out.n6433 0.002
R84679 out.n6996 out.n6995 0.002
R84680 out.n7460 out.n7459 0.002
R84681 out.n5857 out.n5633 0.002
R84682 out.n5602 out.n5601 0.002
R84683 out.n5386 out.n5385 0.002
R84684 out.n3037 out.n3036 0.002
R84685 out.n3035 out.n3033 0.002
R84686 out.n878 out.n876 0.002
R84687 out.n3029 out.n3028 0.002
R84688 out.n2948 out.n2947 0.002
R84689 out.n9465 out.n9425 0.002
R84690 out.n2961 out.n2960 0.002
R84691 out.n9506 out.n9485 0.002
R84692 out.n9506 out.n9481 0.002
R84693 out.n3086 out.n3085 0.002
R84694 out.n12826 out.n12825 0.002
R84695 out.n13247 out.n13246 0.002
R84696 out.n14100 out.n14099 0.002
R84697 out.n13673 out.n13672 0.002
R84698 out.n15413 out.n15412 0.002
R84699 out.n15457 out.n15456 0.002
R84700 out.n9507 out.n9469 0.002
R84701 out.n17185 out.n17176 0.002
R84702 out.n3993 out.n3991 0.002
R84703 out.n119 out.n111 0.002
R84704 out.n185 out.n176 0.002
R84705 out.n251 out.n243 0.002
R84706 out.n313 out.n303 0.002
R84707 out.n381 out.n372 0.002
R84708 out.n444 out.n435 0.002
R84709 out.n511 out.n501 0.002
R84710 out.n572 out.n561 0.002
R84711 out.n638 out.n629 0.002
R84712 out.n705 out.n695 0.002
R84713 out.n768 out.n754 0.002
R84714 out.n828 out.n817 0.002
R84715 out.n919 out.n895 0.002
R84716 out.n4026 out.n4017 0.002
R84717 out.n4092 out.n4083 0.002
R84718 out.n4155 out.n4144 0.002
R84719 out.n4219 out.n4210 0.002
R84720 out.n4282 out.n4274 0.002
R84721 out.n4349 out.n4338 0.002
R84722 out.n4414 out.n4404 0.002
R84723 out.n4478 out.n4469 0.002
R84724 out.n4541 out.n4531 0.002
R84725 out.n4609 out.n4599 0.002
R84726 out.n4673 out.n4664 0.002
R84727 out.n4737 out.n4728 0.002
R84728 out.n4800 out.n4789 0.002
R84729 out.n16233 out.n16232 0.002
R84730 out.n3079 out.n3077 0.002
R84731 out.n3077 out.n3040 0.002
R84732 out.n3185 out.n3183 0.002
R84733 out.n3183 out.n3158 0.002
R84734 out.n3277 out.n3275 0.002
R84735 out.n3275 out.n3199 0.002
R84736 out.n3354 out.n3352 0.002
R84737 out.n3352 out.n3315 0.002
R84738 out.n3431 out.n3429 0.002
R84739 out.n3429 out.n3392 0.002
R84740 out.n3508 out.n3506 0.002
R84741 out.n3506 out.n3469 0.002
R84742 out.n3585 out.n3583 0.002
R84743 out.n3583 out.n3546 0.002
R84744 out.n3662 out.n3660 0.002
R84745 out.n3660 out.n3623 0.002
R84746 out.n3739 out.n3737 0.002
R84747 out.n3737 out.n3700 0.002
R84748 out.n3816 out.n3814 0.002
R84749 out.n3814 out.n3777 0.002
R84750 out.n3893 out.n3891 0.002
R84751 out.n3891 out.n3854 0.002
R84752 out.n3970 out.n3968 0.002
R84753 out.n3968 out.n3931 0.002
R84754 out.n8796 out.n8749 0.002
R84755 out.n8710 out.n8672 0.002
R84756 out.n8712 out.n8710 0.002
R84757 out.n8633 out.n8595 0.002
R84758 out.n8635 out.n8633 0.002
R84759 out.n8556 out.n8518 0.002
R84760 out.n8558 out.n8556 0.002
R84761 out.n8479 out.n8441 0.002
R84762 out.n8481 out.n8479 0.002
R84763 out.n8402 out.n8364 0.002
R84764 out.n8404 out.n8402 0.002
R84765 out.n8325 out.n8287 0.002
R84766 out.n8327 out.n8325 0.002
R84767 out.n8248 out.n8210 0.002
R84768 out.n8250 out.n8248 0.002
R84769 out.n8171 out.n8133 0.002
R84770 out.n8173 out.n8171 0.002
R84771 out.n8094 out.n8056 0.002
R84772 out.n8096 out.n8094 0.002
R84773 out.n8017 out.n7979 0.002
R84774 out.n8019 out.n8017 0.002
R84775 out.n7940 out.n7902 0.002
R84776 out.n7942 out.n7940 0.002
R84777 out.n7863 out.n7825 0.002
R84778 out.n7865 out.n7863 0.002
R84779 out.n5614 out.n5612 0.002
R84780 out.n4838 out.n4802 0.002
R84781 out.n2970 out.n2969 0.002
R84782 out.n56 out.n46 0.002
R84783 out.n15455 out.n15436 0.002
R84784 out.n14103 out.n11137 0.002
R84785 out.n14103 out.n11559 0.002
R84786 out.n15426 out.n15417 0.002
R84787 out.n14147 out.n14126 0.002
R84788 out.n14147 out.n14127 0.002
R84789 out.n14598 out.n14576 0.002
R84790 out.n14598 out.n14577 0.002
R84791 out.n14634 out.n14614 0.002
R84792 out.n14634 out.n14615 0.002
R84793 out.n14669 out.n14649 0.002
R84794 out.n14669 out.n14650 0.002
R84795 out.n14705 out.n14685 0.002
R84796 out.n14705 out.n14686 0.002
R84797 out.n14740 out.n14720 0.002
R84798 out.n14740 out.n14721 0.002
R84799 out.n14776 out.n14756 0.002
R84800 out.n14776 out.n14757 0.002
R84801 out.n14811 out.n14791 0.002
R84802 out.n14811 out.n14792 0.002
R84803 out.n14847 out.n14827 0.002
R84804 out.n14847 out.n14828 0.002
R84805 out.n14882 out.n14862 0.002
R84806 out.n14882 out.n14863 0.002
R84807 out.n14918 out.n14898 0.002
R84808 out.n14918 out.n14899 0.002
R84809 out.n14953 out.n14933 0.002
R84810 out.n14953 out.n14934 0.002
R84811 out.n14989 out.n14969 0.002
R84812 out.n14989 out.n14970 0.002
R84813 out.n15021 out.n15001 0.002
R84814 out.n15021 out.n15002 0.002
R84815 out.n15054 out.n15034 0.002
R84816 out.n15054 out.n15035 0.002
R84817 out.n15086 out.n15066 0.002
R84818 out.n15086 out.n15067 0.002
R84819 out.n15119 out.n15099 0.002
R84820 out.n15119 out.n15100 0.002
R84821 out.n8929 out.n8906 0.002
R84822 out.n8929 out.n8907 0.002
R84823 out.n15157 out.n15137 0.002
R84824 out.n15157 out.n15138 0.002
R84825 out.n8964 out.n8943 0.002
R84826 out.n8964 out.n8944 0.002
R84827 out.n15198 out.n15177 0.002
R84828 out.n15198 out.n15178 0.002
R84829 out.n15229 out.n15209 0.002
R84830 out.n15229 out.n15210 0.002
R84831 out.n15263 out.n15243 0.002
R84832 out.n15263 out.n15244 0.002
R84833 out.n15294 out.n15274 0.002
R84834 out.n15294 out.n15275 0.002
R84835 out.n15328 out.n15308 0.002
R84836 out.n15328 out.n15309 0.002
R84837 out.n15359 out.n15339 0.002
R84838 out.n15359 out.n15340 0.002
R84839 out.n9015 out.n8995 0.002
R84840 out.n16263 out.n16243 0.002
R84841 out.n16263 out.n16245 0.002
R84842 out.n16231 out.n16214 0.002
R84843 out.n16231 out.n16216 0.002
R84844 out.n17277 out.n17253 0.002
R84845 out.n17277 out.n17255 0.002
R84846 out.n16196 out.n16179 0.002
R84847 out.n16196 out.n16181 0.002
R84848 out.n16166 out.n16146 0.002
R84849 out.n16166 out.n16148 0.002
R84850 out.n16135 out.n16118 0.002
R84851 out.n16135 out.n16120 0.002
R84852 out.n16105 out.n16085 0.002
R84853 out.n16105 out.n16087 0.002
R84854 out.n16073 out.n16056 0.002
R84855 out.n16073 out.n16058 0.002
R84856 out.n15978 out.n15954 0.002
R84857 out.n15978 out.n15956 0.002
R84858 out.n15935 out.n15918 0.002
R84859 out.n15935 out.n15920 0.002
R84860 out.n16014 out.n15990 0.002
R84861 out.n16014 out.n15992 0.002
R84862 out.n15899 out.n15882 0.002
R84863 out.n15899 out.n15884 0.002
R84864 out.n15869 out.n15849 0.002
R84865 out.n15869 out.n15851 0.002
R84866 out.n15838 out.n15821 0.002
R84867 out.n15838 out.n15823 0.002
R84868 out.n15808 out.n15788 0.002
R84869 out.n15808 out.n15790 0.002
R84870 out.n15777 out.n15760 0.002
R84871 out.n15777 out.n15762 0.002
R84872 out.n15747 out.n15727 0.002
R84873 out.n15747 out.n15729 0.002
R84874 out.n15711 out.n15694 0.002
R84875 out.n15711 out.n15696 0.002
R84876 out.n15676 out.n15656 0.002
R84877 out.n15676 out.n15658 0.002
R84878 out.n15639 out.n15622 0.002
R84879 out.n15639 out.n15624 0.002
R84880 out.n15605 out.n15581 0.002
R84881 out.n15605 out.n15583 0.002
R84882 out.n15558 out.n15541 0.002
R84883 out.n15558 out.n15543 0.002
R84884 out.n15528 out.n15508 0.002
R84885 out.n15528 out.n15510 0.002
R84886 out.n15492 out.n15474 0.002
R84887 out.n15492 out.n15476 0.002
R84888 out.n15455 out.n15438 0.002
R84889 out.n15426 out.n15421 0.002
R84890 out.n12400 out.n12399 0.002
R84891 out.n12396 out.n12395 0.002
R84892 out.n10290 out.n10289 0.002
R84893 out.n15455 out.n15396 0.002
R84894 out.n15426 out.n15409 0.002
R84895 out.n14103 out.n12827 0.002
R84896 out.n14103 out.n12828 0.002
R84897 out.n14147 out.n14134 0.002
R84898 out.n14147 out.n14138 0.002
R84899 out.n14598 out.n14585 0.002
R84900 out.n14598 out.n14591 0.002
R84901 out.n14634 out.n14622 0.002
R84902 out.n14634 out.n14626 0.002
R84903 out.n14669 out.n14658 0.002
R84904 out.n14669 out.n14662 0.002
R84905 out.n14705 out.n14693 0.002
R84906 out.n14705 out.n14697 0.002
R84907 out.n14740 out.n14729 0.002
R84908 out.n14740 out.n14733 0.002
R84909 out.n14776 out.n14764 0.002
R84910 out.n14776 out.n14768 0.002
R84911 out.n14811 out.n14800 0.002
R84912 out.n14811 out.n14804 0.002
R84913 out.n14847 out.n14835 0.002
R84914 out.n14847 out.n14839 0.002
R84915 out.n14882 out.n14871 0.002
R84916 out.n14882 out.n14875 0.002
R84917 out.n14918 out.n14906 0.002
R84918 out.n14918 out.n14910 0.002
R84919 out.n14953 out.n14942 0.002
R84920 out.n14953 out.n14946 0.002
R84921 out.n14989 out.n14977 0.002
R84922 out.n14989 out.n14981 0.002
R84923 out.n15021 out.n15010 0.002
R84924 out.n15021 out.n15014 0.002
R84925 out.n15054 out.n15042 0.002
R84926 out.n15054 out.n15046 0.002
R84927 out.n15086 out.n15075 0.002
R84928 out.n15086 out.n15079 0.002
R84929 out.n15119 out.n15107 0.002
R84930 out.n15119 out.n15111 0.002
R84931 out.n8929 out.n8915 0.002
R84932 out.n8929 out.n8922 0.002
R84933 out.n15157 out.n15145 0.002
R84934 out.n15157 out.n15149 0.002
R84935 out.n8964 out.n8952 0.002
R84936 out.n8964 out.n8957 0.002
R84937 out.n15198 out.n15185 0.002
R84938 out.n15198 out.n15190 0.002
R84939 out.n15229 out.n15218 0.002
R84940 out.n15229 out.n15222 0.002
R84941 out.n15263 out.n15251 0.002
R84942 out.n15263 out.n15255 0.002
R84943 out.n15294 out.n15283 0.002
R84944 out.n15294 out.n15287 0.002
R84945 out.n15328 out.n15316 0.002
R84946 out.n15328 out.n15320 0.002
R84947 out.n15359 out.n15348 0.002
R84948 out.n15359 out.n15352 0.002
R84949 out.n9015 out.n9002 0.002
R84950 out.n16263 out.n16250 0.002
R84951 out.n16263 out.n16253 0.002
R84952 out.n16231 out.n16220 0.002
R84953 out.n16231 out.n16223 0.002
R84954 out.n17277 out.n17260 0.002
R84955 out.n17277 out.n17267 0.002
R84956 out.n16196 out.n16185 0.002
R84957 out.n16196 out.n16188 0.002
R84958 out.n16166 out.n16153 0.002
R84959 out.n16166 out.n16156 0.002
R84960 out.n16135 out.n16124 0.002
R84961 out.n16135 out.n16127 0.002
R84962 out.n16105 out.n16092 0.002
R84963 out.n16105 out.n16095 0.002
R84964 out.n16073 out.n16062 0.002
R84965 out.n16073 out.n16065 0.002
R84966 out.n15978 out.n15961 0.002
R84967 out.n15978 out.n15968 0.002
R84968 out.n15935 out.n15924 0.002
R84969 out.n15935 out.n15927 0.002
R84970 out.n16014 out.n15997 0.002
R84971 out.n16014 out.n16004 0.002
R84972 out.n15899 out.n15888 0.002
R84973 out.n15899 out.n15891 0.002
R84974 out.n15869 out.n15856 0.002
R84975 out.n15869 out.n15859 0.002
R84976 out.n15838 out.n15827 0.002
R84977 out.n15838 out.n15830 0.002
R84978 out.n15808 out.n15795 0.002
R84979 out.n15808 out.n15798 0.002
R84980 out.n15777 out.n15766 0.002
R84981 out.n15777 out.n15769 0.002
R84982 out.n15747 out.n15734 0.002
R84983 out.n15747 out.n15737 0.002
R84984 out.n15711 out.n15700 0.002
R84985 out.n15711 out.n15703 0.002
R84986 out.n15676 out.n15663 0.002
R84987 out.n15676 out.n15666 0.002
R84988 out.n15639 out.n15628 0.002
R84989 out.n15639 out.n15631 0.002
R84990 out.n15605 out.n15588 0.002
R84991 out.n15605 out.n15595 0.002
R84992 out.n15558 out.n15547 0.002
R84993 out.n15558 out.n15550 0.002
R84994 out.n15528 out.n15515 0.002
R84995 out.n15528 out.n15518 0.002
R84996 out.n15492 out.n15479 0.002
R84997 out.n15492 out.n15482 0.002
R84998 out.n15455 out.n15450 0.002
R84999 out.n15455 out.n15448 0.002
R85000 out.n15528 out.n15513 0.002
R85001 out.n15605 out.n15586 0.002
R85002 out.n15558 out.n15545 0.002
R85003 out.n15676 out.n15661 0.002
R85004 out.n15639 out.n15626 0.002
R85005 out.n15747 out.n15732 0.002
R85006 out.n15711 out.n15698 0.002
R85007 out.n15808 out.n15793 0.002
R85008 out.n15777 out.n15764 0.002
R85009 out.n15869 out.n15854 0.002
R85010 out.n15838 out.n15825 0.002
R85011 out.n16014 out.n15995 0.002
R85012 out.n15899 out.n15886 0.002
R85013 out.n15978 out.n15959 0.002
R85014 out.n15935 out.n15922 0.002
R85015 out.n16105 out.n16090 0.002
R85016 out.n16073 out.n16060 0.002
R85017 out.n16166 out.n16151 0.002
R85018 out.n16135 out.n16122 0.002
R85019 out.n17277 out.n17258 0.002
R85020 out.n16196 out.n16183 0.002
R85021 out.n16263 out.n16248 0.002
R85022 out.n16231 out.n16218 0.002
R85023 out.n15359 out.n15343 0.002
R85024 out.n15294 out.n15278 0.002
R85025 out.n15328 out.n15311 0.002
R85026 out.n15229 out.n15213 0.002
R85027 out.n15263 out.n15246 0.002
R85028 out.n8964 out.n8947 0.002
R85029 out.n15198 out.n15180 0.002
R85030 out.n8929 out.n8910 0.002
R85031 out.n15157 out.n15140 0.002
R85032 out.n15086 out.n15070 0.002
R85033 out.n15119 out.n15102 0.002
R85034 out.n15021 out.n15005 0.002
R85035 out.n15054 out.n15037 0.002
R85036 out.n14953 out.n14937 0.002
R85037 out.n14989 out.n14972 0.002
R85038 out.n14882 out.n14866 0.002
R85039 out.n14918 out.n14901 0.002
R85040 out.n14811 out.n14795 0.002
R85041 out.n14847 out.n14830 0.002
R85042 out.n14740 out.n14724 0.002
R85043 out.n14776 out.n14759 0.002
R85044 out.n14669 out.n14653 0.002
R85045 out.n14705 out.n14688 0.002
R85046 out.n14598 out.n14580 0.002
R85047 out.n14634 out.n14617 0.002
R85048 out.n14147 out.n14129 0.002
R85049 out.n15528 out.n15520 0.002
R85050 out.n15528 out.n15523 0.002
R85051 out.n15492 out.n15484 0.002
R85052 out.n15605 out.n15597 0.002
R85053 out.n15605 out.n15600 0.002
R85054 out.n15558 out.n15552 0.002
R85055 out.n15558 out.n15554 0.002
R85056 out.n15676 out.n15668 0.002
R85057 out.n15676 out.n15671 0.002
R85058 out.n15639 out.n15633 0.002
R85059 out.n15639 out.n15635 0.002
R85060 out.n15747 out.n15739 0.002
R85061 out.n15747 out.n15742 0.002
R85062 out.n15711 out.n15705 0.002
R85063 out.n15711 out.n15707 0.002
R85064 out.n15808 out.n15800 0.002
R85065 out.n15808 out.n15803 0.002
R85066 out.n15777 out.n15771 0.002
R85067 out.n15777 out.n15773 0.002
R85068 out.n15869 out.n15861 0.002
R85069 out.n15869 out.n15864 0.002
R85070 out.n15838 out.n15832 0.002
R85071 out.n15838 out.n15834 0.002
R85072 out.n16014 out.n16006 0.002
R85073 out.n16014 out.n16009 0.002
R85074 out.n15899 out.n15893 0.002
R85075 out.n15899 out.n15895 0.002
R85076 out.n15978 out.n15970 0.002
R85077 out.n15978 out.n15973 0.002
R85078 out.n15935 out.n15929 0.002
R85079 out.n15935 out.n15931 0.002
R85080 out.n16105 out.n16097 0.002
R85081 out.n16105 out.n16100 0.002
R85082 out.n16073 out.n16067 0.002
R85083 out.n16073 out.n16069 0.002
R85084 out.n16166 out.n16158 0.002
R85085 out.n16166 out.n16161 0.002
R85086 out.n16135 out.n16129 0.002
R85087 out.n16135 out.n16131 0.002
R85088 out.n17277 out.n17269 0.002
R85089 out.n17277 out.n17272 0.002
R85090 out.n16196 out.n16190 0.002
R85091 out.n16196 out.n16192 0.002
R85092 out.n16263 out.n16255 0.002
R85093 out.n16263 out.n16258 0.002
R85094 out.n16231 out.n16225 0.002
R85095 out.n16231 out.n16227 0.002
R85096 out.n15359 out.n15354 0.002
R85097 out.n15359 out.n15355 0.002
R85098 out.n9015 out.n9009 0.002
R85099 out.n15294 out.n15289 0.002
R85100 out.n15294 out.n15290 0.002
R85101 out.n15328 out.n15322 0.002
R85102 out.n15328 out.n15323 0.002
R85103 out.n15229 out.n15224 0.002
R85104 out.n15229 out.n15225 0.002
R85105 out.n15263 out.n15257 0.002
R85106 out.n15263 out.n15258 0.002
R85107 out.n8964 out.n8959 0.002
R85108 out.n8964 out.n8960 0.002
R85109 out.n15198 out.n15192 0.002
R85110 out.n15198 out.n15193 0.002
R85111 out.n8929 out.n8924 0.002
R85112 out.n8929 out.n8925 0.002
R85113 out.n15157 out.n15151 0.002
R85114 out.n15157 out.n15152 0.002
R85115 out.n15086 out.n15081 0.002
R85116 out.n15086 out.n15082 0.002
R85117 out.n15119 out.n15113 0.002
R85118 out.n15119 out.n15114 0.002
R85119 out.n15021 out.n15016 0.002
R85120 out.n15021 out.n15017 0.002
R85121 out.n15054 out.n15048 0.002
R85122 out.n15054 out.n15049 0.002
R85123 out.n14953 out.n14948 0.002
R85124 out.n14953 out.n14949 0.002
R85125 out.n14989 out.n14983 0.002
R85126 out.n14989 out.n14984 0.002
R85127 out.n14882 out.n14877 0.002
R85128 out.n14882 out.n14878 0.002
R85129 out.n14918 out.n14912 0.002
R85130 out.n14918 out.n14913 0.002
R85131 out.n14811 out.n14806 0.002
R85132 out.n14811 out.n14807 0.002
R85133 out.n14847 out.n14841 0.002
R85134 out.n14847 out.n14842 0.002
R85135 out.n14740 out.n14735 0.002
R85136 out.n14740 out.n14736 0.002
R85137 out.n14776 out.n14770 0.002
R85138 out.n14776 out.n14771 0.002
R85139 out.n14669 out.n14664 0.002
R85140 out.n14669 out.n14665 0.002
R85141 out.n14705 out.n14699 0.002
R85142 out.n14705 out.n14700 0.002
R85143 out.n14598 out.n14593 0.002
R85144 out.n14598 out.n14594 0.002
R85145 out.n14634 out.n14628 0.002
R85146 out.n14634 out.n14629 0.002
R85147 out.n14103 out.n13674 0.002
R85148 out.n14103 out.n13675 0.002
R85149 out.n14147 out.n14141 0.002
R85150 out.n14147 out.n14142 0.002
R85151 out.n14103 out.n12397 0.002
R85152 out.n15492 out.n15487 0.002
R85153 out.n15455 out.n15444 0.002
R85154 out.n15426 out.n15415 0.002
R85155 out.n14147 out.n14120 0.002
R85156 out.n14598 out.n14579 0.002
R85157 out.n14634 out.n14608 0.002
R85158 out.n14669 out.n14652 0.002
R85159 out.n14705 out.n14679 0.002
R85160 out.n14740 out.n14723 0.002
R85161 out.n14776 out.n14750 0.002
R85162 out.n14811 out.n14794 0.002
R85163 out.n14847 out.n14821 0.002
R85164 out.n14882 out.n14865 0.002
R85165 out.n14918 out.n14892 0.002
R85166 out.n14953 out.n14936 0.002
R85167 out.n14989 out.n14963 0.002
R85168 out.n15021 out.n15004 0.002
R85169 out.n15054 out.n15028 0.002
R85170 out.n15086 out.n15069 0.002
R85171 out.n15119 out.n15093 0.002
R85172 out.n8929 out.n8909 0.002
R85173 out.n15157 out.n15131 0.002
R85174 out.n8964 out.n8946 0.002
R85175 out.n15198 out.n15171 0.002
R85176 out.n15229 out.n15212 0.002
R85177 out.n15263 out.n15237 0.002
R85178 out.n15294 out.n15277 0.002
R85179 out.n15328 out.n15302 0.002
R85180 out.n15359 out.n15342 0.002
R85181 out.n16263 out.n16246 0.002
R85182 out.n16231 out.n16210 0.002
R85183 out.n17277 out.n17256 0.002
R85184 out.n16196 out.n16175 0.002
R85185 out.n16166 out.n16149 0.002
R85186 out.n16135 out.n16114 0.002
R85187 out.n16105 out.n16088 0.002
R85188 out.n16073 out.n16052 0.002
R85189 out.n15978 out.n15957 0.002
R85190 out.n15935 out.n15914 0.002
R85191 out.n16014 out.n15993 0.002
R85192 out.n15899 out.n15878 0.002
R85193 out.n15869 out.n15852 0.002
R85194 out.n15838 out.n15817 0.002
R85195 out.n15808 out.n15791 0.002
R85196 out.n15777 out.n15756 0.002
R85197 out.n15747 out.n15730 0.002
R85198 out.n15711 out.n15690 0.002
R85199 out.n15676 out.n15659 0.002
R85200 out.n15639 out.n15618 0.002
R85201 out.n15605 out.n15584 0.002
R85202 out.n15558 out.n15537 0.002
R85203 out.n15528 out.n15511 0.002
R85204 out.n15492 out.n15470 0.002
R85205 out.n14147 out.n14122 0.002
R85206 out.n14634 out.n14610 0.002
R85207 out.n14705 out.n14681 0.002
R85208 out.n14776 out.n14752 0.002
R85209 out.n14847 out.n14823 0.002
R85210 out.n14918 out.n14894 0.002
R85211 out.n14989 out.n14965 0.002
R85212 out.n15054 out.n15030 0.002
R85213 out.n15119 out.n15095 0.002
R85214 out.n15157 out.n15133 0.002
R85215 out.n15198 out.n15173 0.002
R85216 out.n15263 out.n15239 0.002
R85217 out.n15328 out.n15304 0.002
R85218 out.n9015 out.n8990 0.002
R85219 out.n16231 out.n16211 0.002
R85220 out.n16196 out.n16176 0.002
R85221 out.n16135 out.n16115 0.002
R85222 out.n16073 out.n16053 0.002
R85223 out.n15935 out.n15915 0.002
R85224 out.n15899 out.n15879 0.002
R85225 out.n15838 out.n15818 0.002
R85226 out.n15777 out.n15757 0.002
R85227 out.n15711 out.n15691 0.002
R85228 out.n15639 out.n15619 0.002
R85229 out.n15558 out.n15538 0.002
R85230 out.n15492 out.n15471 0.002
R85231 out.n15455 out.n15440 0.002
R85232 out.n14103 out.n10714 0.002
R85233 out.n14147 out.n14123 0.002
R85234 out.n14598 out.n14572 0.002
R85235 out.n14634 out.n14611 0.002
R85236 out.n14669 out.n14645 0.002
R85237 out.n14705 out.n14682 0.002
R85238 out.n14740 out.n14716 0.002
R85239 out.n14776 out.n14753 0.002
R85240 out.n14811 out.n14787 0.002
R85241 out.n14847 out.n14824 0.002
R85242 out.n14882 out.n14858 0.002
R85243 out.n14918 out.n14895 0.002
R85244 out.n14953 out.n14929 0.002
R85245 out.n14989 out.n14966 0.002
R85246 out.n15021 out.n14997 0.002
R85247 out.n15054 out.n15031 0.002
R85248 out.n15086 out.n15062 0.002
R85249 out.n15119 out.n15096 0.002
R85250 out.n8929 out.n8902 0.002
R85251 out.n15157 out.n15134 0.002
R85252 out.n8964 out.n8939 0.002
R85253 out.n15198 out.n15174 0.002
R85254 out.n15229 out.n15205 0.002
R85255 out.n15263 out.n15240 0.002
R85256 out.n15294 out.n15270 0.002
R85257 out.n15328 out.n15305 0.002
R85258 out.n15359 out.n15335 0.002
R85259 out.n16263 out.n16240 0.002
R85260 out.n16231 out.n16213 0.002
R85261 out.n17277 out.n17250 0.002
R85262 out.n16196 out.n16178 0.002
R85263 out.n16166 out.n16143 0.002
R85264 out.n16135 out.n16117 0.002
R85265 out.n16105 out.n16082 0.002
R85266 out.n16073 out.n16055 0.002
R85267 out.n15978 out.n15951 0.002
R85268 out.n15935 out.n15917 0.002
R85269 out.n16014 out.n15987 0.002
R85270 out.n15899 out.n15881 0.002
R85271 out.n15869 out.n15846 0.002
R85272 out.n15838 out.n15820 0.002
R85273 out.n15808 out.n15785 0.002
R85274 out.n15777 out.n15759 0.002
R85275 out.n15747 out.n15724 0.002
R85276 out.n15711 out.n15693 0.002
R85277 out.n15676 out.n15653 0.002
R85278 out.n15639 out.n15621 0.002
R85279 out.n15605 out.n15578 0.002
R85280 out.n15558 out.n15540 0.002
R85281 out.n15528 out.n15505 0.002
R85282 out.n15492 out.n15473 0.002
R85283 out.n15455 out.n15442 0.002
R85284 out.n15426 out.n15422 0.002
R85285 out.n14103 out.n11136 0.002
R85286 out.n14598 out.n14574 0.002
R85287 out.n14669 out.n14647 0.002
R85288 out.n14740 out.n14718 0.002
R85289 out.n14811 out.n14789 0.002
R85290 out.n14882 out.n14860 0.002
R85291 out.n14953 out.n14931 0.002
R85292 out.n15021 out.n14999 0.002
R85293 out.n15086 out.n15064 0.002
R85294 out.n8929 out.n8904 0.002
R85295 out.n8964 out.n8941 0.002
R85296 out.n15229 out.n15207 0.002
R85297 out.n15294 out.n15272 0.002
R85298 out.n15359 out.n15337 0.002
R85299 out.n16263 out.n16241 0.002
R85300 out.n17277 out.n17251 0.002
R85301 out.n16166 out.n16144 0.002
R85302 out.n16105 out.n16083 0.002
R85303 out.n15978 out.n15952 0.002
R85304 out.n16014 out.n15988 0.002
R85305 out.n15869 out.n15847 0.002
R85306 out.n15808 out.n15786 0.002
R85307 out.n15747 out.n15725 0.002
R85308 out.n15676 out.n15654 0.002
R85309 out.n15605 out.n15579 0.002
R85310 out.n15528 out.n15506 0.002
R85311 out.n15455 out.n15439 0.002
R85312 out.n15455 out.n15435 0.002
R85313 out.n15455 out.n15452 0.002
R85314 out.n15528 out.n15524 0.002
R85315 out.n15528 out.n15527 0.002
R85316 out.n15492 out.n15489 0.002
R85317 out.n15492 out.n15491 0.002
R85318 out.n15605 out.n15601 0.002
R85319 out.n15605 out.n15604 0.002
R85320 out.n15558 out.n15555 0.002
R85321 out.n15558 out.n15557 0.002
R85322 out.n15676 out.n15672 0.002
R85323 out.n15676 out.n15675 0.002
R85324 out.n15639 out.n15636 0.002
R85325 out.n15639 out.n15638 0.002
R85326 out.n15747 out.n15743 0.002
R85327 out.n15747 out.n15746 0.002
R85328 out.n15711 out.n15708 0.002
R85329 out.n15711 out.n15710 0.002
R85330 out.n15808 out.n15804 0.002
R85331 out.n15808 out.n15807 0.002
R85332 out.n15777 out.n15774 0.002
R85333 out.n15777 out.n15776 0.002
R85334 out.n15869 out.n15865 0.002
R85335 out.n15869 out.n15868 0.002
R85336 out.n15838 out.n15835 0.002
R85337 out.n15838 out.n15837 0.002
R85338 out.n16014 out.n16010 0.002
R85339 out.n16014 out.n16013 0.002
R85340 out.n15899 out.n15896 0.002
R85341 out.n15899 out.n15898 0.002
R85342 out.n15978 out.n15974 0.002
R85343 out.n15978 out.n15977 0.002
R85344 out.n15935 out.n15932 0.002
R85345 out.n15935 out.n15934 0.002
R85346 out.n16105 out.n16101 0.002
R85347 out.n16105 out.n16104 0.002
R85348 out.n16073 out.n16070 0.002
R85349 out.n16073 out.n16072 0.002
R85350 out.n16166 out.n16162 0.002
R85351 out.n16166 out.n16165 0.002
R85352 out.n16135 out.n16132 0.002
R85353 out.n16135 out.n16134 0.002
R85354 out.n17277 out.n17273 0.002
R85355 out.n17277 out.n17276 0.002
R85356 out.n16196 out.n16193 0.002
R85357 out.n16196 out.n16195 0.002
R85358 out.n16263 out.n16259 0.002
R85359 out.n16263 out.n16262 0.002
R85360 out.n16231 out.n16228 0.002
R85361 out.n16231 out.n16230 0.002
R85362 out.n15359 out.n15357 0.002
R85363 out.n15359 out.n15358 0.002
R85364 out.n9015 out.n9013 0.002
R85365 out.n15294 out.n15292 0.002
R85366 out.n15294 out.n15293 0.002
R85367 out.n15328 out.n15326 0.002
R85368 out.n15328 out.n15327 0.002
R85369 out.n15229 out.n15227 0.002
R85370 out.n15229 out.n15228 0.002
R85371 out.n15263 out.n15261 0.002
R85372 out.n15263 out.n15262 0.002
R85373 out.n8964 out.n8962 0.002
R85374 out.n8964 out.n8963 0.002
R85375 out.n15198 out.n15196 0.002
R85376 out.n15198 out.n15197 0.002
R85377 out.n8929 out.n8927 0.002
R85378 out.n8929 out.n8928 0.002
R85379 out.n15157 out.n15155 0.002
R85380 out.n15157 out.n15156 0.002
R85381 out.n15086 out.n15084 0.002
R85382 out.n15086 out.n15085 0.002
R85383 out.n15119 out.n15117 0.002
R85384 out.n15119 out.n15118 0.002
R85385 out.n15021 out.n15019 0.002
R85386 out.n15021 out.n15020 0.002
R85387 out.n15054 out.n15052 0.002
R85388 out.n15054 out.n15053 0.002
R85389 out.n14953 out.n14951 0.002
R85390 out.n14953 out.n14952 0.002
R85391 out.n14989 out.n14987 0.002
R85392 out.n14989 out.n14988 0.002
R85393 out.n14882 out.n14880 0.002
R85394 out.n14882 out.n14881 0.002
R85395 out.n14918 out.n14916 0.002
R85396 out.n14918 out.n14917 0.002
R85397 out.n14811 out.n14809 0.002
R85398 out.n14811 out.n14810 0.002
R85399 out.n14847 out.n14845 0.002
R85400 out.n14847 out.n14846 0.002
R85401 out.n14740 out.n14738 0.002
R85402 out.n14740 out.n14739 0.002
R85403 out.n14776 out.n14774 0.002
R85404 out.n14776 out.n14775 0.002
R85405 out.n14669 out.n14667 0.002
R85406 out.n14669 out.n14668 0.002
R85407 out.n14705 out.n14703 0.002
R85408 out.n14705 out.n14704 0.002
R85409 out.n14598 out.n14596 0.002
R85410 out.n14598 out.n14597 0.002
R85411 out.n14634 out.n14632 0.002
R85412 out.n14634 out.n14633 0.002
R85413 out.n14103 out.n14101 0.002
R85414 out.n14103 out.n14102 0.002
R85415 out.n14147 out.n14145 0.002
R85416 out.n14147 out.n14146 0.002
R85417 out.n14103 out.n10709 0.002
R85418 out.n14147 out.n14117 0.002
R85419 out.n14598 out.n14112 0.002
R85420 out.n14634 out.n14602 0.002
R85421 out.n14669 out.n14639 0.002
R85422 out.n14705 out.n14673 0.002
R85423 out.n14740 out.n14710 0.002
R85424 out.n14776 out.n14744 0.002
R85425 out.n14811 out.n14781 0.002
R85426 out.n14847 out.n14815 0.002
R85427 out.n14882 out.n14852 0.002
R85428 out.n14918 out.n14886 0.002
R85429 out.n14953 out.n14923 0.002
R85430 out.n14989 out.n14957 0.002
R85431 out.n15021 out.n14994 0.002
R85432 out.n15054 out.n15025 0.002
R85433 out.n15086 out.n15059 0.002
R85434 out.n15119 out.n15090 0.002
R85435 out.n8929 out.n8899 0.002
R85436 out.n15157 out.n15128 0.002
R85437 out.n8964 out.n8936 0.002
R85438 out.n15198 out.n15168 0.002
R85439 out.n15229 out.n15202 0.002
R85440 out.n15263 out.n15234 0.002
R85441 out.n15294 out.n15267 0.002
R85442 out.n15328 out.n15299 0.002
R85443 out.n15359 out.n15332 0.002
R85444 out.n9015 out.n8984 0.002
R85445 out.n16263 out.n16237 0.002
R85446 out.n16231 out.n16207 0.002
R85447 out.n17277 out.n17247 0.002
R85448 out.n16196 out.n16172 0.002
R85449 out.n16166 out.n16140 0.002
R85450 out.n16135 out.n16111 0.002
R85451 out.n16105 out.n16079 0.002
R85452 out.n16073 out.n15942 0.002
R85453 out.n15978 out.n15948 0.002
R85454 out.n15935 out.n15911 0.002
R85455 out.n16014 out.n15984 0.002
R85456 out.n15899 out.n15875 0.002
R85457 out.n15869 out.n15843 0.002
R85458 out.n15838 out.n15814 0.002
R85459 out.n15808 out.n15782 0.002
R85460 out.n15777 out.n15753 0.002
R85461 out.n15747 out.n15716 0.002
R85462 out.n15711 out.n15682 0.002
R85463 out.n15676 out.n15645 0.002
R85464 out.n15639 out.n15569 0.002
R85465 out.n15605 out.n15575 0.002
R85466 out.n15558 out.n15534 0.002
R85467 out.n15528 out.n15497 0.002
R85468 out.n15492 out.n15462 0.002
R85469 out.n15455 out.n15393 0.002
R85470 out.n2996 out.n2986 0.002
R85471 out.n3057 out.n3050 0.002
R85472 out.n3222 out.n3219 0.002
R85473 out.n3294 out.n3287 0.002
R85474 out.n3238 out.n3226 0.002
R85475 out.n3371 out.n3364 0.002
R85476 out.n3332 out.n3325 0.002
R85477 out.n3448 out.n3441 0.002
R85478 out.n3409 out.n3402 0.002
R85479 out.n3525 out.n3518 0.002
R85480 out.n3486 out.n3479 0.002
R85481 out.n3602 out.n3595 0.002
R85482 out.n3563 out.n3556 0.002
R85483 out.n3679 out.n3672 0.002
R85484 out.n3640 out.n3633 0.002
R85485 out.n3756 out.n3749 0.002
R85486 out.n3717 out.n3710 0.002
R85487 out.n3833 out.n3826 0.002
R85488 out.n3794 out.n3787 0.002
R85489 out.n3910 out.n3903 0.002
R85490 out.n3871 out.n3864 0.002
R85491 out.n3948 out.n3941 0.002
R85492 out.n8732 out.n8726 0.002
R85493 out.n8775 out.n8765 0.002
R85494 out.n8775 out.n8767 0.002
R85495 out.n8655 out.n8649 0.002
R85496 out.n8692 out.n8686 0.002
R85497 out.n8578 out.n8572 0.002
R85498 out.n8615 out.n8609 0.002
R85499 out.n8501 out.n8495 0.002
R85500 out.n8538 out.n8532 0.002
R85501 out.n8424 out.n8418 0.002
R85502 out.n8461 out.n8455 0.002
R85503 out.n8347 out.n8341 0.002
R85504 out.n8384 out.n8378 0.002
R85505 out.n8270 out.n8264 0.002
R85506 out.n8307 out.n8301 0.002
R85507 out.n8193 out.n8187 0.002
R85508 out.n8230 out.n8224 0.002
R85509 out.n8116 out.n8110 0.002
R85510 out.n8153 out.n8147 0.002
R85511 out.n8039 out.n8033 0.002
R85512 out.n8076 out.n8070 0.002
R85513 out.n7962 out.n7956 0.002
R85514 out.n7999 out.n7993 0.002
R85515 out.n7885 out.n7879 0.002
R85516 out.n7922 out.n7916 0.002
R85517 out.n7845 out.n7839 0.002
R85518 out.n2180 out.n1626 0.002
R85519 out.n3121 out.n3089 0.002
R85520 out.n6767 out.n6197 0.002
R85521 out.n2943 out.n2387 0.002
R85522 out.n3070 out.n3059 0.002
R85523 out.n3023 out.n2998 0.002
R85524 out.n3150 out.n3127 0.002
R85525 out.n3307 out.n3296 0.002
R85526 out.n3268 out.n3240 0.002
R85527 out.n3384 out.n3373 0.002
R85528 out.n3345 out.n3334 0.002
R85529 out.n3461 out.n3450 0.002
R85530 out.n3422 out.n3411 0.002
R85531 out.n3538 out.n3527 0.002
R85532 out.n3499 out.n3488 0.002
R85533 out.n3615 out.n3604 0.002
R85534 out.n3576 out.n3565 0.002
R85535 out.n3692 out.n3681 0.002
R85536 out.n3653 out.n3642 0.002
R85537 out.n3769 out.n3758 0.002
R85538 out.n3730 out.n3719 0.002
R85539 out.n3846 out.n3835 0.002
R85540 out.n3807 out.n3796 0.002
R85541 out.n3923 out.n3912 0.002
R85542 out.n3884 out.n3873 0.002
R85543 out.n3961 out.n3950 0.002
R85544 out.n8744 out.n8736 0.002
R85545 out.n8792 out.n8780 0.002
R85546 out.n8667 out.n8659 0.002
R85547 out.n8706 out.n8696 0.002
R85548 out.n8590 out.n8582 0.002
R85549 out.n8629 out.n8619 0.002
R85550 out.n8513 out.n8505 0.002
R85551 out.n8552 out.n8542 0.002
R85552 out.n8436 out.n8428 0.002
R85553 out.n8475 out.n8465 0.002
R85554 out.n8359 out.n8351 0.002
R85555 out.n8398 out.n8388 0.002
R85556 out.n8282 out.n8274 0.002
R85557 out.n8321 out.n8311 0.002
R85558 out.n8205 out.n8197 0.002
R85559 out.n8244 out.n8234 0.002
R85560 out.n8128 out.n8120 0.002
R85561 out.n8167 out.n8157 0.002
R85562 out.n8051 out.n8043 0.002
R85563 out.n8090 out.n8080 0.002
R85564 out.n7974 out.n7966 0.002
R85565 out.n8013 out.n8003 0.002
R85566 out.n7897 out.n7889 0.002
R85567 out.n7936 out.n7926 0.002
R85568 out.n7820 out.n7468 0.002
R85569 out.n7859 out.n7849 0.002
R85570 out.n3133 out.n3131 0.002
R85571 out.n3252 out.n3250 0.002
R85572 out.n8792 out.n8789 0.002
R85573 out.n7820 out.n7474 0.002
R85574 out.n7859 out.n7853 0.002
R85575 out.n7859 out.n7855 0.002
R85576 out.n7897 out.n7892 0.002
R85577 out.n7936 out.n7930 0.002
R85578 out.n7936 out.n7932 0.002
R85579 out.n7974 out.n7969 0.002
R85580 out.n8013 out.n8007 0.002
R85581 out.n8013 out.n8009 0.002
R85582 out.n8051 out.n8046 0.002
R85583 out.n8090 out.n8084 0.002
R85584 out.n8090 out.n8086 0.002
R85585 out.n8128 out.n8123 0.002
R85586 out.n8167 out.n8161 0.002
R85587 out.n8167 out.n8163 0.002
R85588 out.n8205 out.n8200 0.002
R85589 out.n8244 out.n8238 0.002
R85590 out.n8244 out.n8240 0.002
R85591 out.n8282 out.n8277 0.002
R85592 out.n8321 out.n8315 0.002
R85593 out.n8321 out.n8317 0.002
R85594 out.n8359 out.n8354 0.002
R85595 out.n8398 out.n8392 0.002
R85596 out.n8398 out.n8394 0.002
R85597 out.n8436 out.n8431 0.002
R85598 out.n8475 out.n8469 0.002
R85599 out.n8475 out.n8471 0.002
R85600 out.n8513 out.n8508 0.002
R85601 out.n8552 out.n8546 0.002
R85602 out.n8552 out.n8548 0.002
R85603 out.n8590 out.n8585 0.002
R85604 out.n8629 out.n8623 0.002
R85605 out.n8629 out.n8625 0.002
R85606 out.n8667 out.n8662 0.002
R85607 out.n8706 out.n8700 0.002
R85608 out.n8706 out.n8702 0.002
R85609 out.n8744 out.n8739 0.002
R85610 out.n8792 out.n8785 0.002
R85611 out.n3961 out.n3953 0.002
R85612 out.n3961 out.n3957 0.002
R85613 out.n3923 out.n3915 0.002
R85614 out.n3884 out.n3876 0.002
R85615 out.n3884 out.n3880 0.002
R85616 out.n3846 out.n3838 0.002
R85617 out.n3807 out.n3799 0.002
R85618 out.n3807 out.n3803 0.002
R85619 out.n3769 out.n3761 0.002
R85620 out.n3730 out.n3722 0.002
R85621 out.n3730 out.n3726 0.002
R85622 out.n3692 out.n3684 0.002
R85623 out.n3653 out.n3645 0.002
R85624 out.n3653 out.n3649 0.002
R85625 out.n3615 out.n3607 0.002
R85626 out.n3576 out.n3568 0.002
R85627 out.n3576 out.n3572 0.002
R85628 out.n3538 out.n3530 0.002
R85629 out.n3499 out.n3491 0.002
R85630 out.n3499 out.n3495 0.002
R85631 out.n3461 out.n3453 0.002
R85632 out.n3422 out.n3414 0.002
R85633 out.n3422 out.n3418 0.002
R85634 out.n3384 out.n3376 0.002
R85635 out.n3345 out.n3337 0.002
R85636 out.n3345 out.n3341 0.002
R85637 out.n3307 out.n3299 0.002
R85638 out.n3268 out.n3256 0.002
R85639 out.n3268 out.n3263 0.002
R85640 out.n3150 out.n3138 0.002
R85641 out.n3070 out.n3062 0.002
R85642 out.n3070 out.n3066 0.002
R85643 out.n3023 out.n3007 0.002
R85644 out.n2943 out.n2606 0.002
R85645 out.n2943 out.n2715 0.002
R85646 out.n7820 out.n7469 0.002
R85647 out.n7859 out.n7850 0.002
R85648 out.n7897 out.n7890 0.002
R85649 out.n7936 out.n7927 0.002
R85650 out.n7974 out.n7967 0.002
R85651 out.n8013 out.n8004 0.002
R85652 out.n8051 out.n8044 0.002
R85653 out.n8090 out.n8081 0.002
R85654 out.n8128 out.n8121 0.002
R85655 out.n8167 out.n8158 0.002
R85656 out.n8205 out.n8198 0.002
R85657 out.n8244 out.n8235 0.002
R85658 out.n8282 out.n8275 0.002
R85659 out.n8321 out.n8312 0.002
R85660 out.n8359 out.n8352 0.002
R85661 out.n8398 out.n8389 0.002
R85662 out.n8436 out.n8429 0.002
R85663 out.n8475 out.n8466 0.002
R85664 out.n8513 out.n8506 0.002
R85665 out.n8552 out.n8543 0.002
R85666 out.n8590 out.n8583 0.002
R85667 out.n8629 out.n8620 0.002
R85668 out.n8667 out.n8660 0.002
R85669 out.n8706 out.n8697 0.002
R85670 out.n8744 out.n8737 0.002
R85671 out.n8792 out.n8782 0.002
R85672 out.n3984 out.n3975 0.002
R85673 out.n3961 out.n3952 0.002
R85674 out.n3923 out.n3914 0.002
R85675 out.n3884 out.n3875 0.002
R85676 out.n3846 out.n3837 0.002
R85677 out.n3807 out.n3798 0.002
R85678 out.n3769 out.n3760 0.002
R85679 out.n3730 out.n3721 0.002
R85680 out.n3692 out.n3683 0.002
R85681 out.n3653 out.n3644 0.002
R85682 out.n3615 out.n3606 0.002
R85683 out.n3576 out.n3567 0.002
R85684 out.n3538 out.n3529 0.002
R85685 out.n3499 out.n3490 0.002
R85686 out.n3461 out.n3452 0.002
R85687 out.n3422 out.n3413 0.002
R85688 out.n3384 out.n3375 0.002
R85689 out.n3345 out.n3336 0.002
R85690 out.n3307 out.n3298 0.002
R85691 out.n3268 out.n3255 0.002
R85692 out.n3150 out.n3129 0.002
R85693 out.n3070 out.n3061 0.002
R85694 out.n3023 out.n3006 0.002
R85695 out.n2943 out.n2600 0.002
R85696 out.n6767 out.n5866 0.002
R85697 out.n7845 out.n7833 0.002
R85698 out.n7885 out.n7873 0.002
R85699 out.n7922 out.n7910 0.002
R85700 out.n7962 out.n7950 0.002
R85701 out.n7999 out.n7987 0.002
R85702 out.n8039 out.n8027 0.002
R85703 out.n8076 out.n8064 0.002
R85704 out.n8116 out.n8104 0.002
R85705 out.n8153 out.n8141 0.002
R85706 out.n8193 out.n8181 0.002
R85707 out.n8230 out.n8218 0.002
R85708 out.n8270 out.n8258 0.002
R85709 out.n8307 out.n8295 0.002
R85710 out.n8347 out.n8335 0.002
R85711 out.n8384 out.n8372 0.002
R85712 out.n8424 out.n8412 0.002
R85713 out.n8461 out.n8449 0.002
R85714 out.n8501 out.n8489 0.002
R85715 out.n8538 out.n8526 0.002
R85716 out.n8578 out.n8566 0.002
R85717 out.n8615 out.n8603 0.002
R85718 out.n8655 out.n8643 0.002
R85719 out.n8692 out.n8680 0.002
R85720 out.n8732 out.n8720 0.002
R85721 out.n907 out.n897 0.002
R85722 out.n3948 out.n3935 0.002
R85723 out.n3910 out.n3897 0.002
R85724 out.n3871 out.n3858 0.002
R85725 out.n3833 out.n3820 0.002
R85726 out.n3794 out.n3781 0.002
R85727 out.n3756 out.n3743 0.002
R85728 out.n3717 out.n3704 0.002
R85729 out.n3679 out.n3666 0.002
R85730 out.n3640 out.n3627 0.002
R85731 out.n3602 out.n3589 0.002
R85732 out.n3563 out.n3550 0.002
R85733 out.n3525 out.n3512 0.002
R85734 out.n3486 out.n3473 0.002
R85735 out.n3448 out.n3435 0.002
R85736 out.n3409 out.n3396 0.002
R85737 out.n3371 out.n3358 0.002
R85738 out.n3332 out.n3319 0.002
R85739 out.n3294 out.n3281 0.002
R85740 out.n3238 out.n3203 0.002
R85741 out.n3222 out.n3209 0.002
R85742 out.n3121 out.n3083 0.002
R85743 out.n3057 out.n3044 0.002
R85744 out.n2996 out.n2971 0.002
R85745 out.n2180 out.n1620 0.002
R85746 out.n7820 out.n7818 0.002
R85747 out.n7820 out.n7819 0.002
R85748 out.n7859 out.n7857 0.002
R85749 out.n7859 out.n7858 0.002
R85750 out.n7897 out.n7895 0.002
R85751 out.n7897 out.n7896 0.002
R85752 out.n7936 out.n7934 0.002
R85753 out.n7936 out.n7935 0.002
R85754 out.n7974 out.n7972 0.002
R85755 out.n7974 out.n7973 0.002
R85756 out.n8013 out.n8011 0.002
R85757 out.n8013 out.n8012 0.002
R85758 out.n8051 out.n8049 0.002
R85759 out.n8051 out.n8050 0.002
R85760 out.n8090 out.n8088 0.002
R85761 out.n8090 out.n8089 0.002
R85762 out.n8128 out.n8126 0.002
R85763 out.n8128 out.n8127 0.002
R85764 out.n8167 out.n8165 0.002
R85765 out.n8167 out.n8166 0.002
R85766 out.n8205 out.n8203 0.002
R85767 out.n8205 out.n8204 0.002
R85768 out.n8244 out.n8242 0.002
R85769 out.n8244 out.n8243 0.002
R85770 out.n8282 out.n8280 0.002
R85771 out.n8282 out.n8281 0.002
R85772 out.n8321 out.n8319 0.002
R85773 out.n8321 out.n8320 0.002
R85774 out.n8359 out.n8357 0.002
R85775 out.n8359 out.n8358 0.002
R85776 out.n8398 out.n8396 0.002
R85777 out.n8398 out.n8397 0.002
R85778 out.n8436 out.n8434 0.002
R85779 out.n8436 out.n8435 0.002
R85780 out.n8475 out.n8473 0.002
R85781 out.n8475 out.n8474 0.002
R85782 out.n8513 out.n8511 0.002
R85783 out.n8513 out.n8512 0.002
R85784 out.n8552 out.n8550 0.002
R85785 out.n8552 out.n8551 0.002
R85786 out.n8590 out.n8588 0.002
R85787 out.n8590 out.n8589 0.002
R85788 out.n8629 out.n8627 0.002
R85789 out.n8629 out.n8628 0.002
R85790 out.n8667 out.n8665 0.002
R85791 out.n8667 out.n8666 0.002
R85792 out.n8706 out.n8704 0.002
R85793 out.n8706 out.n8705 0.002
R85794 out.n8744 out.n8742 0.002
R85795 out.n8744 out.n8743 0.002
R85796 out.n8792 out.n8791 0.002
R85797 out.n3984 out.n3983 0.002
R85798 out.n3961 out.n3958 0.002
R85799 out.n3961 out.n3960 0.002
R85800 out.n3923 out.n3920 0.002
R85801 out.n3923 out.n3922 0.002
R85802 out.n3884 out.n3881 0.002
R85803 out.n3884 out.n3883 0.002
R85804 out.n3846 out.n3843 0.002
R85805 out.n3846 out.n3845 0.002
R85806 out.n3807 out.n3804 0.002
R85807 out.n3807 out.n3806 0.002
R85808 out.n3769 out.n3766 0.002
R85809 out.n3769 out.n3768 0.002
R85810 out.n3730 out.n3727 0.002
R85811 out.n3730 out.n3729 0.002
R85812 out.n3692 out.n3689 0.002
R85813 out.n3692 out.n3691 0.002
R85814 out.n3653 out.n3650 0.002
R85815 out.n3653 out.n3652 0.002
R85816 out.n3615 out.n3612 0.002
R85817 out.n3615 out.n3614 0.002
R85818 out.n3576 out.n3573 0.002
R85819 out.n3576 out.n3575 0.002
R85820 out.n3538 out.n3535 0.002
R85821 out.n3538 out.n3537 0.002
R85822 out.n3499 out.n3496 0.002
R85823 out.n3499 out.n3498 0.002
R85824 out.n3461 out.n3458 0.002
R85825 out.n3461 out.n3460 0.002
R85826 out.n3422 out.n3419 0.002
R85827 out.n3422 out.n3421 0.002
R85828 out.n3384 out.n3381 0.002
R85829 out.n3384 out.n3383 0.002
R85830 out.n3345 out.n3342 0.002
R85831 out.n3345 out.n3344 0.002
R85832 out.n3307 out.n3304 0.002
R85833 out.n3307 out.n3306 0.002
R85834 out.n3268 out.n3264 0.002
R85835 out.n3268 out.n3267 0.002
R85836 out.n3252 out.n3251 0.002
R85837 out.n3150 out.n3147 0.002
R85838 out.n3150 out.n3149 0.002
R85839 out.n3070 out.n3067 0.002
R85840 out.n3070 out.n3069 0.002
R85841 out.n3023 out.n3018 0.002
R85842 out.n3023 out.n3022 0.002
R85843 out.n2943 out.n2723 0.002
R85844 out.n2943 out.n2942 0.002
R85845 out.n15426 out.n15418 0.002
R85846 out.n15426 out.n15425 0.002
R85847 out.n6191 out.n6190 0.001
R85848 out.n14103 out.n12398 0.001
R85849 out.n14147 out.n14131 0.001
R85850 out.n14598 out.n14583 0.001
R85851 out.n14634 out.n14620 0.001
R85852 out.n14669 out.n14656 0.001
R85853 out.n14705 out.n14691 0.001
R85854 out.n14740 out.n14727 0.001
R85855 out.n14776 out.n14762 0.001
R85856 out.n14811 out.n14798 0.001
R85857 out.n14847 out.n14833 0.001
R85858 out.n14882 out.n14869 0.001
R85859 out.n14918 out.n14904 0.001
R85860 out.n14953 out.n14940 0.001
R85861 out.n14989 out.n14975 0.001
R85862 out.n15021 out.n15008 0.001
R85863 out.n15054 out.n15040 0.001
R85864 out.n15086 out.n15073 0.001
R85865 out.n15119 out.n15105 0.001
R85866 out.n8929 out.n8913 0.001
R85867 out.n15157 out.n15143 0.001
R85868 out.n8964 out.n8950 0.001
R85869 out.n15198 out.n15183 0.001
R85870 out.n15229 out.n15216 0.001
R85871 out.n15263 out.n15249 0.001
R85872 out.n15294 out.n15281 0.001
R85873 out.n15328 out.n15314 0.001
R85874 out.n15359 out.n15346 0.001
R85875 out.n9015 out.n9000 0.001
R85876 out.n16263 out.n16249 0.001
R85877 out.n16231 out.n16219 0.001
R85878 out.n17277 out.n17259 0.001
R85879 out.n16196 out.n16184 0.001
R85880 out.n16166 out.n16152 0.001
R85881 out.n16135 out.n16123 0.001
R85882 out.n16105 out.n16091 0.001
R85883 out.n16073 out.n16061 0.001
R85884 out.n15978 out.n15960 0.001
R85885 out.n15935 out.n15923 0.001
R85886 out.n16014 out.n15996 0.001
R85887 out.n15899 out.n15887 0.001
R85888 out.n15869 out.n15855 0.001
R85889 out.n15838 out.n15826 0.001
R85890 out.n15808 out.n15794 0.001
R85891 out.n15777 out.n15765 0.001
R85892 out.n15747 out.n15733 0.001
R85893 out.n15711 out.n15699 0.001
R85894 out.n15676 out.n15662 0.001
R85895 out.n15639 out.n15627 0.001
R85896 out.n15605 out.n15587 0.001
R85897 out.n15558 out.n15546 0.001
R85898 out.n15528 out.n15514 0.001
R85899 out.n15492 out.n15478 0.001
R85900 out.n15455 out.n15451 0.001
R85901 out.n15455 out.n15446 0.001
R85902 out.n2180 out.n1852 0.001
R85903 out.n2996 out.n2984 0.001
R85904 out.n3121 out.n3093 0.001
R85905 out.n3057 out.n3048 0.001
R85906 out.n3222 out.n3218 0.001
R85907 out.n3294 out.n3285 0.001
R85908 out.n3238 out.n3224 0.001
R85909 out.n3371 out.n3362 0.001
R85910 out.n3332 out.n3323 0.001
R85911 out.n3448 out.n3439 0.001
R85912 out.n3409 out.n3400 0.001
R85913 out.n3525 out.n3516 0.001
R85914 out.n3486 out.n3477 0.001
R85915 out.n3602 out.n3593 0.001
R85916 out.n3563 out.n3554 0.001
R85917 out.n3679 out.n3670 0.001
R85918 out.n3640 out.n3631 0.001
R85919 out.n3756 out.n3747 0.001
R85920 out.n3717 out.n3708 0.001
R85921 out.n3833 out.n3824 0.001
R85922 out.n3794 out.n3785 0.001
R85923 out.n3910 out.n3901 0.001
R85924 out.n3871 out.n3862 0.001
R85925 out.n907 out.n901 0.001
R85926 out.n3948 out.n3939 0.001
R85927 out.n8732 out.n8722 0.001
R85928 out.n8775 out.n8761 0.001
R85929 out.n8655 out.n8645 0.001
R85930 out.n8692 out.n8682 0.001
R85931 out.n8578 out.n8568 0.001
R85932 out.n8615 out.n8605 0.001
R85933 out.n8501 out.n8491 0.001
R85934 out.n8538 out.n8528 0.001
R85935 out.n8424 out.n8414 0.001
R85936 out.n8461 out.n8451 0.001
R85937 out.n8347 out.n8337 0.001
R85938 out.n8384 out.n8374 0.001
R85939 out.n8270 out.n8260 0.001
R85940 out.n8307 out.n8297 0.001
R85941 out.n8193 out.n8183 0.001
R85942 out.n8230 out.n8220 0.001
R85943 out.n8116 out.n8106 0.001
R85944 out.n8153 out.n8143 0.001
R85945 out.n8039 out.n8029 0.001
R85946 out.n8076 out.n8066 0.001
R85947 out.n7962 out.n7952 0.001
R85948 out.n7999 out.n7989 0.001
R85949 out.n7885 out.n7875 0.001
R85950 out.n7922 out.n7912 0.001
R85951 out.n6767 out.n6198 0.001
R85952 out.n7845 out.n7835 0.001
R85953 out.n3984 out.n3976 0.001
R85954 out.n6767 out.n6203 0.001
R85955 out.n7845 out.n7837 0.001
R85956 out.n7885 out.n7877 0.001
R85957 out.n7922 out.n7914 0.001
R85958 out.n7962 out.n7954 0.001
R85959 out.n7999 out.n7991 0.001
R85960 out.n8039 out.n8031 0.001
R85961 out.n8076 out.n8068 0.001
R85962 out.n8116 out.n8108 0.001
R85963 out.n8153 out.n8145 0.001
R85964 out.n8193 out.n8185 0.001
R85965 out.n8230 out.n8222 0.001
R85966 out.n8270 out.n8262 0.001
R85967 out.n8307 out.n8299 0.001
R85968 out.n8347 out.n8339 0.001
R85969 out.n8384 out.n8376 0.001
R85970 out.n8424 out.n8416 0.001
R85971 out.n8461 out.n8453 0.001
R85972 out.n8501 out.n8493 0.001
R85973 out.n8538 out.n8530 0.001
R85974 out.n8578 out.n8570 0.001
R85975 out.n8615 out.n8607 0.001
R85976 out.n8655 out.n8647 0.001
R85977 out.n8692 out.n8684 0.001
R85978 out.n8732 out.n8724 0.001
R85979 out.n8775 out.n8763 0.001
R85980 out.n907 out.n903 0.001
R85981 out.n3948 out.n3940 0.001
R85982 out.n3910 out.n3902 0.001
R85983 out.n3871 out.n3863 0.001
R85984 out.n3833 out.n3825 0.001
R85985 out.n3794 out.n3786 0.001
R85986 out.n3756 out.n3748 0.001
R85987 out.n3717 out.n3709 0.001
R85988 out.n3679 out.n3671 0.001
R85989 out.n3640 out.n3632 0.001
R85990 out.n3602 out.n3594 0.001
R85991 out.n3563 out.n3555 0.001
R85992 out.n3525 out.n3517 0.001
R85993 out.n3486 out.n3478 0.001
R85994 out.n3448 out.n3440 0.001
R85995 out.n3409 out.n3401 0.001
R85996 out.n3371 out.n3363 0.001
R85997 out.n3332 out.n3324 0.001
R85998 out.n3294 out.n3286 0.001
R85999 out.n3238 out.n3225 0.001
R86000 out.n3223 out.n3222 0.001
R86001 out.n3121 out.n3100 0.001
R86002 out.n3057 out.n3049 0.001
R86003 out.n2996 out.n2985 0.001
R86004 out.n2180 out.n1857 0.001
R86005 out.n3984 out.n3981 0.001
R86006 out.n15426 out.n15414 0.001
R86007 out.n12401 out.n12400 0.001
R86008 out.n9540 out.n9524 0.001
R86009 out.n9423 out.n9409 0.001
R86010 out.n9576 out.n9560 0.001
R86011 out.n9390 out.n9377 0.001
R86012 out.n9612 out.n9596 0.001
R86013 out.n9356 out.n9343 0.001
R86014 out.n9651 out.n9635 0.001
R86015 out.n9322 out.n9309 0.001
R86016 out.n9707 out.n9691 0.001
R86017 out.n9289 out.n9276 0.001
R86018 out.n9743 out.n9727 0.001
R86019 out.n9255 out.n9242 0.001
R86020 out.n9779 out.n9763 0.001
R86021 out.n9221 out.n9208 0.001
R86022 out.n9815 out.n9799 0.001
R86023 out.n9187 out.n9174 0.001
R86024 out.n9851 out.n9835 0.001
R86025 out.n9153 out.n9140 0.001
R86026 out.n9890 out.n9874 0.001
R86027 out.n9119 out.n9106 0.001
R86028 out.n9958 out.n9940 0.001
R86029 out.n9922 out.n9909 0.001
R86030 out.n9994 out.n9978 0.001
R86031 out.n9084 out.n9073 0.001
R86032 out.n9052 out.n9040 0.001
R86033 out.n9052 out.n9039 0.001
R86034 out.n16349 out.n16333 0.001
R86035 out.n16318 out.n16305 0.001
R86036 out.n16417 out.n16399 0.001
R86037 out.n16384 out.n16371 0.001
R86038 out.n16483 out.n16465 0.001
R86039 out.n16450 out.n16439 0.001
R86040 out.n16547 out.n16531 0.001
R86041 out.n16516 out.n16505 0.001
R86042 out.n16613 out.n16599 0.001
R86043 out.n16584 out.n16569 0.001
R86044 out.n16679 out.n16663 0.001
R86045 out.n16648 out.n16635 0.001
R86046 out.n16745 out.n16729 0.001
R86047 out.n16714 out.n16701 0.001
R86048 out.n16811 out.n16797 0.001
R86049 out.n16782 out.n16767 0.001
R86050 out.n16877 out.n16863 0.001
R86051 out.n16848 out.n16833 0.001
R86052 out.n16943 out.n16927 0.001
R86053 out.n16912 out.n16899 0.001
R86054 out.n17009 out.n16995 0.001
R86055 out.n16980 out.n16965 0.001
R86056 out.n17075 out.n17059 0.001
R86057 out.n17044 out.n17031 0.001
R86058 out.n17142 out.n17123 0.001
R86059 out.n17110 out.n17097 0.001
R86060 out.n17185 out.n17175 0.001
R86061 out.n9423 out.n9414 0.001
R86062 out.n9423 out.n9416 0.001
R86063 out.n9390 out.n9382 0.001
R86064 out.n9390 out.n9384 0.001
R86065 out.n9540 out.n9529 0.001
R86066 out.n9540 out.n9531 0.001
R86067 out.n9356 out.n9348 0.001
R86068 out.n9356 out.n9350 0.001
R86069 out.n9576 out.n9565 0.001
R86070 out.n9576 out.n9567 0.001
R86071 out.n9322 out.n9314 0.001
R86072 out.n9322 out.n9316 0.001
R86073 out.n9612 out.n9601 0.001
R86074 out.n9612 out.n9603 0.001
R86075 out.n9289 out.n9281 0.001
R86076 out.n9289 out.n9283 0.001
R86077 out.n9651 out.n9640 0.001
R86078 out.n9651 out.n9642 0.001
R86079 out.n9255 out.n9247 0.001
R86080 out.n9255 out.n9249 0.001
R86081 out.n9707 out.n9696 0.001
R86082 out.n9707 out.n9698 0.001
R86083 out.n9221 out.n9213 0.001
R86084 out.n9221 out.n9215 0.001
R86085 out.n9743 out.n9732 0.001
R86086 out.n9743 out.n9734 0.001
R86087 out.n9187 out.n9179 0.001
R86088 out.n9187 out.n9181 0.001
R86089 out.n9779 out.n9768 0.001
R86090 out.n9779 out.n9770 0.001
R86091 out.n9153 out.n9145 0.001
R86092 out.n9153 out.n9147 0.001
R86093 out.n9815 out.n9804 0.001
R86094 out.n9815 out.n9806 0.001
R86095 out.n9119 out.n9111 0.001
R86096 out.n9119 out.n9113 0.001
R86097 out.n9851 out.n9840 0.001
R86098 out.n9851 out.n9842 0.001
R86099 out.n9922 out.n9914 0.001
R86100 out.n9922 out.n9916 0.001
R86101 out.n9890 out.n9879 0.001
R86102 out.n9890 out.n9881 0.001
R86103 out.n9084 out.n9076 0.001
R86104 out.n9084 out.n9078 0.001
R86105 out.n9958 out.n9947 0.001
R86106 out.n9958 out.n9949 0.001
R86107 out.n9052 out.n9047 0.001
R86108 out.n9994 out.n9983 0.001
R86109 out.n9994 out.n9985 0.001
R86110 out.n16318 out.n16310 0.001
R86111 out.n16318 out.n16312 0.001
R86112 out.n16285 out.n16270 0.001
R86113 out.n16384 out.n16376 0.001
R86114 out.n16384 out.n16378 0.001
R86115 out.n16349 out.n16338 0.001
R86116 out.n16349 out.n16340 0.001
R86117 out.n16450 out.n16442 0.001
R86118 out.n16450 out.n16444 0.001
R86119 out.n16417 out.n16406 0.001
R86120 out.n16417 out.n16408 0.001
R86121 out.n16516 out.n16508 0.001
R86122 out.n16516 out.n16510 0.001
R86123 out.n16483 out.n16472 0.001
R86124 out.n16483 out.n16474 0.001
R86125 out.n16584 out.n16576 0.001
R86126 out.n16584 out.n16578 0.001
R86127 out.n16547 out.n16536 0.001
R86128 out.n16547 out.n16538 0.001
R86129 out.n16648 out.n16640 0.001
R86130 out.n16648 out.n16642 0.001
R86131 out.n16613 out.n16602 0.001
R86132 out.n16613 out.n16604 0.001
R86133 out.n16714 out.n16706 0.001
R86134 out.n16714 out.n16708 0.001
R86135 out.n16679 out.n16668 0.001
R86136 out.n16679 out.n16670 0.001
R86137 out.n16782 out.n16774 0.001
R86138 out.n16782 out.n16776 0.001
R86139 out.n16745 out.n16734 0.001
R86140 out.n16745 out.n16736 0.001
R86141 out.n16848 out.n16840 0.001
R86142 out.n16848 out.n16842 0.001
R86143 out.n16811 out.n16800 0.001
R86144 out.n16811 out.n16802 0.001
R86145 out.n16912 out.n16904 0.001
R86146 out.n16912 out.n16906 0.001
R86147 out.n16877 out.n16866 0.001
R86148 out.n16877 out.n16868 0.001
R86149 out.n16980 out.n16972 0.001
R86150 out.n16980 out.n16974 0.001
R86151 out.n16943 out.n16932 0.001
R86152 out.n16943 out.n16934 0.001
R86153 out.n17044 out.n17036 0.001
R86154 out.n17044 out.n17038 0.001
R86155 out.n17009 out.n16998 0.001
R86156 out.n17009 out.n17000 0.001
R86157 out.n17110 out.n17102 0.001
R86158 out.n17110 out.n17104 0.001
R86159 out.n17075 out.n17064 0.001
R86160 out.n17075 out.n17066 0.001
R86161 out.n17185 out.n17170 0.001
R86162 out.n17142 out.n17130 0.001
R86163 out.n17142 out.n17132 0.001
R86164 out.n9540 out.n9521 0.001
R86165 out.n9423 out.n9406 0.001
R86166 out.n9576 out.n9557 0.001
R86167 out.n9390 out.n9374 0.001
R86168 out.n9612 out.n9593 0.001
R86169 out.n9356 out.n9340 0.001
R86170 out.n9651 out.n9632 0.001
R86171 out.n9322 out.n9306 0.001
R86172 out.n9707 out.n9688 0.001
R86173 out.n9289 out.n9273 0.001
R86174 out.n9743 out.n9724 0.001
R86175 out.n9255 out.n9239 0.001
R86176 out.n9779 out.n9760 0.001
R86177 out.n9221 out.n9205 0.001
R86178 out.n9815 out.n9796 0.001
R86179 out.n9187 out.n9171 0.001
R86180 out.n9851 out.n9832 0.001
R86181 out.n9153 out.n9137 0.001
R86182 out.n9890 out.n9871 0.001
R86183 out.n9119 out.n9103 0.001
R86184 out.n9958 out.n9937 0.001
R86185 out.n9922 out.n9906 0.001
R86186 out.n9994 out.n9975 0.001
R86187 out.n9084 out.n9070 0.001
R86188 out.n9052 out.n9037 0.001
R86189 out.n9052 out.n9035 0.001
R86190 out.n16349 out.n16330 0.001
R86191 out.n16318 out.n16302 0.001
R86192 out.n16417 out.n16396 0.001
R86193 out.n16384 out.n16368 0.001
R86194 out.n16483 out.n16462 0.001
R86195 out.n16450 out.n16436 0.001
R86196 out.n16547 out.n16528 0.001
R86197 out.n16516 out.n16502 0.001
R86198 out.n16613 out.n16596 0.001
R86199 out.n16584 out.n16566 0.001
R86200 out.n16679 out.n16660 0.001
R86201 out.n16648 out.n16632 0.001
R86202 out.n16745 out.n16726 0.001
R86203 out.n16714 out.n16698 0.001
R86204 out.n16811 out.n16794 0.001
R86205 out.n16782 out.n16764 0.001
R86206 out.n16877 out.n16860 0.001
R86207 out.n16848 out.n16830 0.001
R86208 out.n16943 out.n16924 0.001
R86209 out.n16912 out.n16896 0.001
R86210 out.n17009 out.n16992 0.001
R86211 out.n16980 out.n16962 0.001
R86212 out.n17075 out.n17056 0.001
R86213 out.n17044 out.n17028 0.001
R86214 out.n17142 out.n17120 0.001
R86215 out.n17110 out.n17094 0.001
R86216 out.n17142 out.n17121 0.001
R86217 out.n17110 out.n17095 0.001
R86218 out.n17075 out.n17057 0.001
R86219 out.n17044 out.n17029 0.001
R86220 out.n17009 out.n16993 0.001
R86221 out.n16980 out.n16963 0.001
R86222 out.n16943 out.n16925 0.001
R86223 out.n16912 out.n16897 0.001
R86224 out.n16877 out.n16861 0.001
R86225 out.n16848 out.n16831 0.001
R86226 out.n16811 out.n16795 0.001
R86227 out.n16782 out.n16765 0.001
R86228 out.n16745 out.n16727 0.001
R86229 out.n16714 out.n16699 0.001
R86230 out.n16679 out.n16661 0.001
R86231 out.n16648 out.n16633 0.001
R86232 out.n16613 out.n16597 0.001
R86233 out.n16584 out.n16567 0.001
R86234 out.n16547 out.n16529 0.001
R86235 out.n16516 out.n16503 0.001
R86236 out.n16483 out.n16463 0.001
R86237 out.n16450 out.n16437 0.001
R86238 out.n16417 out.n16397 0.001
R86239 out.n16384 out.n16369 0.001
R86240 out.n16349 out.n16331 0.001
R86241 out.n16318 out.n16303 0.001
R86242 out.n16285 out.n10031 0.001
R86243 out.n9052 out.n9036 0.001
R86244 out.n9994 out.n9976 0.001
R86245 out.n9084 out.n9071 0.001
R86246 out.n9958 out.n9938 0.001
R86247 out.n9922 out.n9907 0.001
R86248 out.n9890 out.n9872 0.001
R86249 out.n9119 out.n9104 0.001
R86250 out.n9851 out.n9833 0.001
R86251 out.n9153 out.n9138 0.001
R86252 out.n9815 out.n9797 0.001
R86253 out.n9187 out.n9172 0.001
R86254 out.n9779 out.n9761 0.001
R86255 out.n9221 out.n9206 0.001
R86256 out.n9743 out.n9725 0.001
R86257 out.n9255 out.n9240 0.001
R86258 out.n9707 out.n9689 0.001
R86259 out.n9289 out.n9274 0.001
R86260 out.n9651 out.n9633 0.001
R86261 out.n9322 out.n9307 0.001
R86262 out.n9612 out.n9594 0.001
R86263 out.n9356 out.n9341 0.001
R86264 out.n9576 out.n9558 0.001
R86265 out.n9390 out.n9375 0.001
R86266 out.n9540 out.n9522 0.001
R86267 out.n9423 out.n9407 0.001
R86268 out.n9506 out.n9490 0.001
R86269 out.n9540 out.n9532 0.001
R86270 out.n9540 out.n9535 0.001
R86271 out.n9423 out.n9417 0.001
R86272 out.n9423 out.n9419 0.001
R86273 out.n9576 out.n9568 0.001
R86274 out.n9576 out.n9571 0.001
R86275 out.n9390 out.n9385 0.001
R86276 out.n9390 out.n9387 0.001
R86277 out.n9612 out.n9604 0.001
R86278 out.n9612 out.n9607 0.001
R86279 out.n9356 out.n9351 0.001
R86280 out.n9356 out.n9353 0.001
R86281 out.n9651 out.n9643 0.001
R86282 out.n9651 out.n9646 0.001
R86283 out.n9322 out.n9317 0.001
R86284 out.n9322 out.n9319 0.001
R86285 out.n9707 out.n9699 0.001
R86286 out.n9707 out.n9702 0.001
R86287 out.n9289 out.n9284 0.001
R86288 out.n9289 out.n9286 0.001
R86289 out.n9743 out.n9735 0.001
R86290 out.n9743 out.n9738 0.001
R86291 out.n9255 out.n9250 0.001
R86292 out.n9255 out.n9252 0.001
R86293 out.n9779 out.n9771 0.001
R86294 out.n9779 out.n9774 0.001
R86295 out.n9221 out.n9216 0.001
R86296 out.n9221 out.n9218 0.001
R86297 out.n9815 out.n9807 0.001
R86298 out.n9815 out.n9810 0.001
R86299 out.n9187 out.n9182 0.001
R86300 out.n9187 out.n9184 0.001
R86301 out.n9851 out.n9843 0.001
R86302 out.n9851 out.n9846 0.001
R86303 out.n9153 out.n9148 0.001
R86304 out.n9153 out.n9150 0.001
R86305 out.n9890 out.n9882 0.001
R86306 out.n9890 out.n9885 0.001
R86307 out.n9119 out.n9114 0.001
R86308 out.n9119 out.n9116 0.001
R86309 out.n9958 out.n9950 0.001
R86310 out.n9958 out.n9953 0.001
R86311 out.n9922 out.n9917 0.001
R86312 out.n9922 out.n9919 0.001
R86313 out.n9994 out.n9986 0.001
R86314 out.n9994 out.n9989 0.001
R86315 out.n9084 out.n9079 0.001
R86316 out.n9084 out.n9081 0.001
R86317 out.n16285 out.n16275 0.001
R86318 out.n9052 out.n9049 0.001
R86319 out.n16349 out.n16341 0.001
R86320 out.n16349 out.n16344 0.001
R86321 out.n16318 out.n16313 0.001
R86322 out.n16318 out.n16315 0.001
R86323 out.n16417 out.n16409 0.001
R86324 out.n16417 out.n16412 0.001
R86325 out.n16384 out.n16379 0.001
R86326 out.n16384 out.n16381 0.001
R86327 out.n16483 out.n16475 0.001
R86328 out.n16483 out.n16478 0.001
R86329 out.n16450 out.n16445 0.001
R86330 out.n16450 out.n16447 0.001
R86331 out.n16547 out.n16539 0.001
R86332 out.n16547 out.n16542 0.001
R86333 out.n16516 out.n16511 0.001
R86334 out.n16516 out.n16513 0.001
R86335 out.n16613 out.n16605 0.001
R86336 out.n16613 out.n16608 0.001
R86337 out.n16584 out.n16579 0.001
R86338 out.n16584 out.n16581 0.001
R86339 out.n16679 out.n16671 0.001
R86340 out.n16679 out.n16674 0.001
R86341 out.n16648 out.n16643 0.001
R86342 out.n16648 out.n16645 0.001
R86343 out.n16745 out.n16737 0.001
R86344 out.n16745 out.n16740 0.001
R86345 out.n16714 out.n16709 0.001
R86346 out.n16714 out.n16711 0.001
R86347 out.n16811 out.n16803 0.001
R86348 out.n16811 out.n16806 0.001
R86349 out.n16782 out.n16777 0.001
R86350 out.n16782 out.n16779 0.001
R86351 out.n16877 out.n16869 0.001
R86352 out.n16877 out.n16872 0.001
R86353 out.n16848 out.n16843 0.001
R86354 out.n16848 out.n16845 0.001
R86355 out.n16943 out.n16935 0.001
R86356 out.n16943 out.n16938 0.001
R86357 out.n16912 out.n16907 0.001
R86358 out.n16912 out.n16909 0.001
R86359 out.n17009 out.n17001 0.001
R86360 out.n17009 out.n17004 0.001
R86361 out.n16980 out.n16975 0.001
R86362 out.n16980 out.n16977 0.001
R86363 out.n17075 out.n17067 0.001
R86364 out.n17075 out.n17070 0.001
R86365 out.n17044 out.n17039 0.001
R86366 out.n17044 out.n17041 0.001
R86367 out.n17142 out.n17133 0.001
R86368 out.n17142 out.n17136 0.001
R86369 out.n17110 out.n17105 0.001
R86370 out.n17110 out.n17107 0.001
R86371 out.n17185 out.n17166 0.001
R86372 out.n17185 out.n17168 0.001
R86373 out.n17185 out.n17155 0.001
R86374 out.n17142 out.n17118 0.001
R86375 out.n17110 out.n17085 0.001
R86376 out.n17075 out.n17054 0.001
R86377 out.n17044 out.n17019 0.001
R86378 out.n17009 out.n16990 0.001
R86379 out.n16980 out.n16953 0.001
R86380 out.n16943 out.n16922 0.001
R86381 out.n16912 out.n16887 0.001
R86382 out.n16877 out.n16858 0.001
R86383 out.n16848 out.n16821 0.001
R86384 out.n16811 out.n16792 0.001
R86385 out.n16782 out.n16755 0.001
R86386 out.n16745 out.n16724 0.001
R86387 out.n16714 out.n16689 0.001
R86388 out.n16679 out.n16658 0.001
R86389 out.n16648 out.n16623 0.001
R86390 out.n16613 out.n16594 0.001
R86391 out.n16584 out.n16557 0.001
R86392 out.n16547 out.n16526 0.001
R86393 out.n16516 out.n16493 0.001
R86394 out.n16483 out.n16460 0.001
R86395 out.n16450 out.n16427 0.001
R86396 out.n16417 out.n16394 0.001
R86397 out.n16384 out.n16359 0.001
R86398 out.n16349 out.n16328 0.001
R86399 out.n16318 out.n16293 0.001
R86400 out.n16285 out.n10026 0.001
R86401 out.n9052 out.n9025 0.001
R86402 out.n9994 out.n9973 0.001
R86403 out.n9084 out.n9061 0.001
R86404 out.n9958 out.n9935 0.001
R86405 out.n9922 out.n9897 0.001
R86406 out.n9890 out.n9869 0.001
R86407 out.n9119 out.n9094 0.001
R86408 out.n9851 out.n9830 0.001
R86409 out.n9153 out.n9128 0.001
R86410 out.n9815 out.n9794 0.001
R86411 out.n9187 out.n9162 0.001
R86412 out.n9779 out.n9758 0.001
R86413 out.n9221 out.n9196 0.001
R86414 out.n9743 out.n9722 0.001
R86415 out.n9255 out.n9230 0.001
R86416 out.n9707 out.n9686 0.001
R86417 out.n9289 out.n9264 0.001
R86418 out.n9651 out.n9630 0.001
R86419 out.n9322 out.n9297 0.001
R86420 out.n9612 out.n9591 0.001
R86421 out.n9356 out.n9331 0.001
R86422 out.n9576 out.n9555 0.001
R86423 out.n9390 out.n9365 0.001
R86424 out.n9540 out.n9519 0.001
R86425 out.n17110 out.n17086 0.001
R86426 out.n17044 out.n17020 0.001
R86427 out.n16980 out.n16954 0.001
R86428 out.n16912 out.n16888 0.001
R86429 out.n16848 out.n16822 0.001
R86430 out.n16782 out.n16756 0.001
R86431 out.n16714 out.n16690 0.001
R86432 out.n16648 out.n16624 0.001
R86433 out.n16584 out.n16558 0.001
R86434 out.n16516 out.n16494 0.001
R86435 out.n16450 out.n16428 0.001
R86436 out.n16384 out.n16360 0.001
R86437 out.n16318 out.n16294 0.001
R86438 out.n9052 out.n9026 0.001
R86439 out.n9084 out.n9062 0.001
R86440 out.n9922 out.n9898 0.001
R86441 out.n9119 out.n9095 0.001
R86442 out.n9153 out.n9129 0.001
R86443 out.n9187 out.n9163 0.001
R86444 out.n9221 out.n9197 0.001
R86445 out.n9255 out.n9231 0.001
R86446 out.n9289 out.n9265 0.001
R86447 out.n9322 out.n9298 0.001
R86448 out.n9356 out.n9332 0.001
R86449 out.n9390 out.n9366 0.001
R86450 out.n9540 out.n9516 0.001
R86451 out.n17142 out.n17115 0.001
R86452 out.n17075 out.n17051 0.001
R86453 out.n17009 out.n16987 0.001
R86454 out.n16943 out.n16919 0.001
R86455 out.n16877 out.n16855 0.001
R86456 out.n16811 out.n16789 0.001
R86457 out.n16745 out.n16721 0.001
R86458 out.n16679 out.n16655 0.001
R86459 out.n16613 out.n16591 0.001
R86460 out.n16547 out.n16523 0.001
R86461 out.n16483 out.n16457 0.001
R86462 out.n16417 out.n16391 0.001
R86463 out.n16349 out.n16325 0.001
R86464 out.n16285 out.n10021 0.001
R86465 out.n9052 out.n9029 0.001
R86466 out.n9994 out.n9970 0.001
R86467 out.n9958 out.n9932 0.001
R86468 out.n9890 out.n9866 0.001
R86469 out.n9851 out.n9827 0.001
R86470 out.n9815 out.n9791 0.001
R86471 out.n9779 out.n9755 0.001
R86472 out.n9743 out.n9719 0.001
R86473 out.n9707 out.n9683 0.001
R86474 out.n9651 out.n9627 0.001
R86475 out.n9612 out.n9588 0.001
R86476 out.n9576 out.n9552 0.001
R86477 out.n9540 out.n9514 0.001
R86478 out.n9506 out.n9487 0.001
R86479 out.n17185 out.n17159 0.001
R86480 out.n17142 out.n17114 0.001
R86481 out.n17142 out.n17113 0.001
R86482 out.n17110 out.n17090 0.001
R86483 out.n17110 out.n17088 0.001
R86484 out.n17075 out.n17050 0.001
R86485 out.n17075 out.n17049 0.001
R86486 out.n17044 out.n17024 0.001
R86487 out.n17044 out.n17022 0.001
R86488 out.n17009 out.n16986 0.001
R86489 out.n17009 out.n16985 0.001
R86490 out.n16980 out.n16958 0.001
R86491 out.n16980 out.n16956 0.001
R86492 out.n16943 out.n16918 0.001
R86493 out.n16943 out.n16917 0.001
R86494 out.n16912 out.n16892 0.001
R86495 out.n16912 out.n16890 0.001
R86496 out.n16877 out.n16854 0.001
R86497 out.n16877 out.n16853 0.001
R86498 out.n16848 out.n16826 0.001
R86499 out.n16848 out.n16824 0.001
R86500 out.n16811 out.n16788 0.001
R86501 out.n16811 out.n16787 0.001
R86502 out.n16782 out.n16760 0.001
R86503 out.n16782 out.n16758 0.001
R86504 out.n16745 out.n16720 0.001
R86505 out.n16745 out.n16719 0.001
R86506 out.n16714 out.n16694 0.001
R86507 out.n16714 out.n16692 0.001
R86508 out.n16679 out.n16654 0.001
R86509 out.n16679 out.n16653 0.001
R86510 out.n16648 out.n16628 0.001
R86511 out.n16648 out.n16626 0.001
R86512 out.n16613 out.n16590 0.001
R86513 out.n16613 out.n16589 0.001
R86514 out.n16584 out.n16562 0.001
R86515 out.n16584 out.n16560 0.001
R86516 out.n16547 out.n16522 0.001
R86517 out.n16547 out.n16521 0.001
R86518 out.n16516 out.n16498 0.001
R86519 out.n16516 out.n16496 0.001
R86520 out.n16483 out.n16456 0.001
R86521 out.n16483 out.n16455 0.001
R86522 out.n16450 out.n16432 0.001
R86523 out.n16450 out.n16430 0.001
R86524 out.n16417 out.n16390 0.001
R86525 out.n16417 out.n16389 0.001
R86526 out.n16384 out.n16364 0.001
R86527 out.n16384 out.n16362 0.001
R86528 out.n16349 out.n16324 0.001
R86529 out.n16349 out.n16323 0.001
R86530 out.n16318 out.n16298 0.001
R86531 out.n16318 out.n16296 0.001
R86532 out.n16285 out.n10010 0.001
R86533 out.n9052 out.n9028 0.001
R86534 out.n9994 out.n9969 0.001
R86535 out.n9994 out.n9968 0.001
R86536 out.n9084 out.n9066 0.001
R86537 out.n9084 out.n9064 0.001
R86538 out.n9958 out.n9931 0.001
R86539 out.n9958 out.n9930 0.001
R86540 out.n9922 out.n9902 0.001
R86541 out.n9922 out.n9900 0.001
R86542 out.n9890 out.n9865 0.001
R86543 out.n9890 out.n9864 0.001
R86544 out.n9119 out.n9099 0.001
R86545 out.n9119 out.n9097 0.001
R86546 out.n9851 out.n9826 0.001
R86547 out.n9851 out.n9825 0.001
R86548 out.n9153 out.n9133 0.001
R86549 out.n9153 out.n9131 0.001
R86550 out.n9815 out.n9790 0.001
R86551 out.n9815 out.n9789 0.001
R86552 out.n9187 out.n9167 0.001
R86553 out.n9187 out.n9165 0.001
R86554 out.n9779 out.n9754 0.001
R86555 out.n9779 out.n9753 0.001
R86556 out.n9221 out.n9201 0.001
R86557 out.n9221 out.n9199 0.001
R86558 out.n9743 out.n9718 0.001
R86559 out.n9743 out.n9717 0.001
R86560 out.n9255 out.n9235 0.001
R86561 out.n9255 out.n9233 0.001
R86562 out.n9707 out.n9682 0.001
R86563 out.n9707 out.n9681 0.001
R86564 out.n9289 out.n9269 0.001
R86565 out.n9289 out.n9267 0.001
R86566 out.n9651 out.n9626 0.001
R86567 out.n9651 out.n9625 0.001
R86568 out.n9322 out.n9302 0.001
R86569 out.n9322 out.n9300 0.001
R86570 out.n9612 out.n9587 0.001
R86571 out.n9612 out.n9586 0.001
R86572 out.n9356 out.n9336 0.001
R86573 out.n9356 out.n9334 0.001
R86574 out.n9576 out.n9551 0.001
R86575 out.n9576 out.n9550 0.001
R86576 out.n9390 out.n9370 0.001
R86577 out.n9390 out.n9368 0.001
R86578 out.n9540 out.n9513 0.001
R86579 out.n9423 out.n9404 0.001
R86580 out.n9423 out.n9402 0.001
R86581 out.n9423 out.n9401 0.001
R86582 out.n9423 out.n9397 0.001
R86583 out.n17185 out.n17164 0.001
R86584 out.n17142 out.n17117 0.001
R86585 out.n17110 out.n17092 0.001
R86586 out.n17075 out.n17053 0.001
R86587 out.n17044 out.n17026 0.001
R86588 out.n17009 out.n16989 0.001
R86589 out.n16980 out.n16960 0.001
R86590 out.n16943 out.n16921 0.001
R86591 out.n16912 out.n16894 0.001
R86592 out.n16877 out.n16857 0.001
R86593 out.n16848 out.n16828 0.001
R86594 out.n16811 out.n16791 0.001
R86595 out.n16782 out.n16762 0.001
R86596 out.n16745 out.n16723 0.001
R86597 out.n16714 out.n16696 0.001
R86598 out.n16679 out.n16657 0.001
R86599 out.n16648 out.n16630 0.001
R86600 out.n16613 out.n16593 0.001
R86601 out.n16584 out.n16564 0.001
R86602 out.n16547 out.n16525 0.001
R86603 out.n16516 out.n16500 0.001
R86604 out.n16483 out.n16459 0.001
R86605 out.n16450 out.n16434 0.001
R86606 out.n16417 out.n16393 0.001
R86607 out.n16384 out.n16366 0.001
R86608 out.n16349 out.n16327 0.001
R86609 out.n16318 out.n16300 0.001
R86610 out.n9052 out.n9031 0.001
R86611 out.n9052 out.n9033 0.001
R86612 out.n9994 out.n9972 0.001
R86613 out.n9084 out.n9068 0.001
R86614 out.n9958 out.n9934 0.001
R86615 out.n9922 out.n9904 0.001
R86616 out.n9890 out.n9868 0.001
R86617 out.n9119 out.n9101 0.001
R86618 out.n9851 out.n9829 0.001
R86619 out.n9153 out.n9135 0.001
R86620 out.n9815 out.n9793 0.001
R86621 out.n9187 out.n9169 0.001
R86622 out.n9779 out.n9757 0.001
R86623 out.n9221 out.n9203 0.001
R86624 out.n9743 out.n9721 0.001
R86625 out.n9255 out.n9237 0.001
R86626 out.n9707 out.n9685 0.001
R86627 out.n9289 out.n9271 0.001
R86628 out.n9651 out.n9629 0.001
R86629 out.n9322 out.n9304 0.001
R86630 out.n9612 out.n9590 0.001
R86631 out.n9356 out.n9338 0.001
R86632 out.n9576 out.n9554 0.001
R86633 out.n9390 out.n9372 0.001
R86634 out.n9540 out.n9518 0.001
R86635 out.n9506 out.n9477 0.001
R86636 out.n9506 out.n9478 0.001
R86637 out.n9540 out.n9536 0.001
R86638 out.n9576 out.n9572 0.001
R86639 out.n9390 out.n9389 0.001
R86640 out.n9612 out.n9608 0.001
R86641 out.n9356 out.n9355 0.001
R86642 out.n9651 out.n9647 0.001
R86643 out.n9322 out.n9321 0.001
R86644 out.n9707 out.n9703 0.001
R86645 out.n9289 out.n9288 0.001
R86646 out.n9743 out.n9739 0.001
R86647 out.n9255 out.n9254 0.001
R86648 out.n9779 out.n9775 0.001
R86649 out.n9221 out.n9220 0.001
R86650 out.n9815 out.n9811 0.001
R86651 out.n9187 out.n9186 0.001
R86652 out.n9851 out.n9847 0.001
R86653 out.n9153 out.n9152 0.001
R86654 out.n9890 out.n9886 0.001
R86655 out.n9119 out.n9118 0.001
R86656 out.n9958 out.n9954 0.001
R86657 out.n9922 out.n9921 0.001
R86658 out.n9994 out.n9990 0.001
R86659 out.n9084 out.n9083 0.001
R86660 out.n16285 out.n16280 0.001
R86661 out.n9052 out.n9051 0.001
R86662 out.n16349 out.n16345 0.001
R86663 out.n16318 out.n16317 0.001
R86664 out.n16417 out.n16413 0.001
R86665 out.n16384 out.n16383 0.001
R86666 out.n16483 out.n16479 0.001
R86667 out.n16450 out.n16449 0.001
R86668 out.n16547 out.n16543 0.001
R86669 out.n16516 out.n16515 0.001
R86670 out.n16613 out.n16609 0.001
R86671 out.n16584 out.n16583 0.001
R86672 out.n16679 out.n16675 0.001
R86673 out.n16648 out.n16647 0.001
R86674 out.n16745 out.n16741 0.001
R86675 out.n16714 out.n16713 0.001
R86676 out.n16811 out.n16807 0.001
R86677 out.n16782 out.n16781 0.001
R86678 out.n16877 out.n16873 0.001
R86679 out.n16848 out.n16847 0.001
R86680 out.n16943 out.n16939 0.001
R86681 out.n16912 out.n16911 0.001
R86682 out.n17009 out.n17005 0.001
R86683 out.n16980 out.n16979 0.001
R86684 out.n17075 out.n17071 0.001
R86685 out.n17044 out.n17043 0.001
R86686 out.n17142 out.n17138 0.001
R86687 out.n17110 out.n17109 0.001
R86688 out.n17142 out.n17140 0.001
R86689 out.n17110 out.n17083 0.001
R86690 out.n17075 out.n17073 0.001
R86691 out.n17044 out.n17017 0.001
R86692 out.n17009 out.n17007 0.001
R86693 out.n16980 out.n16951 0.001
R86694 out.n16943 out.n16941 0.001
R86695 out.n16912 out.n16885 0.001
R86696 out.n16877 out.n16875 0.001
R86697 out.n16848 out.n16819 0.001
R86698 out.n16811 out.n16809 0.001
R86699 out.n16782 out.n16753 0.001
R86700 out.n16745 out.n16743 0.001
R86701 out.n16714 out.n16687 0.001
R86702 out.n16679 out.n16677 0.001
R86703 out.n16648 out.n16621 0.001
R86704 out.n16613 out.n16611 0.001
R86705 out.n16584 out.n16555 0.001
R86706 out.n16547 out.n16545 0.001
R86707 out.n16516 out.n16491 0.001
R86708 out.n16483 out.n16481 0.001
R86709 out.n16450 out.n16425 0.001
R86710 out.n16417 out.n16415 0.001
R86711 out.n16384 out.n16357 0.001
R86712 out.n16349 out.n16347 0.001
R86713 out.n16318 out.n16291 0.001
R86714 out.n9994 out.n9992 0.001
R86715 out.n9084 out.n9059 0.001
R86716 out.n9958 out.n9956 0.001
R86717 out.n9922 out.n9895 0.001
R86718 out.n9890 out.n9888 0.001
R86719 out.n9119 out.n9092 0.001
R86720 out.n9851 out.n9849 0.001
R86721 out.n9153 out.n9126 0.001
R86722 out.n9815 out.n9813 0.001
R86723 out.n9187 out.n9160 0.001
R86724 out.n9779 out.n9777 0.001
R86725 out.n9221 out.n9194 0.001
R86726 out.n9743 out.n9741 0.001
R86727 out.n9255 out.n9228 0.001
R86728 out.n9707 out.n9705 0.001
R86729 out.n9289 out.n9262 0.001
R86730 out.n9651 out.n9649 0.001
R86731 out.n9322 out.n9295 0.001
R86732 out.n9612 out.n9610 0.001
R86733 out.n9356 out.n9329 0.001
R86734 out.n9576 out.n9574 0.001
R86735 out.n9390 out.n9363 0.001
R86736 out.n9540 out.n9538 0.001
R86737 out.n9423 out.n9398 0.001
R86738 out.n9423 out.n9421 0.001
R86739 out.n17185 out.n17184 0.001
R86740 out.n17110 out.n17082 0.001
R86741 out.n17075 out.n17047 0.001
R86742 out.n17044 out.n17016 0.001
R86743 out.n17009 out.n16983 0.001
R86744 out.n16980 out.n16950 0.001
R86745 out.n16943 out.n16915 0.001
R86746 out.n16912 out.n16884 0.001
R86747 out.n16877 out.n16851 0.001
R86748 out.n16848 out.n16818 0.001
R86749 out.n16811 out.n16785 0.001
R86750 out.n16782 out.n16752 0.001
R86751 out.n16745 out.n16717 0.001
R86752 out.n16714 out.n16686 0.001
R86753 out.n16679 out.n16651 0.001
R86754 out.n16648 out.n16620 0.001
R86755 out.n16613 out.n16587 0.001
R86756 out.n16584 out.n16554 0.001
R86757 out.n16547 out.n16519 0.001
R86758 out.n16516 out.n16490 0.001
R86759 out.n16483 out.n16453 0.001
R86760 out.n16450 out.n16424 0.001
R86761 out.n16417 out.n16387 0.001
R86762 out.n16384 out.n16356 0.001
R86763 out.n16349 out.n16321 0.001
R86764 out.n16318 out.n16290 0.001
R86765 out.n16285 out.n10003 0.001
R86766 out.n9052 out.n9023 0.001
R86767 out.n9994 out.n9966 0.001
R86768 out.n9084 out.n9058 0.001
R86769 out.n9958 out.n9928 0.001
R86770 out.n9922 out.n9894 0.001
R86771 out.n9890 out.n9862 0.001
R86772 out.n9119 out.n9091 0.001
R86773 out.n9851 out.n9823 0.001
R86774 out.n9153 out.n9125 0.001
R86775 out.n9815 out.n9787 0.001
R86776 out.n9187 out.n9159 0.001
R86777 out.n9779 out.n9751 0.001
R86778 out.n9221 out.n9193 0.001
R86779 out.n9743 out.n9715 0.001
R86780 out.n9255 out.n9227 0.001
R86781 out.n9707 out.n9679 0.001
R86782 out.n9289 out.n9261 0.001
R86783 out.n9651 out.n9623 0.001
R86784 out.n9322 out.n9294 0.001
R86785 out.n9612 out.n9584 0.001
R86786 out.n9356 out.n9328 0.001
R86787 out.n9576 out.n9548 0.001
R86788 out.n9390 out.n9362 0.001
R86789 out.n9540 out.n9512 0.001
R86790 out.n9423 out.n9395 0.001
R86791 out.n9506 out.n9471 0.001
R86792 out.n56 out.n40 0.001
R86793 out.n119 out.n107 0.001
R86794 out.n185 out.n171 0.001
R86795 out.n251 out.n238 0.001
R86796 out.n313 out.n299 0.001
R86797 out.n381 out.n368 0.001
R86798 out.n444 out.n431 0.001
R86799 out.n511 out.n496 0.001
R86800 out.n572 out.n558 0.001
R86801 out.n638 out.n624 0.001
R86802 out.n705 out.n690 0.001
R86803 out.n768 out.n750 0.001
R86804 out.n828 out.n813 0.001
R86805 out.n919 out.n891 0.001
R86806 out.n919 out.n889 0.001
R86807 out.n4026 out.n4012 0.001
R86808 out.n4092 out.n4078 0.001
R86809 out.n4155 out.n4139 0.001
R86810 out.n4219 out.n4205 0.001
R86811 out.n4282 out.n4270 0.001
R86812 out.n4349 out.n4335 0.001
R86813 out.n4414 out.n4400 0.001
R86814 out.n4478 out.n4465 0.001
R86815 out.n4541 out.n4527 0.001
R86816 out.n4609 out.n4594 0.001
R86817 out.n4673 out.n4659 0.001
R86818 out.n4737 out.n4723 0.001
R86819 out.n4800 out.n4785 0.001
R86820 out.n4800 out.n4794 0.001
R86821 out.n4763 out.n4755 0.001
R86822 out.n4737 out.n4731 0.001
R86823 out.n4699 out.n4692 0.001
R86824 out.n4673 out.n4667 0.001
R86825 out.n4637 out.n4630 0.001
R86826 out.n4609 out.n4603 0.001
R86827 out.n4570 out.n4562 0.001
R86828 out.n4541 out.n4536 0.001
R86829 out.n4506 out.n4496 0.001
R86830 out.n4478 out.n4472 0.001
R86831 out.n4441 out.n4435 0.001
R86832 out.n4414 out.n4407 0.001
R86833 out.n4378 out.n4370 0.001
R86834 out.n4349 out.n4344 0.001
R86835 out.n4313 out.n4303 0.001
R86836 out.n4282 out.n4276 0.001
R86837 out.n4247 out.n4240 0.001
R86838 out.n4219 out.n4213 0.001
R86839 out.n4183 out.n4177 0.001
R86840 out.n4155 out.n4148 0.001
R86841 out.n4120 out.n4113 0.001
R86842 out.n4092 out.n4086 0.001
R86843 out.n4054 out.n4047 0.001
R86844 out.n4026 out.n4020 0.001
R86845 out.n4942 out.n4935 0.001
R86846 out.n4942 out.n4928 0.001
R86847 out.n858 out.n848 0.001
R86848 out.n828 out.n821 0.001
R86849 out.n791 out.n784 0.001
R86850 out.n768 out.n760 0.001
R86851 out.n729 out.n723 0.001
R86852 out.n705 out.n699 0.001
R86853 out.n664 out.n656 0.001
R86854 out.n638 out.n632 0.001
R86855 out.n601 out.n593 0.001
R86856 out.n572 out.n566 0.001
R86857 out.n533 out.n525 0.001
R86858 out.n511 out.n505 0.001
R86859 out.n472 out.n464 0.001
R86860 out.n444 out.n438 0.001
R86861 out.n409 out.n402 0.001
R86862 out.n381 out.n375 0.001
R86863 out.n344 out.n337 0.001
R86864 out.n313 out.n307 0.001
R86865 out.n274 out.n266 0.001
R86866 out.n251 out.n246 0.001
R86867 out.n213 out.n205 0.001
R86868 out.n185 out.n180 0.001
R86869 out.n148 out.n140 0.001
R86870 out.n119 out.n114 0.001
R86871 out.n88 out.n80 0.001
R86872 out.n56 out.n51 0.001
R86873 out.n56 out.n43 0.001
R86874 out.n919 out.n915 0.001
R86875 out.n4835 out.n4817 0.001
R86876 out.n4800 out.n4795 0.001
R86877 out.n4763 out.n4757 0.001
R86878 out.n4763 out.n4750 0.001
R86879 out.n4737 out.n4732 0.001
R86880 out.n4699 out.n4693 0.001
R86881 out.n4699 out.n4686 0.001
R86882 out.n4673 out.n4668 0.001
R86883 out.n4637 out.n4631 0.001
R86884 out.n4637 out.n4624 0.001
R86885 out.n4609 out.n4604 0.001
R86886 out.n4570 out.n4563 0.001
R86887 out.n4570 out.n4556 0.001
R86888 out.n4541 out.n4537 0.001
R86889 out.n4506 out.n4498 0.001
R86890 out.n4506 out.n4491 0.001
R86891 out.n4478 out.n4473 0.001
R86892 out.n4441 out.n4436 0.001
R86893 out.n4441 out.n4428 0.001
R86894 out.n4414 out.n4409 0.001
R86895 out.n4378 out.n4371 0.001
R86896 out.n4378 out.n4364 0.001
R86897 out.n4349 out.n4345 0.001
R86898 out.n4313 out.n4305 0.001
R86899 out.n4313 out.n4296 0.001
R86900 out.n4282 out.n4277 0.001
R86901 out.n4247 out.n4241 0.001
R86902 out.n4247 out.n4234 0.001
R86903 out.n4219 out.n4214 0.001
R86904 out.n4183 out.n4178 0.001
R86905 out.n4183 out.n4171 0.001
R86906 out.n4155 out.n4150 0.001
R86907 out.n4120 out.n4114 0.001
R86908 out.n4120 out.n4108 0.001
R86909 out.n4092 out.n4087 0.001
R86910 out.n4054 out.n4048 0.001
R86911 out.n4054 out.n4041 0.001
R86912 out.n4026 out.n4021 0.001
R86913 out.n4942 out.n4936 0.001
R86914 out.n4942 out.n4926 0.001
R86915 out.n858 out.n850 0.001
R86916 out.n858 out.n842 0.001
R86917 out.n828 out.n822 0.001
R86918 out.n791 out.n785 0.001
R86919 out.n791 out.n779 0.001
R86920 out.n768 out.n762 0.001
R86921 out.n729 out.n724 0.001
R86922 out.n729 out.n719 0.001
R86923 out.n705 out.n701 0.001
R86924 out.n664 out.n657 0.001
R86925 out.n664 out.n651 0.001
R86926 out.n638 out.n633 0.001
R86927 out.n601 out.n594 0.001
R86928 out.n601 out.n586 0.001
R86929 out.n572 out.n567 0.001
R86930 out.n533 out.n526 0.001
R86931 out.n533 out.n521 0.001
R86932 out.n511 out.n507 0.001
R86933 out.n472 out.n465 0.001
R86934 out.n472 out.n457 0.001
R86935 out.n444 out.n439 0.001
R86936 out.n409 out.n403 0.001
R86937 out.n409 out.n395 0.001
R86938 out.n381 out.n376 0.001
R86939 out.n344 out.n338 0.001
R86940 out.n344 out.n329 0.001
R86941 out.n313 out.n308 0.001
R86942 out.n274 out.n268 0.001
R86943 out.n274 out.n262 0.001
R86944 out.n251 out.n247 0.001
R86945 out.n213 out.n206 0.001
R86946 out.n213 out.n199 0.001
R86947 out.n185 out.n181 0.001
R86948 out.n148 out.n141 0.001
R86949 out.n148 out.n134 0.001
R86950 out.n119 out.n115 0.001
R86951 out.n88 out.n82 0.001
R86952 out.n88 out.n73 0.001
R86953 out.n56 out.n52 0.001
R86954 out.n88 out.n71 0.001
R86955 out.n56 out.n36 0.001
R86956 out.n251 out.n236 0.001
R86957 out.n4942 out.n4939 0.001
R86958 out.n88 out.n85 0.001
R86959 out.n148 out.n145 0.001
R86960 out.n213 out.n210 0.001
R86961 out.n274 out.n271 0.001
R86962 out.n344 out.n341 0.001
R86963 out.n409 out.n406 0.001
R86964 out.n472 out.n469 0.001
R86965 out.n533 out.n530 0.001
R86966 out.n601 out.n598 0.001
R86967 out.n664 out.n661 0.001
R86968 out.n729 out.n726 0.001
R86969 out.n791 out.n788 0.001
R86970 out.n858 out.n855 0.001
R86971 out.n4054 out.n4051 0.001
R86972 out.n4120 out.n4117 0.001
R86973 out.n4183 out.n4180 0.001
R86974 out.n4247 out.n4244 0.001
R86975 out.n4313 out.n4310 0.001
R86976 out.n4378 out.n4375 0.001
R86977 out.n4441 out.n4438 0.001
R86978 out.n4506 out.n4503 0.001
R86979 out.n4570 out.n4567 0.001
R86980 out.n4637 out.n4634 0.001
R86981 out.n4699 out.n4696 0.001
R86982 out.n4763 out.n4760 0.001
R86983 out.n4835 out.n4833 0.001
R86984 out.n4800 out.n4783 0.001
R86985 out.n4800 out.n4799 0.001
R86986 out.n4763 out.n4748 0.001
R86987 out.n4763 out.n4762 0.001
R86988 out.n4737 out.n4720 0.001
R86989 out.n4737 out.n4736 0.001
R86990 out.n4699 out.n4683 0.001
R86991 out.n4699 out.n4698 0.001
R86992 out.n4673 out.n4656 0.001
R86993 out.n4673 out.n4672 0.001
R86994 out.n4637 out.n4621 0.001
R86995 out.n4637 out.n4636 0.001
R86996 out.n4609 out.n4591 0.001
R86997 out.n4609 out.n4608 0.001
R86998 out.n4570 out.n4553 0.001
R86999 out.n4570 out.n4569 0.001
R87000 out.n4541 out.n4525 0.001
R87001 out.n4541 out.n4540 0.001
R87002 out.n4506 out.n4489 0.001
R87003 out.n4506 out.n4505 0.001
R87004 out.n4478 out.n4463 0.001
R87005 out.n4478 out.n4477 0.001
R87006 out.n4441 out.n4425 0.001
R87007 out.n4441 out.n4440 0.001
R87008 out.n4414 out.n4397 0.001
R87009 out.n4414 out.n4413 0.001
R87010 out.n4378 out.n4361 0.001
R87011 out.n4378 out.n4377 0.001
R87012 out.n4349 out.n4333 0.001
R87013 out.n4349 out.n4348 0.001
R87014 out.n4313 out.n4294 0.001
R87015 out.n4313 out.n4312 0.001
R87016 out.n4282 out.n4268 0.001
R87017 out.n4282 out.n4281 0.001
R87018 out.n4247 out.n4231 0.001
R87019 out.n4247 out.n4246 0.001
R87020 out.n4219 out.n4202 0.001
R87021 out.n4219 out.n4218 0.001
R87022 out.n4183 out.n4168 0.001
R87023 out.n4183 out.n4182 0.001
R87024 out.n4155 out.n4136 0.001
R87025 out.n4155 out.n4154 0.001
R87026 out.n4120 out.n4105 0.001
R87027 out.n4120 out.n4119 0.001
R87028 out.n4092 out.n4075 0.001
R87029 out.n4092 out.n4091 0.001
R87030 out.n4054 out.n4038 0.001
R87031 out.n4054 out.n4053 0.001
R87032 out.n4026 out.n4009 0.001
R87033 out.n4026 out.n4025 0.001
R87034 out.n4942 out.n4923 0.001
R87035 out.n4942 out.n4941 0.001
R87036 out.n919 out.n917 0.001
R87037 out.n858 out.n839 0.001
R87038 out.n858 out.n857 0.001
R87039 out.n828 out.n811 0.001
R87040 out.n828 out.n827 0.001
R87041 out.n791 out.n777 0.001
R87042 out.n791 out.n790 0.001
R87043 out.n768 out.n748 0.001
R87044 out.n768 out.n767 0.001
R87045 out.n729 out.n717 0.001
R87046 out.n729 out.n728 0.001
R87047 out.n705 out.n687 0.001
R87048 out.n705 out.n704 0.001
R87049 out.n664 out.n648 0.001
R87050 out.n664 out.n663 0.001
R87051 out.n638 out.n621 0.001
R87052 out.n638 out.n637 0.001
R87053 out.n601 out.n583 0.001
R87054 out.n601 out.n600 0.001
R87055 out.n572 out.n556 0.001
R87056 out.n572 out.n571 0.001
R87057 out.n533 out.n519 0.001
R87058 out.n533 out.n532 0.001
R87059 out.n511 out.n494 0.001
R87060 out.n511 out.n510 0.001
R87061 out.n472 out.n454 0.001
R87062 out.n472 out.n471 0.001
R87063 out.n444 out.n428 0.001
R87064 out.n444 out.n443 0.001
R87065 out.n409 out.n392 0.001
R87066 out.n409 out.n408 0.001
R87067 out.n381 out.n365 0.001
R87068 out.n381 out.n380 0.001
R87069 out.n344 out.n326 0.001
R87070 out.n344 out.n343 0.001
R87071 out.n313 out.n296 0.001
R87072 out.n313 out.n312 0.001
R87073 out.n274 out.n260 0.001
R87074 out.n274 out.n273 0.001
R87075 out.n251 out.n250 0.001
R87076 out.n213 out.n196 0.001
R87077 out.n213 out.n212 0.001
R87078 out.n185 out.n168 0.001
R87079 out.n185 out.n184 0.001
R87080 out.n148 out.n131 0.001
R87081 out.n148 out.n147 0.001
R87082 out.n119 out.n104 0.001
R87083 out.n119 out.n118 0.001
R87084 out.n88 out.n87 0.001
R87085 out.n56 out.n32 0.001
R87086 out.n56 out.n23 0.001
R87087 out.n119 out.n98 0.001
R87088 out.n185 out.n162 0.001
R87089 out.n251 out.n228 0.001
R87090 out.n313 out.n289 0.001
R87091 out.n381 out.n358 0.001
R87092 out.n444 out.n422 0.001
R87093 out.n511 out.n488 0.001
R87094 out.n572 out.n550 0.001
R87095 out.n638 out.n615 0.001
R87096 out.n705 out.n680 0.001
R87097 out.n768 out.n742 0.001
R87098 out.n828 out.n805 0.001
R87099 out.n919 out.n873 0.001
R87100 out.n4026 out.n4003 0.001
R87101 out.n4092 out.n4068 0.001
R87102 out.n4155 out.n4130 0.001
R87103 out.n4219 out.n4196 0.001
R87104 out.n4282 out.n4262 0.001
R87105 out.n4349 out.n4327 0.001
R87106 out.n4414 out.n4391 0.001
R87107 out.n4478 out.n4457 0.001
R87108 out.n4541 out.n4519 0.001
R87109 out.n4609 out.n4584 0.001
R87110 out.n4673 out.n4649 0.001
R87111 out.n4737 out.n4714 0.001
R87112 out.n4800 out.n4777 0.001
R87113 out.n4835 out.n4806 0.001
R87114 out.n4800 out.n4774 0.001
R87115 out.n4800 out.n4775 0.001
R87116 out.n4763 out.n4741 0.001
R87117 out.n4763 out.n4743 0.001
R87118 out.n4737 out.n4710 0.001
R87119 out.n4737 out.n4712 0.001
R87120 out.n4699 out.n4676 0.001
R87121 out.n4699 out.n4678 0.001
R87122 out.n4673 out.n4646 0.001
R87123 out.n4673 out.n4647 0.001
R87124 out.n4637 out.n4613 0.001
R87125 out.n4637 out.n4615 0.001
R87126 out.n4609 out.n4581 0.001
R87127 out.n4609 out.n4582 0.001
R87128 out.n4570 out.n4544 0.001
R87129 out.n4570 out.n4546 0.001
R87130 out.n4541 out.n4516 0.001
R87131 out.n4541 out.n4517 0.001
R87132 out.n4506 out.n4483 0.001
R87133 out.n4506 out.n4484 0.001
R87134 out.n4478 out.n4454 0.001
R87135 out.n4478 out.n4455 0.001
R87136 out.n4441 out.n4418 0.001
R87137 out.n4441 out.n4419 0.001
R87138 out.n4414 out.n4388 0.001
R87139 out.n4414 out.n4389 0.001
R87140 out.n4378 out.n4353 0.001
R87141 out.n4378 out.n4355 0.001
R87142 out.n4349 out.n4324 0.001
R87143 out.n4349 out.n4325 0.001
R87144 out.n4313 out.n4287 0.001
R87145 out.n4313 out.n4289 0.001
R87146 out.n4282 out.n4259 0.001
R87147 out.n4282 out.n4261 0.001
R87148 out.n4247 out.n4224 0.001
R87149 out.n4247 out.n4226 0.001
R87150 out.n4219 out.n4194 0.001
R87151 out.n4219 out.n4195 0.001
R87152 out.n4183 out.n4160 0.001
R87153 out.n4183 out.n4162 0.001
R87154 out.n4155 out.n4128 0.001
R87155 out.n4155 out.n4129 0.001
R87156 out.n4120 out.n4097 0.001
R87157 out.n4120 out.n4099 0.001
R87158 out.n4092 out.n4066 0.001
R87159 out.n4092 out.n4067 0.001
R87160 out.n4054 out.n4031 0.001
R87161 out.n4054 out.n4033 0.001
R87162 out.n4026 out.n4000 0.001
R87163 out.n4026 out.n4002 0.001
R87164 out.n4942 out.n4915 0.001
R87165 out.n4942 out.n4917 0.001
R87166 out.n919 out.n871 0.001
R87167 out.n858 out.n832 0.001
R87168 out.n858 out.n833 0.001
R87169 out.n828 out.n801 0.001
R87170 out.n828 out.n803 0.001
R87171 out.n791 out.n772 0.001
R87172 out.n791 out.n773 0.001
R87173 out.n768 out.n738 0.001
R87174 out.n768 out.n739 0.001
R87175 out.n729 out.n709 0.001
R87176 out.n729 out.n711 0.001
R87177 out.n705 out.n676 0.001
R87178 out.n705 out.n678 0.001
R87179 out.n664 out.n642 0.001
R87180 out.n664 out.n644 0.001
R87181 out.n638 out.n612 0.001
R87182 out.n638 out.n613 0.001
R87183 out.n601 out.n576 0.001
R87184 out.n601 out.n577 0.001
R87185 out.n572 out.n545 0.001
R87186 out.n572 out.n547 0.001
R87187 out.n533 out.n514 0.001
R87188 out.n533 out.n515 0.001
R87189 out.n511 out.n483 0.001
R87190 out.n511 out.n485 0.001
R87191 out.n472 out.n448 0.001
R87192 out.n472 out.n450 0.001
R87193 out.n444 out.n419 0.001
R87194 out.n444 out.n420 0.001
R87195 out.n409 out.n384 0.001
R87196 out.n409 out.n386 0.001
R87197 out.n381 out.n355 0.001
R87198 out.n381 out.n356 0.001
R87199 out.n344 out.n318 0.001
R87200 out.n344 out.n320 0.001
R87201 out.n313 out.n286 0.001
R87202 out.n313 out.n288 0.001
R87203 out.n274 out.n254 0.001
R87204 out.n274 out.n256 0.001
R87205 out.n251 out.n224 0.001
R87206 out.n251 out.n226 0.001
R87207 out.n213 out.n190 0.001
R87208 out.n213 out.n192 0.001
R87209 out.n185 out.n159 0.001
R87210 out.n185 out.n161 0.001
R87211 out.n148 out.n124 0.001
R87212 out.n148 out.n126 0.001
R87213 out.n119 out.n96 0.001
R87214 out.n119 out.n97 0.001
R87215 out.n88 out.n61 0.001
R87216 out.n88 out.n63 0.001
R87217 out.n56 out.n19 0.001
R87218 out.n56 out.n22 0.001
R87219 out.n4800 out.n4772 0.001
R87220 out.n4737 out.n4708 0.001
R87221 out.n4673 out.n4645 0.001
R87222 out.n4609 out.n4580 0.001
R87223 out.n4541 out.n4515 0.001
R87224 out.n4478 out.n4452 0.001
R87225 out.n4414 out.n4387 0.001
R87226 out.n4349 out.n4323 0.001
R87227 out.n4282 out.n4257 0.001
R87228 out.n4219 out.n4193 0.001
R87229 out.n4155 out.n4127 0.001
R87230 out.n4092 out.n4064 0.001
R87231 out.n4026 out.n3998 0.001
R87232 out.n4942 out.n4913 0.001
R87233 out.n919 out.n869 0.001
R87234 out.n828 out.n800 0.001
R87235 out.n768 out.n736 0.001
R87236 out.n705 out.n674 0.001
R87237 out.n638 out.n610 0.001
R87238 out.n572 out.n544 0.001
R87239 out.n511 out.n481 0.001
R87240 out.n444 out.n417 0.001
R87241 out.n381 out.n353 0.001
R87242 out.n313 out.n284 0.001
R87243 out.n251 out.n222 0.001
R87244 out.n185 out.n157 0.001
R87245 out.n119 out.n95 0.001
R87246 out.n56 out.n18 0.001
R87247 out.n9506 out.n9499 0.001
R87248 out.n9506 out.n9500 0.001
R87249 out.n8796 out.n8795 0.001
R87250 out.n7 out.n6 0.001
R87251 out.n17308 out.n17307 0.001
R87252 out.n12403 out.n12402 0.001
R87253 out.n3145 out.n3144 0.001
R87254 out.n17187 out.n17186 0.001
R87255 out.n17190 out.n17189 0.001
R87256 out.n17191 out.n17190 0.001
R87257 out.n17194 out.n17193 0.001
R87258 out.n17195 out.n17194 0.001
R87259 out.n17198 out.n17197 0.001
R87260 out.n17199 out.n17198 0.001
R87261 out.n17202 out.n17201 0.001
R87262 out.n17203 out.n17202 0.001
R87263 out.n17206 out.n17205 0.001
R87264 out.n17207 out.n17206 0.001
R87265 out.n17210 out.n17209 0.001
R87266 out.n17211 out.n17210 0.001
R87267 out.n17214 out.n17213 0.001
R87268 out.n17215 out.n17214 0.001
R87269 out.n17218 out.n17217 0.001
R87270 out.n17219 out.n17218 0.001
R87271 out.n17222 out.n17221 0.001
R87272 out.n17223 out.n17222 0.001
R87273 out.n17226 out.n17225 0.001
R87274 out.n17227 out.n17226 0.001
R87275 out.n17230 out.n17229 0.001
R87276 out.n17231 out.n17230 0.001
R87277 out.n17234 out.n17233 0.001
R87278 out.n17235 out.n17234 0.001
R87279 out.n17238 out.n17237 0.001
R87280 out.n17239 out.n17238 0.001
R87281 out.n10001 out.n9999 0.001
R87282 out.n9999 out.n9998 0.001
R87283 out.n9964 out.n9963 0.001
R87284 out.n9963 out.n9962 0.001
R87285 out.n9926 out.n9925 0.001
R87286 out.n9892 out.n9891 0.001
R87287 out.n9858 out.n9856 0.001
R87288 out.n9856 out.n9855 0.001
R87289 out.n9821 out.n9820 0.001
R87290 out.n9820 out.n9819 0.001
R87291 out.n9785 out.n9784 0.001
R87292 out.n9784 out.n9783 0.001
R87293 out.n9749 out.n9748 0.001
R87294 out.n9748 out.n9747 0.001
R87295 out.n9713 out.n9712 0.001
R87296 out.n9712 out.n9711 0.001
R87297 out.n9677 out.n9676 0.001
R87298 out.n9676 out.n9675 0.001
R87299 out.n9619 out.n9617 0.001
R87300 out.n9617 out.n9616 0.001
R87301 out.n9582 out.n9581 0.001
R87302 out.n9581 out.n9580 0.001
R87303 out.n9546 out.n9545 0.001
R87304 out.n9545 out.n9544 0.001
R87305 out.n9510 out.n9509 0.001
R87306 out.n16285 out.n10007 0.001
R87307 out.n16285 out.n10036 0.001
R87308 out.n17142 out.n17124 0.001
R87309 out.n17110 out.n17098 0.001
R87310 out.n17075 out.n17060 0.001
R87311 out.n17044 out.n17032 0.001
R87312 out.n17009 out.n16996 0.001
R87313 out.n16980 out.n16966 0.001
R87314 out.n16943 out.n16928 0.001
R87315 out.n16912 out.n16900 0.001
R87316 out.n16877 out.n16864 0.001
R87317 out.n16848 out.n16834 0.001
R87318 out.n16811 out.n16798 0.001
R87319 out.n16782 out.n16768 0.001
R87320 out.n16745 out.n16730 0.001
R87321 out.n16714 out.n16702 0.001
R87322 out.n16679 out.n16664 0.001
R87323 out.n16648 out.n16636 0.001
R87324 out.n16613 out.n16600 0.001
R87325 out.n16584 out.n16570 0.001
R87326 out.n16547 out.n16532 0.001
R87327 out.n16516 out.n16506 0.001
R87328 out.n16483 out.n16466 0.001
R87329 out.n16450 out.n16440 0.001
R87330 out.n16417 out.n16400 0.001
R87331 out.n16384 out.n16372 0.001
R87332 out.n16349 out.n16334 0.001
R87333 out.n16318 out.n16306 0.001
R87334 out.n16285 out.n10037 0.001
R87335 out.n9994 out.n9979 0.001
R87336 out.n9084 out.n9074 0.001
R87337 out.n9958 out.n9941 0.001
R87338 out.n9922 out.n9910 0.001
R87339 out.n9890 out.n9875 0.001
R87340 out.n9119 out.n9107 0.001
R87341 out.n9851 out.n9836 0.001
R87342 out.n9153 out.n9141 0.001
R87343 out.n9815 out.n9800 0.001
R87344 out.n9187 out.n9175 0.001
R87345 out.n9779 out.n9764 0.001
R87346 out.n9221 out.n9209 0.001
R87347 out.n9743 out.n9728 0.001
R87348 out.n9255 out.n9243 0.001
R87349 out.n9707 out.n9692 0.001
R87350 out.n9289 out.n9277 0.001
R87351 out.n9651 out.n9636 0.001
R87352 out.n9322 out.n9310 0.001
R87353 out.n9612 out.n9597 0.001
R87354 out.n9356 out.n9344 0.001
R87355 out.n9576 out.n9561 0.001
R87356 out.n9390 out.n9378 0.001
R87357 out.n9540 out.n9525 0.001
R87358 out.n9423 out.n9410 0.001
R87359 out.n9506 out.n9494 0.001
R87360 out.n16285 out.n16274 0.001
R87361 out.n16285 out.n10030 0.001
R87362 out.n16285 out.n16279 0.001
R87363 out.n16285 out.n10025 0.001
R87364 out.n16285 out.n10020 0.001
R87365 out.n16285 out.n16284 0.001
R87366 out.n4763 out.n4746 0.001
R87367 out.n4699 out.n4681 0.001
R87368 out.n4637 out.n4619 0.001
R87369 out.n4570 out.n4551 0.001
R87370 out.n4506 out.n4487 0.001
R87371 out.n4441 out.n4423 0.001
R87372 out.n4378 out.n4359 0.001
R87373 out.n4313 out.n4292 0.001
R87374 out.n4247 out.n4229 0.001
R87375 out.n4183 out.n4166 0.001
R87376 out.n4120 out.n4103 0.001
R87377 out.n4054 out.n4036 0.001
R87378 out.n4942 out.n4921 0.001
R87379 out.n919 out.n881 0.001
R87380 out.n858 out.n837 0.001
R87381 out.n791 out.n775 0.001
R87382 out.n729 out.n715 0.001
R87383 out.n664 out.n646 0.001
R87384 out.n601 out.n581 0.001
R87385 out.n533 out.n517 0.001
R87386 out.n472 out.n452 0.001
R87387 out.n409 out.n390 0.001
R87388 out.n344 out.n324 0.001
R87389 out.n274 out.n258 0.001
R87390 out.n213 out.n194 0.001
R87391 out.n148 out.n129 0.001
R87392 out.n88 out.n68 0.001
R87393 out.n4800 out.n4781 0.001
R87394 out.n4737 out.n4718 0.001
R87395 out.n4673 out.n4653 0.001
R87396 out.n4609 out.n4588 0.001
R87397 out.n4541 out.n4523 0.001
R87398 out.n4478 out.n4461 0.001
R87399 out.n4414 out.n4395 0.001
R87400 out.n4349 out.n4331 0.001
R87401 out.n4282 out.n4266 0.001
R87402 out.n4219 out.n4200 0.001
R87403 out.n4155 out.n4134 0.001
R87404 out.n4092 out.n4072 0.001
R87405 out.n4026 out.n4007 0.001
R87406 out.n4942 out.n4919 0.001
R87407 out.n919 out.n875 0.001
R87408 out.n828 out.n809 0.001
R87409 out.n768 out.n746 0.001
R87410 out.n705 out.n684 0.001
R87411 out.n638 out.n619 0.001
R87412 out.n572 out.n554 0.001
R87413 out.n511 out.n492 0.001
R87414 out.n444 out.n426 0.001
R87415 out.n381 out.n362 0.001
R87416 out.n313 out.n293 0.001
R87417 out.n251 out.n232 0.001
R87418 out.n185 out.n166 0.001
R87419 out.n119 out.n102 0.001
R87420 out.n8869 out.n91 0.001
R87421 out.n8869 out.n58 0.001
R87422 out.n8863 out.n152 0.001
R87423 out.n8863 out.n121 0.001
R87424 out.n8857 out.n217 0.001
R87425 out.n8857 out.n187 0.001
R87426 out.n8851 out.n277 0.001
R87427 out.n8851 out.n253 0.001
R87428 out.n8846 out.n347 0.001
R87429 out.n8846 out.n315 0.001
R87430 out.n8842 out.n412 0.001
R87431 out.n8842 out.n383 0.001
R87432 out.n8836 out.n476 0.001
R87433 out.n8836 out.n446 0.001
R87434 out.n8830 out.n537 0.001
R87435 out.n8830 out.n513 0.001
R87436 out.n8825 out.n605 0.001
R87437 out.n8825 out.n574 0.001
R87438 out.n8819 out.n668 0.001
R87439 out.n8819 out.n640 0.001
R87440 out.n8814 out.n732 0.001
R87441 out.n8814 out.n707 0.001
R87442 out.n8808 out.n795 0.001
R87443 out.n8808 out.n770 0.001
R87444 out.n8802 out.n862 0.001
R87445 out.n8802 out.n830 0.001
R87446 out.n8796 out.n4910 0.001
R87447 out.n4904 out.n4058 0.001
R87448 out.n4904 out.n4028 0.001
R87449 out.n4899 out.n4123 0.001
R87450 out.n4899 out.n4094 0.001
R87451 out.n4893 out.n4187 0.001
R87452 out.n4893 out.n4157 0.001
R87453 out.n4888 out.n4251 0.001
R87454 out.n4888 out.n4221 0.001
R87455 out.n4883 out.n4317 0.001
R87456 out.n4883 out.n4284 0.001
R87457 out.n4878 out.n4382 0.001
R87458 out.n4878 out.n4351 0.001
R87459 out.n4872 out.n4445 0.001
R87460 out.n4872 out.n4416 0.001
R87461 out.n4867 out.n4510 0.001
R87462 out.n4867 out.n4480 0.001
R87463 out.n4861 out.n4574 0.001
R87464 out.n4861 out.n4543 0.001
R87465 out.n4856 out.n4640 0.001
R87466 out.n4856 out.n4611 0.001
R87467 out.n4850 out.n4702 0.001
R87468 out.n4850 out.n4675 0.001
R87469 out.n4844 out.n4767 0.001
R87470 out.n4844 out.n4739 0.001
R87471 out.n4838 out.n4804 0.001
R87472 out.n4835 out.n4813 0.001
R87473 out.n4800 out.n4779 0.001
R87474 out.n4763 out.n4744 0.001
R87475 out.n4737 out.n4716 0.001
R87476 out.n4699 out.n4680 0.001
R87477 out.n4673 out.n4651 0.001
R87478 out.n4637 out.n4617 0.001
R87479 out.n4609 out.n4586 0.001
R87480 out.n4570 out.n4549 0.001
R87481 out.n4541 out.n4521 0.001
R87482 out.n4506 out.n4485 0.001
R87483 out.n4478 out.n4459 0.001
R87484 out.n4441 out.n4421 0.001
R87485 out.n4414 out.n4393 0.001
R87486 out.n4378 out.n4357 0.001
R87487 out.n4349 out.n4329 0.001
R87488 out.n4313 out.n4290 0.001
R87489 out.n4282 out.n4264 0.001
R87490 out.n4247 out.n4228 0.001
R87491 out.n4219 out.n4198 0.001
R87492 out.n4183 out.n4164 0.001
R87493 out.n4155 out.n4132 0.001
R87494 out.n4120 out.n4101 0.001
R87495 out.n4092 out.n4070 0.001
R87496 out.n4054 out.n4034 0.001
R87497 out.n4026 out.n4005 0.001
R87498 out.n858 out.n836 0.001
R87499 out.n828 out.n807 0.001
R87500 out.n791 out.n774 0.001
R87501 out.n768 out.n744 0.001
R87502 out.n729 out.n713 0.001
R87503 out.n705 out.n682 0.001
R87504 out.n664 out.n645 0.001
R87505 out.n638 out.n617 0.001
R87506 out.n601 out.n579 0.001
R87507 out.n572 out.n552 0.001
R87508 out.n533 out.n516 0.001
R87509 out.n511 out.n490 0.001
R87510 out.n472 out.n451 0.001
R87511 out.n444 out.n424 0.001
R87512 out.n409 out.n388 0.001
R87513 out.n381 out.n360 0.001
R87514 out.n344 out.n322 0.001
R87515 out.n313 out.n291 0.001
R87516 out.n274 out.n257 0.001
R87517 out.n251 out.n230 0.001
R87518 out.n213 out.n193 0.001
R87519 out.n185 out.n164 0.001
R87520 out.n148 out.n128 0.001
R87521 out.n119 out.n100 0.001
R87522 out.n88 out.n66 0.001
R87523 out.n56 out.n25 0.001
R87524 out.n56 out.n30 0.001
R87525 out.n4835 out.n4824 0.001
R87526 out.n4800 out.n4787 0.001
R87527 out.n4800 out.n4791 0.001
R87528 out.n4763 out.n4753 0.001
R87529 out.n4737 out.n4726 0.001
R87530 out.n4737 out.n4729 0.001
R87531 out.n4699 out.n4690 0.001
R87532 out.n4673 out.n4662 0.001
R87533 out.n4673 out.n4665 0.001
R87534 out.n4637 out.n4628 0.001
R87535 out.n4609 out.n4597 0.001
R87536 out.n4609 out.n4601 0.001
R87537 out.n4570 out.n4561 0.001
R87538 out.n4541 out.n4529 0.001
R87539 out.n4541 out.n4534 0.001
R87540 out.n4506 out.n4495 0.001
R87541 out.n4478 out.n4467 0.001
R87542 out.n4478 out.n4470 0.001
R87543 out.n4441 out.n4433 0.001
R87544 out.n4414 out.n4402 0.001
R87545 out.n4414 out.n4405 0.001
R87546 out.n4378 out.n4368 0.001
R87547 out.n4349 out.n4336 0.001
R87548 out.n4349 out.n4341 0.001
R87549 out.n4313 out.n4301 0.001
R87550 out.n4282 out.n4272 0.001
R87551 out.n4282 out.n4275 0.001
R87552 out.n4247 out.n4238 0.001
R87553 out.n4219 out.n4208 0.001
R87554 out.n4219 out.n4211 0.001
R87555 out.n4183 out.n4175 0.001
R87556 out.n4155 out.n4142 0.001
R87557 out.n4155 out.n4146 0.001
R87558 out.n4120 out.n4112 0.001
R87559 out.n4092 out.n4081 0.001
R87560 out.n4092 out.n4084 0.001
R87561 out.n4054 out.n4045 0.001
R87562 out.n4026 out.n4015 0.001
R87563 out.n4026 out.n4018 0.001
R87564 out.n919 out.n893 0.001
R87565 out.n919 out.n913 0.001
R87566 out.n858 out.n847 0.001
R87567 out.n828 out.n815 0.001
R87568 out.n828 out.n820 0.001
R87569 out.n791 out.n782 0.001
R87570 out.n768 out.n752 0.001
R87571 out.n768 out.n757 0.001
R87572 out.n729 out.n722 0.001
R87573 out.n705 out.n693 0.001
R87574 out.n705 out.n697 0.001
R87575 out.n664 out.n655 0.001
R87576 out.n638 out.n627 0.001
R87577 out.n638 out.n630 0.001
R87578 out.n601 out.n591 0.001
R87579 out.n572 out.n559 0.001
R87580 out.n572 out.n564 0.001
R87581 out.n533 out.n523 0.001
R87582 out.n511 out.n499 0.001
R87583 out.n511 out.n502 0.001
R87584 out.n472 out.n462 0.001
R87585 out.n444 out.n433 0.001
R87586 out.n444 out.n436 0.001
R87587 out.n409 out.n400 0.001
R87588 out.n381 out.n370 0.001
R87589 out.n381 out.n373 0.001
R87590 out.n344 out.n335 0.001
R87591 out.n313 out.n301 0.001
R87592 out.n313 out.n306 0.001
R87593 out.n274 out.n265 0.001
R87594 out.n251 out.n241 0.001
R87595 out.n251 out.n244 0.001
R87596 out.n213 out.n203 0.001
R87597 out.n185 out.n174 0.001
R87598 out.n185 out.n178 0.001
R87599 out.n148 out.n138 0.001
R87600 out.n119 out.n109 0.001
R87601 out.n119 out.n112 0.001
R87602 out.n88 out.n78 0.001
R87603 out.n56 out.n44 0.001
R87604 out.n56 out.n55 0.001
R87605 out.n119 out.n116 0.001
R87606 out.n185 out.n183 0.001
R87607 out.n251 out.n249 0.001
R87608 out.n313 out.n310 0.001
R87609 out.n381 out.n378 0.001
R87610 out.n444 out.n441 0.001
R87611 out.n511 out.n509 0.001
R87612 out.n572 out.n570 0.001
R87613 out.n638 out.n635 0.001
R87614 out.n705 out.n703 0.001
R87615 out.n768 out.n765 0.001
R87616 out.n828 out.n825 0.001
R87617 out.n919 out.n916 0.001
R87618 out.n4026 out.n4023 0.001
R87619 out.n4092 out.n4089 0.001
R87620 out.n4155 out.n4152 0.001
R87621 out.n4219 out.n4216 0.001
R87622 out.n4282 out.n4279 0.001
R87623 out.n4349 out.n4347 0.001
R87624 out.n4414 out.n4411 0.001
R87625 out.n4478 out.n4475 0.001
R87626 out.n4541 out.n4539 0.001
R87627 out.n4609 out.n4606 0.001
R87628 out.n4673 out.n4670 0.001
R87629 out.n4737 out.n4734 0.001
R87630 out.n4800 out.n4797 0.001
R87631 out.n919 out.n887 0.001
R87632 out.n4835 out.n4829 0.001
R87633 out.n4763 out.n4759 0.001
R87634 out.n4699 out.n4695 0.001
R87635 out.n4637 out.n4633 0.001
R87636 out.n4570 out.n4566 0.001
R87637 out.n4506 out.n4501 0.001
R87638 out.n4441 out.n4437 0.001
R87639 out.n4378 out.n4374 0.001
R87640 out.n4313 out.n4308 0.001
R87641 out.n4247 out.n4243 0.001
R87642 out.n4183 out.n4179 0.001
R87643 out.n4120 out.n4116 0.001
R87644 out.n4054 out.n4050 0.001
R87645 out.n4942 out.n4938 0.001
R87646 out.n858 out.n853 0.001
R87647 out.n791 out.n787 0.001
R87648 out.n729 out.n725 0.001
R87649 out.n664 out.n659 0.001
R87650 out.n601 out.n597 0.001
R87651 out.n533 out.n528 0.001
R87652 out.n472 out.n467 0.001
R87653 out.n409 out.n405 0.001
R87654 out.n344 out.n340 0.001
R87655 out.n274 out.n270 0.001
R87656 out.n213 out.n208 0.001
R87657 out.n148 out.n143 0.001
R87658 out.n88 out.n84 0.001
R87659 out.n919 out.n884 0.001
R87660 out.n8871 out.n11 0.001
R87661 out.n8866 out.n93 0.001
R87662 out.n8860 out.n154 0.001
R87663 out.n8854 out.n219 0.001
R87664 out.n8848 out.n280 0.001
R87665 out.n8844 out.n351 0.001
R87666 out.n8839 out.n414 0.001
R87667 out.n8833 out.n478 0.001
R87668 out.n8827 out.n540 0.001
R87669 out.n8822 out.n607 0.001
R87670 out.n8817 out.n671 0.001
R87671 out.n8811 out.n734 0.001
R87672 out.n8805 out.n797 0.001
R87673 out.n4906 out.n3996 0.001
R87674 out.n4902 out.n4061 0.001
R87675 out.n4896 out.n4125 0.001
R87676 out.n4890 out.n4190 0.001
R87677 out.n4886 out.n4254 0.001
R87678 out.n4881 out.n4320 0.001
R87679 out.n4875 out.n4384 0.001
R87680 out.n4870 out.n4448 0.001
R87681 out.n4864 out.n4512 0.001
R87682 out.n4859 out.n4577 0.001
R87683 out.n4853 out.n4642 0.001
R87684 out.n4847 out.n4704 0.001
R87685 out.n4841 out.n4769 0.001
R87686 out.n4841 out.n4768 0.001
R87687 out.n4847 out.n4703 0.001
R87688 out.n4853 out.n4641 0.001
R87689 out.n4859 out.n4576 0.001
R87690 out.n4864 out.n4511 0.001
R87691 out.n4870 out.n4447 0.001
R87692 out.n4875 out.n4383 0.001
R87693 out.n4881 out.n4319 0.001
R87694 out.n4886 out.n4253 0.001
R87695 out.n4890 out.n4188 0.001
R87696 out.n4896 out.n4124 0.001
R87697 out.n4902 out.n4060 0.001
R87698 out.n4906 out.n3994 0.001
R87699 out.n8799 out.n867 0.001
R87700 out.n8799 out.n921 0.001
R87701 out.n8805 out.n796 0.001
R87702 out.n8811 out.n733 0.001
R87703 out.n8817 out.n670 0.001
R87704 out.n8822 out.n606 0.001
R87705 out.n8827 out.n538 0.001
R87706 out.n8833 out.n477 0.001
R87707 out.n8839 out.n413 0.001
R87708 out.n8844 out.n349 0.001
R87709 out.n8848 out.n278 0.001
R87710 out.n8854 out.n218 0.001
R87711 out.n8860 out.n153 0.001
R87712 out.n8866 out.n92 0.001
R87713 out.n8871 out.n9 0.001
R87714 out.n8796 out.n3993 0.001
R87715 out.n16077 out.n15941 0.001
R87716 out.n15121 out.n15120 0.001
R87717 out.n14105 out.n14104 0.001
R87718 out.n9506 out.n9473 0.001
R87719 out.n1531 out.n1530 0.001
R87720 out.n2378 out.n2377 0.001
R87721 out.n14137 out.n14136 0.001
R87722 out.n3085 out.n3084 0.001
R87723 out.n15426 out.n15413 0.001
R87724 out.n10009 out.n10008 0.001
R87725 out.n15433 out.n15432 0.001
R87726 out.n8981 out.n8980 0.001
R87727 out.n17306 out.n17305 0.001
R87728 out.n16075 out.n16074 0.001
R87729 out.n8918 out.n8917 0.001
R87730 out.n9437 out.n9430 0.001
R87731 out.n10270 out.n10265 0.001
R87732 out.n10259 out.n10256 0.001
R87733 out.n10246 out.n10245 0.001
R87734 out.n10239 out.n10238 0.001
R87735 out.n10235 out.n10233 0.001
R87736 out.n10221 out.n10216 0.001
R87737 out.n10205 out.n10204 0.001
R87738 out.n10199 out.n10196 0.001
R87739 out.n10164 out.n10161 0.001
R87740 out.n10159 out.n10158 0.001
R87741 out.n10144 out.n10142 0.001
R87742 out.n10139 out.n10135 0.001
R87743 out.n13230 out.n13229 0.001
R87744 out.n13229 out.n13226 0.001
R87745 out.n13224 out.n13223 0.001
R87746 out.n13078 out.n13075 0.001
R87747 out.n12967 out.n12964 0.001
R87748 out.n12963 out.n12961 0.001
R87749 out.n12798 out.n12797 0.001
R87750 out.n12656 out.n12653 0.001
R87751 out.n12652 out.n12650 0.001
R87752 out.n12540 out.n12537 0.001
R87753 out.n12536 out.n12535 0.001
R87754 out.n12365 out.n12364 0.001
R87755 out.n12364 out.n12361 0.001
R87756 out.n12359 out.n12358 0.001
R87757 out.n12213 out.n12210 0.001
R87758 out.n12102 out.n12099 0.001
R87759 out.n12098 out.n12096 0.001
R87760 out.n13632 out.n13631 0.001
R87761 out.n13489 out.n13486 0.001
R87762 out.n13485 out.n13483 0.001
R87763 out.n13373 out.n13370 0.001
R87764 out.n13369 out.n13368 0.001
R87765 out.n11534 out.n11533 0.001
R87766 out.n11533 out.n11530 0.001
R87767 out.n11528 out.n11527 0.001
R87768 out.n11387 out.n11384 0.001
R87769 out.n11279 out.n11276 0.001
R87770 out.n11275 out.n11273 0.001
R87771 out.n11107 out.n11106 0.001
R87772 out.n11106 out.n11103 0.001
R87773 out.n11101 out.n11100 0.001
R87774 out.n10960 out.n10957 0.001
R87775 out.n10849 out.n10846 0.001
R87776 out.n10845 out.n10843 0.001
R87777 out.n11945 out.n11944 0.001
R87778 out.n11944 out.n11941 0.001
R87779 out.n11939 out.n11938 0.001
R87780 out.n11793 out.n11790 0.001
R87781 out.n11682 out.n11679 0.001
R87782 out.n11678 out.n11676 0.001
R87783 out.n14087 out.n14086 0.001
R87784 out.n13944 out.n13941 0.001
R87785 out.n13940 out.n13938 0.001
R87786 out.n13828 out.n13825 0.001
R87787 out.n13824 out.n13823 0.001
R87788 out.n10678 out.n10677 0.001
R87789 out.n10677 out.n10674 0.001
R87790 out.n10672 out.n10671 0.001
R87791 out.n10526 out.n10523 0.001
R87792 out.n10415 out.n10412 0.001
R87793 out.n10411 out.n10409 0.001
R87794 out.n14539 out.n14536 0.001
R87795 out.n14534 out.n14533 0.001
R87796 out.n14491 out.n14488 0.001
R87797 out.n14486 out.n14485 0.001
R87798 out.n14422 out.n14419 0.001
R87799 out.n14561 out.n14560 0.001
R87800 out.n14553 out.n14552 0.001
R87801 out.n14552 out.n14551 0.001
R87802 out.n15567 out.n15566 0.001
R87803 out.n15373 out.n15372 0.001
R87804 out.n16205 out.n16204 0.001
R87805 out.n15125 out.n15124 0.001
R87806 out.n14109 out.n14108 0.001
R87807 out.n16285 out.n16269 0.001
R87808 out.n9506 out.n9493 0.001
R87809 out.n14104 out.n14103 0.001
R87810 out.n14589 out.n14588 0.001
R87811 out.n14599 out.n14598 0.001
R87812 out.n14624 out.n14623 0.001
R87813 out.n14635 out.n14634 0.001
R87814 out.n14660 out.n14659 0.001
R87815 out.n14670 out.n14669 0.001
R87816 out.n14695 out.n14694 0.001
R87817 out.n14706 out.n14705 0.001
R87818 out.n14731 out.n14730 0.001
R87819 out.n14741 out.n14740 0.001
R87820 out.n14766 out.n14765 0.001
R87821 out.n14777 out.n14776 0.001
R87822 out.n14802 out.n14801 0.001
R87823 out.n14812 out.n14811 0.001
R87824 out.n14837 out.n14836 0.001
R87825 out.n14848 out.n14847 0.001
R87826 out.n14873 out.n14872 0.001
R87827 out.n14883 out.n14882 0.001
R87828 out.n14908 out.n14907 0.001
R87829 out.n14919 out.n14918 0.001
R87830 out.n14944 out.n14943 0.001
R87831 out.n14954 out.n14953 0.001
R87832 out.n14979 out.n14978 0.001
R87833 out.n14990 out.n14989 0.001
R87834 out.n15012 out.n15011 0.001
R87835 out.n15022 out.n15021 0.001
R87836 out.n15044 out.n15043 0.001
R87837 out.n15055 out.n15054 0.001
R87838 out.n15077 out.n15076 0.001
R87839 out.n15087 out.n15086 0.001
R87840 out.n15109 out.n15108 0.001
R87841 out.n15120 out.n15119 0.001
R87842 out.n15147 out.n15146 0.001
R87843 out.n15158 out.n15157 0.001
R87844 out.n15188 out.n15187 0.001
R87845 out.n15199 out.n15198 0.001
R87846 out.n15220 out.n15219 0.001
R87847 out.n15230 out.n15229 0.001
R87848 out.n15253 out.n15252 0.001
R87849 out.n15264 out.n15263 0.001
R87850 out.n15285 out.n15284 0.001
R87851 out.n15295 out.n15294 0.001
R87852 out.n15318 out.n15317 0.001
R87853 out.n15329 out.n15328 0.001
R87854 out.n15350 out.n15349 0.001
R87855 out.n15360 out.n15359 0.001
R87856 out.n9005 out.n9004 0.001
R87857 out.n10034 out.n10033 0.001
R87858 out.n16266 out.n16263 0.001
R87859 out.n16265 out.n16264 0.001
R87860 out.n16235 out.n16231 0.001
R87861 out.n17264 out.n17263 0.001
R87862 out.n16199 out.n16196 0.001
R87863 out.n16198 out.n16197 0.001
R87864 out.n16169 out.n16166 0.001
R87865 out.n16168 out.n16167 0.001
R87866 out.n16138 out.n16135 0.001
R87867 out.n16137 out.n16136 0.001
R87868 out.n16108 out.n16105 0.001
R87869 out.n16107 out.n16106 0.001
R87870 out.n16077 out.n16073 0.001
R87871 out.n15965 out.n15964 0.001
R87872 out.n15938 out.n15935 0.001
R87873 out.n16001 out.n16000 0.001
R87874 out.n15902 out.n15899 0.001
R87875 out.n15901 out.n15900 0.001
R87876 out.n15872 out.n15869 0.001
R87877 out.n15871 out.n15870 0.001
R87878 out.n15841 out.n15838 0.001
R87879 out.n15840 out.n15839 0.001
R87880 out.n15811 out.n15808 0.001
R87881 out.n15810 out.n15809 0.001
R87882 out.n15780 out.n15777 0.001
R87883 out.n15779 out.n15778 0.001
R87884 out.n15750 out.n15747 0.001
R87885 out.n15749 out.n15748 0.001
R87886 out.n15714 out.n15711 0.001
R87887 out.n15713 out.n15712 0.001
R87888 out.n15679 out.n15676 0.001
R87889 out.n15678 out.n15677 0.001
R87890 out.n15643 out.n15639 0.001
R87891 out.n15592 out.n15591 0.001
R87892 out.n15561 out.n15558 0.001
R87893 out.n15560 out.n15559 0.001
R87894 out.n15531 out.n15528 0.001
R87895 out.n15530 out.n15529 0.001
R87896 out.n15495 out.n15492 0.001
R87897 out.n15494 out.n15493 0.001
R87898 out.n15459 out.n15455 0.001
R87899 out.n10711 out.n10710 0.001
R87900 out.n10712 out.n10711 0.001
R87901 out.n15428 out.n15426 0.001
R87902 out.n17186 out.n17185 0.001
R87903 out.n17147 out.n17146 0.001
R87904 out.n17188 out.n17142 0.001
R87905 out.n17144 out.n17143 0.001
R87906 out.n17190 out.n17110 0.001
R87907 out.n17080 out.n17079 0.001
R87908 out.n17192 out.n17075 0.001
R87909 out.n17077 out.n17076 0.001
R87910 out.n17194 out.n17044 0.001
R87911 out.n17014 out.n17013 0.001
R87912 out.n17196 out.n17009 0.001
R87913 out.n17011 out.n17010 0.001
R87914 out.n17198 out.n16980 0.001
R87915 out.n16948 out.n16947 0.001
R87916 out.n17200 out.n16943 0.001
R87917 out.n16945 out.n16944 0.001
R87918 out.n17202 out.n16912 0.001
R87919 out.n16882 out.n16881 0.001
R87920 out.n17204 out.n16877 0.001
R87921 out.n16879 out.n16878 0.001
R87922 out.n17206 out.n16848 0.001
R87923 out.n16816 out.n16815 0.001
R87924 out.n17208 out.n16811 0.001
R87925 out.n16813 out.n16812 0.001
R87926 out.n17210 out.n16782 0.001
R87927 out.n16750 out.n16749 0.001
R87928 out.n17212 out.n16745 0.001
R87929 out.n16747 out.n16746 0.001
R87930 out.n17214 out.n16714 0.001
R87931 out.n16684 out.n16683 0.001
R87932 out.n17216 out.n16679 0.001
R87933 out.n16681 out.n16680 0.001
R87934 out.n17218 out.n16648 0.001
R87935 out.n16618 out.n16617 0.001
R87936 out.n17220 out.n16613 0.001
R87937 out.n16615 out.n16614 0.001
R87938 out.n17222 out.n16584 0.001
R87939 out.n16552 out.n16551 0.001
R87940 out.n17224 out.n16547 0.001
R87941 out.n16549 out.n16548 0.001
R87942 out.n17226 out.n16516 0.001
R87943 out.n16488 out.n16487 0.001
R87944 out.n17228 out.n16483 0.001
R87945 out.n16485 out.n16484 0.001
R87946 out.n17230 out.n16450 0.001
R87947 out.n16422 out.n16421 0.001
R87948 out.n17232 out.n16417 0.001
R87949 out.n16419 out.n16418 0.001
R87950 out.n17234 out.n16384 0.001
R87951 out.n16354 out.n16353 0.001
R87952 out.n17236 out.n16349 0.001
R87953 out.n16351 out.n16350 0.001
R87954 out.n17238 out.n16318 0.001
R87955 out.n16288 out.n16287 0.001
R87956 out.n17307 out.n16285 0.001
R87957 out.n9020 out.n9017 0.001
R87958 out.n9999 out.n9052 0.001
R87959 out.n9022 out.n9021 0.001
R87960 out.n9997 out.n9994 0.001
R87961 out.n9996 out.n9995 0.001
R87962 out.n9963 out.n9084 0.001
R87963 out.n9056 out.n9055 0.001
R87964 out.n9961 out.n9958 0.001
R87965 out.n9960 out.n9959 0.001
R87966 out.n9925 out.n9922 0.001
R87967 out.n9924 out.n9923 0.001
R87968 out.n9891 out.n9890 0.001
R87969 out.n9860 out.n9859 0.001
R87970 out.n9856 out.n9119 0.001
R87971 out.n9089 out.n9088 0.001
R87972 out.n9854 out.n9851 0.001
R87973 out.n9853 out.n9852 0.001
R87974 out.n9820 out.n9153 0.001
R87975 out.n9123 out.n9122 0.001
R87976 out.n9818 out.n9815 0.001
R87977 out.n9817 out.n9816 0.001
R87978 out.n9784 out.n9187 0.001
R87979 out.n9157 out.n9156 0.001
R87980 out.n9782 out.n9779 0.001
R87981 out.n9781 out.n9780 0.001
R87982 out.n9748 out.n9221 0.001
R87983 out.n9191 out.n9190 0.001
R87984 out.n9746 out.n9743 0.001
R87985 out.n9745 out.n9744 0.001
R87986 out.n9712 out.n9255 0.001
R87987 out.n9225 out.n9224 0.001
R87988 out.n9710 out.n9707 0.001
R87989 out.n9709 out.n9708 0.001
R87990 out.n9676 out.n9289 0.001
R87991 out.n9259 out.n9258 0.001
R87992 out.n9674 out.n9651 0.001
R87993 out.n9621 out.n9620 0.001
R87994 out.n9617 out.n9322 0.001
R87995 out.n9292 out.n9291 0.001
R87996 out.n9615 out.n9612 0.001
R87997 out.n9614 out.n9613 0.001
R87998 out.n9581 out.n9356 0.001
R87999 out.n9326 out.n9325 0.001
R88000 out.n9579 out.n9576 0.001
R88001 out.n9578 out.n9577 0.001
R88002 out.n9545 out.n9390 0.001
R88003 out.n9360 out.n9359 0.001
R88004 out.n9543 out.n9540 0.001
R88005 out.n9542 out.n9541 0.001
R88006 out.n9509 out.n9423 0.001
R88007 out.n12394 out.n12393 0.001
R88008 out.n13671 out.n13670 0.001
R88009 out.n11133 out.n11132 0.001
R88010 out.n14098 out.n13703 0.001
R88011 out.n14564 out.n14149 0.001
R88012 out.n9469 out.n9468 0.001
R88013 out.n9468 out.n9467 0.001
R88014 out.n5165 out.n5162 0.001
R88015 out.n5160 out.n5159 0.001
R88016 out.n5096 out.n5093 0.001
R88017 out.n1067 out.n1066 0.001
R88018 out.n1071 out.n1069 0.001
R88019 out.n5706 out.n5702 0.001
R88020 out.n5831 out.n5828 0.001
R88021 out.n5827 out.n5825 0.001
R88022 out.n5587 out.n5584 0.001
R88023 out.n5583 out.n5581 0.001
R88024 out.n5246 out.n5243 0.001
R88025 out.n5242 out.n5240 0.001
R88026 out.n5356 out.n5353 0.001
R88027 out.n5173 out.n5172 0.001
R88028 out.n1275 out.n1274 0.001
R88029 out.n4838 out.n4835 0.001
R88030 out.n4837 out.n4836 0.001
R88031 out.n4841 out.n4800 0.001
R88032 out.n4771 out.n4770 0.001
R88033 out.n4844 out.n4763 0.001
R88034 out.n4765 out.n4764 0.001
R88035 out.n4847 out.n4737 0.001
R88036 out.n4706 out.n4705 0.001
R88037 out.n4850 out.n4699 0.001
R88038 out.n4853 out.n4673 0.001
R88039 out.n4644 out.n4643 0.001
R88040 out.n4856 out.n4637 0.001
R88041 out.n4859 out.n4609 0.001
R88042 out.n4861 out.n4570 0.001
R88043 out.n4572 out.n4571 0.001
R88044 out.n4864 out.n4541 0.001
R88045 out.n4514 out.n4513 0.001
R88046 out.n4867 out.n4506 0.001
R88047 out.n4508 out.n4507 0.001
R88048 out.n4870 out.n4478 0.001
R88049 out.n4450 out.n4449 0.001
R88050 out.n4872 out.n4441 0.001
R88051 out.n4443 out.n4442 0.001
R88052 out.n4875 out.n4414 0.001
R88053 out.n4386 out.n4385 0.001
R88054 out.n4878 out.n4378 0.001
R88055 out.n4380 out.n4379 0.001
R88056 out.n4881 out.n4349 0.001
R88057 out.n4322 out.n4321 0.001
R88058 out.n4883 out.n4313 0.001
R88059 out.n4315 out.n4314 0.001
R88060 out.n4886 out.n4282 0.001
R88061 out.n4256 out.n4255 0.001
R88062 out.n4888 out.n4247 0.001
R88063 out.n4249 out.n4248 0.001
R88064 out.n4890 out.n4219 0.001
R88065 out.n4192 out.n4191 0.001
R88066 out.n4893 out.n4183 0.001
R88067 out.n4185 out.n4184 0.001
R88068 out.n4896 out.n4155 0.001
R88069 out.n4899 out.n4120 0.001
R88070 out.n4902 out.n4092 0.001
R88071 out.n4063 out.n4062 0.001
R88072 out.n4904 out.n4054 0.001
R88073 out.n4056 out.n4055 0.001
R88074 out.n4906 out.n4026 0.001
R88075 out.n8796 out.n4942 0.001
R88076 out.n8799 out.n919 0.001
R88077 out.n8802 out.n858 0.001
R88078 out.n860 out.n859 0.001
R88079 out.n8805 out.n828 0.001
R88080 out.n799 out.n798 0.001
R88081 out.n8808 out.n791 0.001
R88082 out.n793 out.n792 0.001
R88083 out.n8811 out.n768 0.001
R88084 out.n8814 out.n729 0.001
R88085 out.n8817 out.n705 0.001
R88086 out.n673 out.n672 0.001
R88087 out.n8819 out.n664 0.001
R88088 out.n666 out.n665 0.001
R88089 out.n8822 out.n638 0.001
R88090 out.n609 out.n608 0.001
R88091 out.n8825 out.n601 0.001
R88092 out.n603 out.n602 0.001
R88093 out.n8827 out.n572 0.001
R88094 out.n542 out.n541 0.001
R88095 out.n8830 out.n533 0.001
R88096 out.n535 out.n534 0.001
R88097 out.n8833 out.n511 0.001
R88098 out.n480 out.n479 0.001
R88099 out.n8836 out.n472 0.001
R88100 out.n474 out.n473 0.001
R88101 out.n8839 out.n444 0.001
R88102 out.n8842 out.n409 0.001
R88103 out.n8844 out.n381 0.001
R88104 out.n8846 out.n344 0.001
R88105 out.n8848 out.n313 0.001
R88106 out.n282 out.n281 0.001
R88107 out.n8851 out.n274 0.001
R88108 out.n8854 out.n251 0.001
R88109 out.n221 out.n220 0.001
R88110 out.n8857 out.n213 0.001
R88111 out.n215 out.n214 0.001
R88112 out.n8860 out.n185 0.001
R88113 out.n156 out.n155 0.001
R88114 out.n8863 out.n148 0.001
R88115 out.n150 out.n149 0.001
R88116 out.n8866 out.n119 0.001
R88117 out.n8869 out.n88 0.001
R88118 out.n8871 out.n56 0.001
R88119 out.n15 out.n14 0.001
R88120 out.n6741 out.n6738 0.001
R88121 out.n6737 out.n6735 0.001
R88122 out.n3230 out.n3229 0.001
R88123 out.n919 out.n911 0.001
R88124 out.n6283 out.n6279 0.001
R88125 out.n6403 out.n6400 0.001
R88126 out.n6399 out.n6397 0.001
R88127 out.n6065 out.n6062 0.001
R88128 out.n6061 out.n6059 0.001
R88129 out.n6170 out.n6167 0.001
R88130 out.n6188 out.n6185 0.001
R88131 out.n1622 out.n1621 0.001
R88132 out.n3087 out.n3086 0.001
R88133 out.n6194 out.n6193 0.001
R88134 out.n6840 out.n6836 0.001
R88135 out.n6965 out.n6962 0.001
R88136 out.n6961 out.n6959 0.001
R88137 out.n7445 out.n7442 0.001
R88138 out.n7441 out.n7439 0.001
R88139 out.n7102 out.n7098 0.001
R88140 out.n7215 out.n7212 0.001
R88141 out.n7211 out.n7209 0.001
R88142 out.n7687 out.n7683 0.001
R88143 out.n7786 out.n7783 0.001
R88144 out.n7782 out.n7780 0.001
R88145 out.n2722 out.n2721 0.001
R88146 out.n2618 out.n2617 0.001
R88147 out.n883 out.n882 0.001
R88148 out.n7000 out.n6999 0.001
R88149 out.n7012 out.n7011 0.001
R88150 out.n7820 out.n6767 0.001
R88151 out.n7847 out.n7846 0.001
R88152 out.n7859 out.n7845 0.001
R88153 out.n7887 out.n7886 0.001
R88154 out.n7897 out.n7885 0.001
R88155 out.n7924 out.n7923 0.001
R88156 out.n7936 out.n7922 0.001
R88157 out.n7964 out.n7963 0.001
R88158 out.n7974 out.n7962 0.001
R88159 out.n8001 out.n8000 0.001
R88160 out.n8013 out.n7999 0.001
R88161 out.n8041 out.n8040 0.001
R88162 out.n8051 out.n8039 0.001
R88163 out.n8078 out.n8077 0.001
R88164 out.n8090 out.n8076 0.001
R88165 out.n8118 out.n8117 0.001
R88166 out.n8128 out.n8116 0.001
R88167 out.n8155 out.n8154 0.001
R88168 out.n8167 out.n8153 0.001
R88169 out.n8195 out.n8194 0.001
R88170 out.n8205 out.n8193 0.001
R88171 out.n8232 out.n8231 0.001
R88172 out.n8244 out.n8230 0.001
R88173 out.n8272 out.n8271 0.001
R88174 out.n8282 out.n8270 0.001
R88175 out.n8309 out.n8308 0.001
R88176 out.n8321 out.n8307 0.001
R88177 out.n8349 out.n8348 0.001
R88178 out.n8359 out.n8347 0.001
R88179 out.n8386 out.n8385 0.001
R88180 out.n8398 out.n8384 0.001
R88181 out.n8426 out.n8425 0.001
R88182 out.n8436 out.n8424 0.001
R88183 out.n8463 out.n8462 0.001
R88184 out.n8475 out.n8461 0.001
R88185 out.n8503 out.n8502 0.001
R88186 out.n8513 out.n8501 0.001
R88187 out.n8540 out.n8539 0.001
R88188 out.n8552 out.n8538 0.001
R88189 out.n8580 out.n8579 0.001
R88190 out.n8590 out.n8578 0.001
R88191 out.n8617 out.n8616 0.001
R88192 out.n8629 out.n8615 0.001
R88193 out.n8657 out.n8656 0.001
R88194 out.n8667 out.n8655 0.001
R88195 out.n8694 out.n8693 0.001
R88196 out.n8706 out.n8692 0.001
R88197 out.n8734 out.n8733 0.001
R88198 out.n8744 out.n8732 0.001
R88199 out.n8777 out.n8776 0.001
R88200 out.n8792 out.n8775 0.001
R88201 out.n886 out.n885 0.001
R88202 out.n899 out.n898 0.001
R88203 out.n3961 out.n3948 0.001
R88204 out.n3937 out.n3936 0.001
R88205 out.n3923 out.n3910 0.001
R88206 out.n3899 out.n3898 0.001
R88207 out.n3884 out.n3871 0.001
R88208 out.n3860 out.n3859 0.001
R88209 out.n3846 out.n3833 0.001
R88210 out.n3822 out.n3821 0.001
R88211 out.n3807 out.n3794 0.001
R88212 out.n3783 out.n3782 0.001
R88213 out.n3769 out.n3756 0.001
R88214 out.n3745 out.n3744 0.001
R88215 out.n3730 out.n3717 0.001
R88216 out.n3706 out.n3705 0.001
R88217 out.n3692 out.n3679 0.001
R88218 out.n3668 out.n3667 0.001
R88219 out.n3653 out.n3640 0.001
R88220 out.n3629 out.n3628 0.001
R88221 out.n3615 out.n3602 0.001
R88222 out.n3591 out.n3590 0.001
R88223 out.n3576 out.n3563 0.001
R88224 out.n3552 out.n3551 0.001
R88225 out.n3538 out.n3525 0.001
R88226 out.n3514 out.n3513 0.001
R88227 out.n3499 out.n3486 0.001
R88228 out.n3475 out.n3474 0.001
R88229 out.n3461 out.n3448 0.001
R88230 out.n3437 out.n3436 0.001
R88231 out.n3422 out.n3409 0.001
R88232 out.n3398 out.n3397 0.001
R88233 out.n3384 out.n3371 0.001
R88234 out.n3360 out.n3359 0.001
R88235 out.n3345 out.n3332 0.001
R88236 out.n3321 out.n3320 0.001
R88237 out.n3307 out.n3294 0.001
R88238 out.n3283 out.n3282 0.001
R88239 out.n3268 out.n3238 0.001
R88240 out.n3207 out.n3206 0.001
R88241 out.n3214 out.n3213 0.001
R88242 out.n3123 out.n3122 0.001
R88243 out.n3150 out.n3121 0.001
R88244 out.n3091 out.n3090 0.001
R88245 out.n3070 out.n3057 0.001
R88246 out.n3046 out.n3045 0.001
R88247 out.n3023 out.n2996 0.001
R88248 out.n2976 out.n2975 0.001
R88249 out.n2184 out.n2183 0.001
R88250 out.n2943 out.n2180 0.001
R88251 out.n1633 out.n1632 0.001
R88252 out.n1630 out.n1629 0.001
R88253 out.n1849 out.n1848 0.001
R88254 out.n1617 out.n1616 0.001
R88255 out.n6444 out.n6443 0.001
R88256 out.n6449 out.n6448 0.001
R88257 out.n6767 out.n6766 0.001
R88258 out.n7843 out.n7842 0.001
R88259 out.n7845 out.n7844 0.001
R88260 out.n7881 out.n7880 0.001
R88261 out.n7885 out.n7884 0.001
R88262 out.n7920 out.n7919 0.001
R88263 out.n7922 out.n7921 0.001
R88264 out.n7958 out.n7957 0.001
R88265 out.n7962 out.n7961 0.001
R88266 out.n7997 out.n7996 0.001
R88267 out.n7999 out.n7998 0.001
R88268 out.n8035 out.n8034 0.001
R88269 out.n8039 out.n8038 0.001
R88270 out.n8074 out.n8073 0.001
R88271 out.n8076 out.n8075 0.001
R88272 out.n8112 out.n8111 0.001
R88273 out.n8116 out.n8115 0.001
R88274 out.n8151 out.n8150 0.001
R88275 out.n8153 out.n8152 0.001
R88276 out.n8189 out.n8188 0.001
R88277 out.n8193 out.n8192 0.001
R88278 out.n8228 out.n8227 0.001
R88279 out.n8230 out.n8229 0.001
R88280 out.n8266 out.n8265 0.001
R88281 out.n8270 out.n8269 0.001
R88282 out.n8305 out.n8304 0.001
R88283 out.n8307 out.n8306 0.001
R88284 out.n8343 out.n8342 0.001
R88285 out.n8347 out.n8346 0.001
R88286 out.n8382 out.n8381 0.001
R88287 out.n8384 out.n8383 0.001
R88288 out.n8420 out.n8419 0.001
R88289 out.n8424 out.n8423 0.001
R88290 out.n8459 out.n8458 0.001
R88291 out.n8461 out.n8460 0.001
R88292 out.n8497 out.n8496 0.001
R88293 out.n8501 out.n8500 0.001
R88294 out.n8536 out.n8535 0.001
R88295 out.n8538 out.n8537 0.001
R88296 out.n8574 out.n8573 0.001
R88297 out.n8578 out.n8577 0.001
R88298 out.n8613 out.n8612 0.001
R88299 out.n8615 out.n8614 0.001
R88300 out.n8651 out.n8650 0.001
R88301 out.n8655 out.n8654 0.001
R88302 out.n8690 out.n8689 0.001
R88303 out.n8692 out.n8691 0.001
R88304 out.n8728 out.n8727 0.001
R88305 out.n8732 out.n8731 0.001
R88306 out.n8771 out.n8770 0.001
R88307 out.n8775 out.n8774 0.001
R88308 out.n4933 out.n4932 0.001
R88309 out.n910 out.n907 0.001
R88310 out.n906 out.n905 0.001
R88311 out.n3948 out.n3945 0.001
R88312 out.n3947 out.n3946 0.001
R88313 out.n3910 out.n3907 0.001
R88314 out.n3909 out.n3908 0.001
R88315 out.n3871 out.n3868 0.001
R88316 out.n3870 out.n3869 0.001
R88317 out.n3833 out.n3830 0.001
R88318 out.n3832 out.n3831 0.001
R88319 out.n3794 out.n3791 0.001
R88320 out.n3793 out.n3792 0.001
R88321 out.n3756 out.n3753 0.001
R88322 out.n3755 out.n3754 0.001
R88323 out.n3717 out.n3714 0.001
R88324 out.n3716 out.n3715 0.001
R88325 out.n3679 out.n3676 0.001
R88326 out.n3678 out.n3677 0.001
R88327 out.n3640 out.n3637 0.001
R88328 out.n3639 out.n3638 0.001
R88329 out.n3602 out.n3599 0.001
R88330 out.n3601 out.n3600 0.001
R88331 out.n3563 out.n3560 0.001
R88332 out.n3562 out.n3561 0.001
R88333 out.n3525 out.n3522 0.001
R88334 out.n3524 out.n3523 0.001
R88335 out.n3486 out.n3483 0.001
R88336 out.n3485 out.n3484 0.001
R88337 out.n3448 out.n3445 0.001
R88338 out.n3447 out.n3446 0.001
R88339 out.n3409 out.n3406 0.001
R88340 out.n3408 out.n3407 0.001
R88341 out.n3371 out.n3368 0.001
R88342 out.n3370 out.n3369 0.001
R88343 out.n3332 out.n3329 0.001
R88344 out.n3331 out.n3330 0.001
R88345 out.n3294 out.n3291 0.001
R88346 out.n3293 out.n3292 0.001
R88347 out.n3238 out.n3233 0.001
R88348 out.n3237 out.n3236 0.001
R88349 out.n3111 out.n3110 0.001
R88350 out.n3113 out.n3109 0.001
R88351 out.n3104 out.n3103 0.001
R88352 out.n3121 out.n3118 0.001
R88353 out.n3120 out.n3119 0.001
R88354 out.n3057 out.n3054 0.001
R88355 out.n3056 out.n3055 0.001
R88356 out.n2996 out.n2991 0.001
R88357 out.n2995 out.n2994 0.001
R88358 out.n2072 out.n2071 0.001
R88359 out.n2180 out.n2172 0.001
R88360 out.n2179 out.n2178 0.001
R88361 out.n2176 out.n2175 0.001
R88362 out.n7242 out.n7241 0.001
R88363 out.n2957 out.n1134 0.001
R88364 out.n5612 out.n5611 0.001
R88365 out.n5617 out.n5616 0.001
R88366 out.n7824 out.n7823 0.001
R88367 out.n7828 out.n7827 0.001
R88368 out.n7863 out.n7862 0.001
R88369 out.n7868 out.n7867 0.001
R88370 out.n7901 out.n7900 0.001
R88371 out.n7905 out.n7904 0.001
R88372 out.n7940 out.n7939 0.001
R88373 out.n7945 out.n7944 0.001
R88374 out.n7978 out.n7977 0.001
R88375 out.n7982 out.n7981 0.001
R88376 out.n8017 out.n8016 0.001
R88377 out.n8022 out.n8021 0.001
R88378 out.n8055 out.n8054 0.001
R88379 out.n8059 out.n8058 0.001
R88380 out.n8094 out.n8093 0.001
R88381 out.n8099 out.n8098 0.001
R88382 out.n8132 out.n8131 0.001
R88383 out.n8136 out.n8135 0.001
R88384 out.n8171 out.n8170 0.001
R88385 out.n8176 out.n8175 0.001
R88386 out.n8209 out.n8208 0.001
R88387 out.n8213 out.n8212 0.001
R88388 out.n8248 out.n8247 0.001
R88389 out.n8253 out.n8252 0.001
R88390 out.n8286 out.n8285 0.001
R88391 out.n8290 out.n8289 0.001
R88392 out.n8325 out.n8324 0.001
R88393 out.n8330 out.n8329 0.001
R88394 out.n8363 out.n8362 0.001
R88395 out.n8367 out.n8366 0.001
R88396 out.n8402 out.n8401 0.001
R88397 out.n8407 out.n8406 0.001
R88398 out.n8440 out.n8439 0.001
R88399 out.n8444 out.n8443 0.001
R88400 out.n8479 out.n8478 0.001
R88401 out.n8484 out.n8483 0.001
R88402 out.n8517 out.n8516 0.001
R88403 out.n8521 out.n8520 0.001
R88404 out.n8556 out.n8555 0.001
R88405 out.n8561 out.n8560 0.001
R88406 out.n8594 out.n8593 0.001
R88407 out.n8598 out.n8597 0.001
R88408 out.n8633 out.n8632 0.001
R88409 out.n8638 out.n8637 0.001
R88410 out.n8671 out.n8670 0.001
R88411 out.n8675 out.n8674 0.001
R88412 out.n8710 out.n8709 0.001
R88413 out.n8715 out.n8714 0.001
R88414 out.n8748 out.n8747 0.001
R88415 out.n8752 out.n8751 0.001
R88416 out.n8796 out.n8794 0.001
R88417 out.n865 out.n864 0.001
R88418 out.n864 out.n863 0.001
R88419 out.n3991 out.n3988 0.001
R88420 out.n3990 out.n3989 0.001
R88421 out.n3968 out.n3965 0.001
R88422 out.n3967 out.n3966 0.001
R88423 out.n3930 out.n3927 0.001
R88424 out.n3929 out.n3928 0.001
R88425 out.n3891 out.n3888 0.001
R88426 out.n3890 out.n3889 0.001
R88427 out.n3853 out.n3850 0.001
R88428 out.n3852 out.n3851 0.001
R88429 out.n3814 out.n3811 0.001
R88430 out.n3813 out.n3812 0.001
R88431 out.n3776 out.n3773 0.001
R88432 out.n3775 out.n3774 0.001
R88433 out.n3737 out.n3734 0.001
R88434 out.n3736 out.n3735 0.001
R88435 out.n3699 out.n3696 0.001
R88436 out.n3698 out.n3697 0.001
R88437 out.n3660 out.n3657 0.001
R88438 out.n3659 out.n3658 0.001
R88439 out.n3622 out.n3619 0.001
R88440 out.n3621 out.n3620 0.001
R88441 out.n3583 out.n3580 0.001
R88442 out.n3582 out.n3581 0.001
R88443 out.n3545 out.n3542 0.001
R88444 out.n3544 out.n3543 0.001
R88445 out.n3506 out.n3503 0.001
R88446 out.n3505 out.n3504 0.001
R88447 out.n3468 out.n3465 0.001
R88448 out.n3467 out.n3466 0.001
R88449 out.n3429 out.n3426 0.001
R88450 out.n3428 out.n3427 0.001
R88451 out.n3391 out.n3388 0.001
R88452 out.n3390 out.n3389 0.001
R88453 out.n3352 out.n3349 0.001
R88454 out.n3351 out.n3350 0.001
R88455 out.n3314 out.n3311 0.001
R88456 out.n3313 out.n3312 0.001
R88457 out.n3275 out.n3272 0.001
R88458 out.n3274 out.n3273 0.001
R88459 out.n3198 out.n3195 0.001
R88460 out.n3197 out.n3196 0.001
R88461 out.n3183 out.n3180 0.001
R88462 out.n3182 out.n3181 0.001
R88463 out.n3157 out.n3154 0.001
R88464 out.n3156 out.n3155 0.001
R88465 out.n3077 out.n3074 0.001
R88466 out.n3076 out.n3075 0.001
R88467 out.n3039 out.n3031 0.001
R88468 out.n1138 out.n1137 0.001
R88469 out.n2957 out.n2952 0.001
R88470 out.n878 out.n877 0.001
R88471 out.n3195 out.n3194 0.001
R88472 out.n5626 out.n5625 0.001
R88473 out.n5865 out.n5864 0.001
R88474 out.n7821 out.n7820 0.001
R88475 out.n7832 out.n7831 0.001
R88476 out.n7860 out.n7859 0.001
R88477 out.n7872 out.n7871 0.001
R88478 out.n7898 out.n7897 0.001
R88479 out.n7909 out.n7908 0.001
R88480 out.n7937 out.n7936 0.001
R88481 out.n7949 out.n7948 0.001
R88482 out.n7975 out.n7974 0.001
R88483 out.n7986 out.n7985 0.001
R88484 out.n8014 out.n8013 0.001
R88485 out.n8026 out.n8025 0.001
R88486 out.n8052 out.n8051 0.001
R88487 out.n8063 out.n8062 0.001
R88488 out.n8091 out.n8090 0.001
R88489 out.n8103 out.n8102 0.001
R88490 out.n8129 out.n8128 0.001
R88491 out.n8140 out.n8139 0.001
R88492 out.n8168 out.n8167 0.001
R88493 out.n8180 out.n8179 0.001
R88494 out.n8206 out.n8205 0.001
R88495 out.n8217 out.n8216 0.001
R88496 out.n8245 out.n8244 0.001
R88497 out.n8257 out.n8256 0.001
R88498 out.n8283 out.n8282 0.001
R88499 out.n8294 out.n8293 0.001
R88500 out.n8322 out.n8321 0.001
R88501 out.n8334 out.n8333 0.001
R88502 out.n8360 out.n8359 0.001
R88503 out.n8371 out.n8370 0.001
R88504 out.n8399 out.n8398 0.001
R88505 out.n8411 out.n8410 0.001
R88506 out.n8437 out.n8436 0.001
R88507 out.n8448 out.n8447 0.001
R88508 out.n8476 out.n8475 0.001
R88509 out.n8488 out.n8487 0.001
R88510 out.n8514 out.n8513 0.001
R88511 out.n8525 out.n8524 0.001
R88512 out.n8553 out.n8552 0.001
R88513 out.n8565 out.n8564 0.001
R88514 out.n8591 out.n8590 0.001
R88515 out.n8602 out.n8601 0.001
R88516 out.n8630 out.n8629 0.001
R88517 out.n8642 out.n8641 0.001
R88518 out.n8668 out.n8667 0.001
R88519 out.n8679 out.n8678 0.001
R88520 out.n8707 out.n8706 0.001
R88521 out.n8719 out.n8718 0.001
R88522 out.n8745 out.n8744 0.001
R88523 out.n8758 out.n8757 0.001
R88524 out.n8793 out.n8792 0.001
R88525 out.n880 out.n879 0.001
R88526 out.n3985 out.n3984 0.001
R88527 out.n3978 out.n3977 0.001
R88528 out.n3962 out.n3961 0.001
R88529 out.n3955 out.n3954 0.001
R88530 out.n3924 out.n3923 0.001
R88531 out.n3917 out.n3916 0.001
R88532 out.n3885 out.n3884 0.001
R88533 out.n3878 out.n3877 0.001
R88534 out.n3847 out.n3846 0.001
R88535 out.n3840 out.n3839 0.001
R88536 out.n3808 out.n3807 0.001
R88537 out.n3801 out.n3800 0.001
R88538 out.n3770 out.n3769 0.001
R88539 out.n3763 out.n3762 0.001
R88540 out.n3731 out.n3730 0.001
R88541 out.n3724 out.n3723 0.001
R88542 out.n3693 out.n3692 0.001
R88543 out.n3686 out.n3685 0.001
R88544 out.n3654 out.n3653 0.001
R88545 out.n3647 out.n3646 0.001
R88546 out.n3616 out.n3615 0.001
R88547 out.n3609 out.n3608 0.001
R88548 out.n3577 out.n3576 0.001
R88549 out.n3570 out.n3569 0.001
R88550 out.n3539 out.n3538 0.001
R88551 out.n3532 out.n3531 0.001
R88552 out.n3500 out.n3499 0.001
R88553 out.n3493 out.n3492 0.001
R88554 out.n3462 out.n3461 0.001
R88555 out.n3455 out.n3454 0.001
R88556 out.n3423 out.n3422 0.001
R88557 out.n3416 out.n3415 0.001
R88558 out.n3385 out.n3384 0.001
R88559 out.n3378 out.n3377 0.001
R88560 out.n3346 out.n3345 0.001
R88561 out.n3339 out.n3338 0.001
R88562 out.n3308 out.n3307 0.001
R88563 out.n3301 out.n3300 0.001
R88564 out.n3269 out.n3268 0.001
R88565 out.n3260 out.n3259 0.001
R88566 out.n3167 out.n3166 0.001
R88567 out.n3177 out.n3176 0.001
R88568 out.n3170 out.n3169 0.001
R88569 out.n3151 out.n3150 0.001
R88570 out.n3140 out.n3139 0.001
R88571 out.n3071 out.n3070 0.001
R88572 out.n3064 out.n3063 0.001
R88573 out.n3024 out.n3023 0.001
R88574 out.n3012 out.n3011 0.001
R88575 out.n1537 out.n1536 0.001
R88576 out.n2944 out.n2943 0.001
R88577 out.n2614 out.n2613 0.001
R88578 out.n2611 out.n2610 0.001
R88579 out.n2727 out.n2726 0.001
R88580 out.n10292 out.n10291 0.001
R88581 out.n10294 out.n10293 0.001
R88582 out.n15199 out.n15166 0.001
R88583 out.n16268 out.n16266 0.001
R88584 out.n16200 out.n16199 0.001
R88585 out.n15903 out.n15902 0.001
R88586 out.n15562 out.n15561 0.001
R88587 out.n11977 out.n11976 0.001
R88588 out.n3233 out.n3232 0.001
R88589 out.n8774 out.n8773 0.001
R88590 out.n6766 out.n6765 0.001
R88591 out.n3113 out.n3112 0.001
R88592 out.n2991 out.n2990 0.001
R88593 out.n2172 out.n2075 0.001
R88594 out.n2172 out.n2171 0.001
R88595 out.n9052 out.n9044 0.001
R88596 out.n9423 out.n9412 0.001
R88597 out.n8872 out.n8871 0.001
R88598 out.n10016 out.n10015 0.001
R88599 out.n9544 out.n9543 0.001
R88600 out.n9543 out.n9510 0.001
R88601 out.n9580 out.n9579 0.001
R88602 out.n9579 out.n9546 0.001
R88603 out.n9616 out.n9615 0.001
R88604 out.n9615 out.n9582 0.001
R88605 out.n9674 out.n9619 0.001
R88606 out.n9675 out.n9674 0.001
R88607 out.n9711 out.n9710 0.001
R88608 out.n9710 out.n9677 0.001
R88609 out.n9747 out.n9746 0.001
R88610 out.n9746 out.n9713 0.001
R88611 out.n9783 out.n9782 0.001
R88612 out.n9782 out.n9749 0.001
R88613 out.n9819 out.n9818 0.001
R88614 out.n9818 out.n9785 0.001
R88615 out.n9855 out.n9854 0.001
R88616 out.n9854 out.n9821 0.001
R88617 out.n9891 out.n9858 0.001
R88618 out.n9925 out.n9892 0.001
R88619 out.n9962 out.n9961 0.001
R88620 out.n9961 out.n9926 0.001
R88621 out.n9998 out.n9997 0.001
R88622 out.n9997 out.n9964 0.001
R88623 out.n17307 out.n10001 0.001
R88624 out.n17307 out.n17239 0.001
R88625 out.n17236 out.n17235 0.001
R88626 out.n17237 out.n17236 0.001
R88627 out.n17232 out.n17231 0.001
R88628 out.n17233 out.n17232 0.001
R88629 out.n17228 out.n17227 0.001
R88630 out.n17229 out.n17228 0.001
R88631 out.n17224 out.n17223 0.001
R88632 out.n17225 out.n17224 0.001
R88633 out.n17220 out.n17219 0.001
R88634 out.n17221 out.n17220 0.001
R88635 out.n17216 out.n17215 0.001
R88636 out.n17217 out.n17216 0.001
R88637 out.n17212 out.n17211 0.001
R88638 out.n17213 out.n17212 0.001
R88639 out.n17208 out.n17207 0.001
R88640 out.n17209 out.n17208 0.001
R88641 out.n17204 out.n17203 0.001
R88642 out.n17205 out.n17204 0.001
R88643 out.n17200 out.n17199 0.001
R88644 out.n17201 out.n17200 0.001
R88645 out.n17196 out.n17195 0.001
R88646 out.n17197 out.n17196 0.001
R88647 out.n17192 out.n17191 0.001
R88648 out.n17193 out.n17192 0.001
R88649 out.n17188 out.n17187 0.001
R88650 out.n17189 out.n17188 0.001
R88651 out.n3146 out.n3145 0.001
R88652 out.n4835 out.n4823 0.001
R88653 out.n4763 out.n4752 0.001
R88654 out.n4699 out.n4689 0.001
R88655 out.n4637 out.n4627 0.001
R88656 out.n4570 out.n4559 0.001
R88657 out.n4506 out.n4494 0.001
R88658 out.n4441 out.n4432 0.001
R88659 out.n4378 out.n4367 0.001
R88660 out.n4313 out.n4299 0.001
R88661 out.n4247 out.n4237 0.001
R88662 out.n4183 out.n4174 0.001
R88663 out.n4120 out.n4111 0.001
R88664 out.n4054 out.n4044 0.001
R88665 out.n4942 out.n4931 0.001
R88666 out.n858 out.n845 0.001
R88667 out.n791 out.n781 0.001
R88668 out.n729 out.n721 0.001
R88669 out.n664 out.n654 0.001
R88670 out.n601 out.n589 0.001
R88671 out.n533 out.n522 0.001
R88672 out.n472 out.n461 0.001
R88673 out.n409 out.n399 0.001
R88674 out.n344 out.n333 0.001
R88675 out.n274 out.n264 0.001
R88676 out.n213 out.n202 0.001
R88677 out.n148 out.n137 0.001
R88678 out.n88 out.n77 0.001
R88679 out.n2074 out.n2073 0.001
R88680 out.n2960 out.n2957 0.001
R88681 out.n9508 out.n9507 0.001
R88682 out.n9509 out.n9508 0.001
R88683 out.n8871 out.n8870 0.001
R88684 out.n8868 out.n8866 0.001
R88685 out.n8866 out.n8865 0.001
R88686 out.n8862 out.n8860 0.001
R88687 out.n8860 out.n8859 0.001
R88688 out.n8856 out.n8854 0.001
R88689 out.n8854 out.n8853 0.001
R88690 out.n8850 out.n8848 0.001
R88691 out.n8848 out.n8847 0.001
R88692 out.n8845 out.n8844 0.001
R88693 out.n8844 out.n8843 0.001
R88694 out.n8841 out.n8839 0.001
R88695 out.n8839 out.n8838 0.001
R88696 out.n8835 out.n8833 0.001
R88697 out.n8833 out.n8832 0.001
R88698 out.n8829 out.n8827 0.001
R88699 out.n8827 out.n8826 0.001
R88700 out.n8824 out.n8822 0.001
R88701 out.n8822 out.n8821 0.001
R88702 out.n8818 out.n8817 0.001
R88703 out.n8817 out.n8816 0.001
R88704 out.n8813 out.n8811 0.001
R88705 out.n8811 out.n8810 0.001
R88706 out.n8807 out.n8805 0.001
R88707 out.n8805 out.n8804 0.001
R88708 out.n8801 out.n8799 0.001
R88709 out.n8798 out.n8796 0.001
R88710 out.n4908 out.n4906 0.001
R88711 out.n4906 out.n4905 0.001
R88712 out.n4903 out.n4902 0.001
R88713 out.n4902 out.n4901 0.001
R88714 out.n4898 out.n4896 0.001
R88715 out.n4896 out.n4895 0.001
R88716 out.n4892 out.n4890 0.001
R88717 out.n4890 out.n4889 0.001
R88718 out.n4887 out.n4886 0.001
R88719 out.n4886 out.n4885 0.001
R88720 out.n4882 out.n4881 0.001
R88721 out.n4881 out.n4880 0.001
R88722 out.n4877 out.n4875 0.001
R88723 out.n4875 out.n4874 0.001
R88724 out.n4871 out.n4870 0.001
R88725 out.n4870 out.n4869 0.001
R88726 out.n4866 out.n4864 0.001
R88727 out.n4864 out.n4863 0.001
R88728 out.n4860 out.n4859 0.001
R88729 out.n4859 out.n4858 0.001
R88730 out.n4855 out.n4853 0.001
R88731 out.n4853 out.n4852 0.001
R88732 out.n4849 out.n4847 0.001
R88733 out.n4847 out.n4846 0.001
R88734 out.n4843 out.n4841 0.001
R88735 out.n4841 out.n4840 0.001
R88736 out.n4840 out.n4838 0.001
R88737 out.n4844 out.n4843 0.001
R88738 out.n4846 out.n4844 0.001
R88739 out.n4850 out.n4849 0.001
R88740 out.n4852 out.n4850 0.001
R88741 out.n4856 out.n4855 0.001
R88742 out.n4858 out.n4856 0.001
R88743 out.n4861 out.n4860 0.001
R88744 out.n4863 out.n4861 0.001
R88745 out.n4867 out.n4866 0.001
R88746 out.n4869 out.n4867 0.001
R88747 out.n4872 out.n4871 0.001
R88748 out.n4874 out.n4872 0.001
R88749 out.n4878 out.n4877 0.001
R88750 out.n4880 out.n4878 0.001
R88751 out.n4883 out.n4882 0.001
R88752 out.n4885 out.n4883 0.001
R88753 out.n4888 out.n4887 0.001
R88754 out.n4889 out.n4888 0.001
R88755 out.n4893 out.n4892 0.001
R88756 out.n4895 out.n4893 0.001
R88757 out.n4899 out.n4898 0.001
R88758 out.n4901 out.n4899 0.001
R88759 out.n4904 out.n4903 0.001
R88760 out.n4905 out.n4904 0.001
R88761 out.n8796 out.n4908 0.001
R88762 out.n8799 out.n8798 0.001
R88763 out.n8802 out.n8801 0.001
R88764 out.n8804 out.n8802 0.001
R88765 out.n8808 out.n8807 0.001
R88766 out.n8810 out.n8808 0.001
R88767 out.n8814 out.n8813 0.001
R88768 out.n8816 out.n8814 0.001
R88769 out.n8819 out.n8818 0.001
R88770 out.n8821 out.n8819 0.001
R88771 out.n8825 out.n8824 0.001
R88772 out.n8826 out.n8825 0.001
R88773 out.n8830 out.n8829 0.001
R88774 out.n8832 out.n8830 0.001
R88775 out.n8836 out.n8835 0.001
R88776 out.n8838 out.n8836 0.001
R88777 out.n8842 out.n8841 0.001
R88778 out.n8843 out.n8842 0.001
R88779 out.n8846 out.n8845 0.001
R88780 out.n8847 out.n8846 0.001
R88781 out.n8851 out.n8850 0.001
R88782 out.n8853 out.n8851 0.001
R88783 out.n8857 out.n8856 0.001
R88784 out.n8859 out.n8857 0.001
R88785 out.n8863 out.n8862 0.001
R88786 out.n8865 out.n8863 0.001
R88787 out.n8869 out.n8868 0.001
R88788 out.n8870 out.n8869 0.001
R88789 out.n2 out.n0 0.001
R88790 ldomc_0.otaldom_0.pcascodeupm_0.o1.n27 ldomc_0.otaldom_0.pcascodeupm_0.o1.t12 13.847
R88791 ldomc_0.otaldom_0.pcascodeupm_0.o1.n27 ldomc_0.otaldom_0.pcascodeupm_0.o1.t14 13.847
R88792 ldomc_0.otaldom_0.pcascodeupm_0.o1.n21 ldomc_0.otaldom_0.pcascodeupm_0.o1.t11 13.847
R88793 ldomc_0.otaldom_0.pcascodeupm_0.o1.n21 ldomc_0.otaldom_0.pcascodeupm_0.o1.t10 13.847
R88794 ldomc_0.otaldom_0.pcascodeupm_0.o1.n32 ldomc_0.otaldom_0.pcascodeupm_0.o1.t13 13.847
R88795 ldomc_0.otaldom_0.pcascodeupm_0.o1.n32 ldomc_0.otaldom_0.pcascodeupm_0.o1.t9 13.847
R88796 ldomc_0.otaldom_0.pcascodeupm_0.o1.n31 ldomc_0.otaldom_0.pcascodeupm_0.o1.t8 13.847
R88797 ldomc_0.otaldom_0.pcascodeupm_0.o1.n31 ldomc_0.otaldom_0.pcascodeupm_0.o1.t15 13.847
R88798 ldomc_0.otaldom_0.pcascodeupm_0.o1.n39 ldomc_0.otaldom_0.pcascodeupm_0.o1.t2 13.847
R88799 ldomc_0.otaldom_0.pcascodeupm_0.o1.n39 ldomc_0.otaldom_0.pcascodeupm_0.o1.t0 13.847
R88800 ldomc_0.otaldom_0.pcascodeupm_0.o1.n16 ldomc_0.otaldom_0.pcascodeupm_0.o1.t5 13.847
R88801 ldomc_0.otaldom_0.pcascodeupm_0.o1.n16 ldomc_0.otaldom_0.pcascodeupm_0.o1.t3 13.847
R88802 ldomc_0.otaldom_0.pcascodeupm_0.o1.n8 ldomc_0.otaldom_0.pcascodeupm_0.o1.t4 13.847
R88803 ldomc_0.otaldom_0.pcascodeupm_0.o1.n8 ldomc_0.otaldom_0.pcascodeupm_0.o1.t1 13.847
R88804 ldomc_0.otaldom_0.pcascodeupm_0.o1.n34 ldomc_0.otaldom_0.pcascodeupm_0.o1.t6 13.847
R88805 ldomc_0.otaldom_0.pcascodeupm_0.o1.n34 ldomc_0.otaldom_0.pcascodeupm_0.o1.t7 13.847
R88806 ldomc_0.otaldom_0.pcascodeupm_0.o1.n1 ldomc_0.otaldom_0.pcascodeupm_0.o1.n31 10.814
R88807 ldomc_0.otaldom_0.pcascodeupm_0.o1.n0 ldomc_0.otaldom_0.pcascodeupm_0.o1.n8 6.881
R88808 ldomc_0.otaldom_0.pcascodeupm_0.o1.n5 ldomc_0.otaldom_0.pcascodeupm_0.o1.n27 6.881
R88809 ldomc_0.otaldom_0.pcascodeupm_0.o1.n10 ldomc_0.otaldom_0.pcascodeupm_0.o1.n21 6.881
R88810 ldomc_0.otaldom_0.pcascodeupm_0.o1.n17 ldomc_0.otaldom_0.pcascodeupm_0.o1.n16 5.76
R88811 ldomc_0.otaldom_0.pcascodeupm_0.o1.n2 ldomc_0.otaldom_0.pcascodeupm_0.o1.n24 5.698
R88812 ldomc_0.otaldom_0.pcascodeupm_0.o1.n29 ldomc_0.otaldom_0.pcascodeupm_0.o1.n28 5.646
R88813 ldomc_0.otaldom_0.pcascodeupm_0.o1.n20 ldomc_0.otaldom_0.pcascodeupm_0.o1.n19 5.646
R88814 ldomc_0.otaldom_0.pcascodeupm_0.o1.n40 ldomc_0.otaldom_0.pcascodeupm_0.o1.n39 5.621
R88815 ldomc_0.otaldom_0.pcascodeupm_0.o1.n35 ldomc_0.otaldom_0.pcascodeupm_0.o1.n34 5.6
R88816 ldomc_0.otaldom_0.pcascodeupm_0.o1.n7 ldomc_0.otaldom_0.pcascodeupm_0.o1.n26 4.5
R88817 ldomc_0.otaldom_0.pcascodeupm_0.o1.n7 ldomc_0.otaldom_0.pcascodeupm_0.o1.n29 4.5
R88818 ldomc_0.otaldom_0.pcascodeupm_0.o1.n12 ldomc_0.otaldom_0.pcascodeupm_0.o1.n22 4.5
R88819 ldomc_0.otaldom_0.pcascodeupm_0.o1.n12 ldomc_0.otaldom_0.pcascodeupm_0.o1.n20 4.5
R88820 ldomc_0.otaldom_0.pcascodeupm_0.o1.n13 ldomc_0.otaldom_0.pcascodeupm_0.o1.n41 4.5
R88821 ldomc_0.otaldom_0.pcascodeupm_0.o1.n0 ldomc_0.otaldom_0.pcascodeupm_0.o1.n44 4.5
R88822 ldomc_0.otaldom_0.pcascodeupm_0.o1.n33 ldomc_0.otaldom_0.pcascodeupm_0.o1 3.616
R88823 ldomc_0.otaldom_0.pcascodeupm_0.o1.n4 ldomc_0.otaldom_0.pcascodeupm_0.o1.n15 3.03
R88824 ldomc_0.otaldom_0.pcascodeupm_0.o1.n2 ldomc_0.otaldom_0.pcascodeupm_0.o1.n25 2.252
R88825 ldomc_0.otaldom_0.pcascodeupm_0.o1.n3 ldomc_0.otaldom_0.pcascodeupm_0.o1.n7 2.25
R88826 ldomc_0.otaldom_0.pcascodeupm_0.o1.n3 ldomc_0.otaldom_0.pcascodeupm_0.o1.n30 2.25
R88827 ldomc_0.otaldom_0.pcascodeupm_0.o1.n0 ldomc_0.otaldom_0.pcascodeupm_0.o1.n43 2.182
R88828 ldomc_0.otaldom_0.pcascodeupm_0.o1.n45 ldomc_0.otaldom_0.pcascodeupm_0.o1.n42 2.039
R88829 ldomc_0.otaldom_0.pcascodeupm_0.o1.n35 ldomc_0.otaldom_0.pcascodeupm_0.o1.n33 1.377
R88830 ldomc_0.otaldom_0.pmoslm_0.o1 ldomc_0.otaldom_0.pcascodeupm_0.o1.n45 1.235
R88831 ldomc_0.otaldom_0.pcascodeupm_0.o1.n13 ldomc_0.otaldom_0.pcascodeupm_0.o1.n40 1.033
R88832 ldomc_0.otaldom_0.pcascodeupm_0.o1.n4 ldomc_0.otaldom_0.pcascodeupm_0.o1.n17 0.999
R88833 ldomc_0.otaldom_0.pmoslm_0.o1 ldomc_0.otaldom_0.pcascodeupm_0.o1.n37 0.89
R88834 ldomc_0.otaldom_0.pcascodeupm_0.o1.n24 ldomc_0.otaldom_0.pcascodeupm_0.o1.n23 0.866
R88835 ldomc_0.otaldom_0.pcascodeupm_0.o1.n42 ldomc_0.otaldom_0.pcascodeupm_0.o1.n13 0.865
R88836 ldomc_0.otaldom_0.pcascodeupm_0.o1.n37 ldomc_0.otaldom_0.pcascodeupm_0.o1.n4 0.766
R88837 ldomc_0.otaldom_0.pcascodeupm_0.o1.n33 ldomc_0.otaldom_0.pcascodeupm_0.o1.n3 0.668
R88838 ldomc_0.otaldom_0.pcascodeupm_0.o1.n13 ldomc_0.otaldom_0.pcascodeupm_0.o1.n38 0.613
R88839 ldomc_0.otaldom_0.pcascodeupm_0.o1.n23 ldomc_0.otaldom_0.pcascodeupm_0.o1.n18 0.613
R88840 ldomc_0.otaldom_0.pcascodeupm_0.o1.n23 ldomc_0.otaldom_0.pcascodeupm_0.o1.n12 0.589
R88841 ldomc_0.otaldom_0.pcascodeupm_0.o1.n36 ldomc_0.otaldom_0.pcascodeupm_0.o1.n35 0.344
R88842 ldomc_0.otaldom_0.pcascodeupm_0.o1.n12 ldomc_0.otaldom_0.pcascodeupm_0.o1.n9 0.171
R88843 ldomc_0.otaldom_0.pcascodeupm_0.o1.n12 ldomc_0.otaldom_0.pcascodeupm_0.o1.n11 0.133
R88844 ldomc_0.otaldom_0.pcascodeupm_0.o1.n1 ldomc_0.otaldom_0.pcascodeupm_0.o1.n32 5.124
R88845 ldomc_0.otaldom_0.pcascodeupm_0.o1.n4 ldomc_0.otaldom_0.pcascodeupm_0.o1.n14 0.626
R88846 ldomc_0.otaldom_0.pcascodeupm_0.o1.n7 ldomc_0.otaldom_0.pcascodeupm_0.o1.n5 0.135
R88847 ldomc_0.otaldom_0.pcascodeupm_0.o1.n3 ldomc_0.otaldom_0.pcascodeupm_0.o1.n2 0.127
R88848 ldomc_0.otaldom_0.pcascodeupm_0.o1.n12 ldomc_0.otaldom_0.pcascodeupm_0.o1.n10 0.11
R88849 ldomc_0.otaldom_0.pcascodeupm_0.o1.n7 ldomc_0.otaldom_0.pcascodeupm_0.o1.n6 0.108
R88850 ldomc_0.otaldom_0.pcascodeupm_0.o1.n37 ldomc_0.otaldom_0.pcascodeupm_0.o1.n36 0.097
R88851 ldomc_0.otaldom_0.pcascodeupm_0.o1 ldomc_0.otaldom_0.pcascodeupm_0.o1.n1 1.326
R88852 ldomc_0.otaldom_0.pcascodeupm_0.o1.n45 ldomc_0.otaldom_0.pcascodeupm_0.o1.n0 1.216
R88853 bandgapmd_0.otam_1.pdiffm_0.inp.n3 bandgapmd_0.otam_1.pdiffm_0.inp.t4 110.471
R88854 bandgapmd_0.otam_1.pdiffm_0.inp.n4 bandgapmd_0.otam_1.pdiffm_0.inp.t6 110.471
R88855 bandgapmd_0.otam_1.pdiffm_0.inp.n5 bandgapmd_0.otam_1.pdiffm_0.inp.t9 110.471
R88856 bandgapmd_0.otam_1.pdiffm_0.inp.n6 bandgapmd_0.otam_1.pdiffm_0.inp.t3 110.471
R88857 bandgapmd_0.otam_1.pdiffm_0.inp.n1 bandgapmd_0.otam_1.pdiffm_0.inp.t10 110.47
R88858 bandgapmd_0.otam_1.pdiffm_0.inp.n3 bandgapmd_0.otam_1.pdiffm_0.inp.t2 110.47
R88859 bandgapmd_0.otam_1.pdiffm_0.inp.n4 bandgapmd_0.otam_1.pdiffm_0.inp.t5 110.47
R88860 bandgapmd_0.otam_1.pdiffm_0.inp.n5 bandgapmd_0.otam_1.pdiffm_0.inp.t7 110.47
R88861 bandgapmd_0.otam_1.pdiffm_0.inp.n6 bandgapmd_0.otam_1.pdiffm_0.inp.t11 110.47
R88862 bandgapmd_0.otam_1.pdiffm_0.inp.n1 bandgapmd_0.otam_1.pdiffm_0.inp.t8 110.469
R88863 bandgapmd_0.otam_1.pdiffm_0.inp.n15 bandgapmd_0.otam_1.pdiffm_0.inp.n14 5.796
R88864 bandgapmd_0.otam_1.pdiffm_0.inp.n8 bandgapmd_0.otam_1.pdiffm_0.inp.n7 2.039
R88865 bandgapmd_0.otam_1.pdiffm_0.inp.n11 bandgapmd_0.otam_1.pdiffm_0.inp.n2 1.353
R88866 bandgapmd_0.otam_1.pdiffm_0.inp.n10 bandgapmd_0.otam_1.pdiffm_0.inp.n9 1.317
R88867 bandgapmd_0.otam_1.pdiffm_0.inp.n9 bandgapmd_0.otam_1.pdiffm_0.inp.n8 1.288
R88868 bandgapmd_0.otam_1.pdiffm_0.inp.n11 bandgapmd_0.otam_1.pdiffm_0.inp.n10 1.195
R88869 bandgapmd_0.otam_1.pdiffm_0.inp.n10 bandgapmd_0.otam_1.pdiffm_0.inp.n3 0.857
R88870 bandgapmd_0.otam_1.pdiffm_0.inp.n8 bandgapmd_0.otam_1.pdiffm_0.inp.n5 0.854
R88871 bandgapmd_0.otam_1.pdiffm_0.inp.n9 bandgapmd_0.otam_1.pdiffm_0.inp.n4 0.854
R88872 bandgapmd_0.bg_resm_0.vp bandgapmd_0.otam_1.pdiffm_0.inp.t0 0.425
R88873 bandgapmd_0.otam_1.pdiffm_0.inp.n2 bandgapmd_0.otam_1.pdiffm_0.inp.n1 0.139
R88874 bandgapmd_0.otam_1.pdiffm_0.inp.n7 bandgapmd_0.otam_1.pdiffm_0.inp 0.071
R88875 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.otam_1.pdiffm_0.inp.n6 0.066
R88876 bandgapmd_0.otam_1.pdiffm_0.inp.n12 bandgapmd_0.otam_1.pdiffm_0.inp.n11 0.022
R88877 bandgapmd_0.otam_1.pdiffm_0.inp.n14 bandgapmd_0.otam_1.pdiffm_0.inp.n13 0.019
R88878 bandgapmd_0.bg_resm_0.vp bandgapmd_0.otam_1.pdiffm_0.inp.n15 0.017
R88879 bandgapmd_0.otam_1.pdiffm_0.inp.n13 bandgapmd_0.otam_1.pdiffm_0.inp.n12 0.016
R88880 bandgapmd_0.otam_1.pdiffm_0.inp.n15 bandgapmd_0.bg_resm_0.vp 0.016
R88881 bandgapmd_0.otam_1.pdiffm_0.inp.n7 bandgapmd_0.otam_1.inp 0.008
R88882 bandgapmd_0.otam_1.pdiffm_0.inp.n14 bandgapmd_0.otam_1.pdiffm_0.inp.n0 0.001
R88883 bandgapmd_0.bg_stupm_0.vs2 bandgapmd_0.bg_stupm_0.vs2.t0 40.126
R88884 bandgapmd_0.bg_stupm_0.vs2 bandgapmd_0.bg_stupm_0.vs2.t1 40.123
R88885 bandgapmd_0.bg_pmosm_0.vbg.n67 bandgapmd_0.bg_pmosm_0.vbg.t9 110.493
R88886 bandgapmd_0.bg_pmosm_0.vbg.n55 bandgapmd_0.bg_pmosm_0.vbg.t10 110.492
R88887 bandgapmd_0.bg_pmosm_0.vbg.n44 bandgapmd_0.bg_pmosm_0.vbg.t11 110.49
R88888 bandgapmd_0.bg_pmosm_0.vbg.n52 bandgapmd_0.bg_pmosm_0.vbg.t3 110.489
R88889 bandgapmd_0.bg_pmosm_0.vbg.n62 bandgapmd_0.bg_pmosm_0.vbg.t12 110.488
R88890 bandgapmd_0.bg_pmosm_0.vbg.n60 bandgapmd_0.bg_pmosm_0.vbg.t8 110.485
R88891 bandgapmd_0.bg_pmosm_0.vbg.n50 bandgapmd_0.bg_pmosm_0.vbg.t14 110.484
R88892 bandgapmd_0.bg_pmosm_0.vbg.n47 bandgapmd_0.bg_pmosm_0.vbg.t4 110.483
R88893 bandgapmd_0.bg_pmosm_0.vbg.n57 bandgapmd_0.bg_pmosm_0.vbg.t6 110.481
R88894 bandgapmd_0.bg_pmosm_0.vbg.n65 bandgapmd_0.bg_pmosm_0.vbg.t13 110.48
R88895 bandgapmd_0.bg_pmosm_0.vbg.n35 bandgapmd_0.bg_pmosm_0.vbg.t5 37.358
R88896 bandgapmd_0.bg_pmosm_0.vbg.n19 bandgapmd_0.bg_pmosm_0.vbg.n18 22.445
R88897 bandgapmd_0.bg_pmosm_0.vbg.n10 bandgapmd_0.bg_pmosm_0.vbg.n9 12.759
R88898 bandgapmd_0.bg_pmosm_0.vbg.n37 bandgapmd_0.bg_pmosm_0.vbg.n36 10.617
R88899 bandgapmd_0.bg_pmosm_0.vbg.n13 bandgapmd_0.bg_pmosm_0.vbg.n6 10.285
R88900 bandgapmd_0.bg_pmosm_0.vbg.n20 bandgapmd_0.bg_pmosm_0.vbg.n19 9.3
R88901 bandgapmd_0.bg_pmosm_0.vbg.n19 bandgapmd_0.bg_pmosm_0.vbg.n3 9.3
R88902 bandgapmd_0.bg_pmosm_0.vbg.n11 bandgapmd_0.bg_pmosm_0.vbg.n5 9.3
R88903 bandgapmd_0.bg_pmosm_0.vbg.n17 bandgapmd_0.bg_pmosm_0.vbg.n10 9.122
R88904 bandgapmd_0.bg_pmosm_0.vbg.n16 bandgapmd_0.bg_pmosm_0.vbg.n13 7.106
R88905 bandgapmd_0.bg_pmosm_0.vbg.n17 bandgapmd_0.bg_pmosm_0.vbg.t0 6.923
R88906 bandgapmd_0.bg_pmosm_0.vbg.n17 bandgapmd_0.bg_pmosm_0.vbg.t1 6.923
R88907 bandgapmd_0.bg_pmosm_0.vbg.n36 bandgapmd_0.bg_pmosm_0.vbg.n33 5.571
R88908 bandgapmd_0.bg_pmosm_0.vbg.n69 bandgapmd_0.bg_pmosm_0.vbg.n68 5.461
R88909 bandgapmd_0.bg_pmosm_0.vbg.n30 bandgapmd_0.bg_pmosm_0.vbg.n0 4.5
R88910 bandgapmd_0.bg_pmosm_0.vbg.n28 bandgapmd_0.bg_pmosm_0.vbg.n27 4.5
R88911 bandgapmd_0.bg_pmosm_0.vbg.n26 bandgapmd_0.bg_pmosm_0.vbg.n21 4.5
R88912 bandgapmd_0.bg_pmosm_0.vbg.n22 bandgapmd_0.bg_pmosm_0.vbg.n4 4.5
R88913 bandgapmd_0.bg_pmosm_0.vbg.n23 bandgapmd_0.bg_pmosm_0.vbg.n2 4.5
R88914 bandgapmd_0.bg_pmosm_0.vbg.n32 bandgapmd_0.bg_pmosm_0.vbg.n31 4.5
R88915 bandgapmd_0.bg_pmosm_0.vbg.n17 bandgapmd_0.bg_pmosm_0.vbg.n16 3.097
R88916 bandgapmd_0.bg_pmosm_0.vbg.n25 bandgapmd_0.bg_pmosm_0.vbg.n24 2.337
R88917 bandgapmd_0.bg_pmosm_0.vbg.n45 bandgapmd_0.bg_pmosm_0.vbg.n44 2.331
R88918 bandgapmd_0.bg_pmosm_0.vbg.n65 bandgapmd_0.bg_pmosm_0.vbg.n64 2.251
R88919 bandgapmd_0.bg_pmosm_0.vbg.n60 bandgapmd_0.bg_pmosm_0.vbg.n59 2.25
R88920 bandgapmd_0.bg_pmosm_0.vbg.n58 bandgapmd_0.bg_pmosm_0.vbg.n57 2.25
R88921 bandgapmd_0.bg_pmosm_0.vbg.n56 bandgapmd_0.bg_pmosm_0.vbg.n42 2.25
R88922 bandgapmd_0.bg_pmosm_0.vbg.n55 bandgapmd_0.bg_pmosm_0.vbg.n54 2.25
R88923 bandgapmd_0.bg_pmosm_0.vbg.n46 bandgapmd_0.bg_pmosm_0.vbg.n45 2.25
R88924 bandgapmd_0.bg_pmosm_0.vbg.n48 bandgapmd_0.bg_pmosm_0.vbg.n47 2.25
R88925 bandgapmd_0.bg_pmosm_0.vbg.n50 bandgapmd_0.bg_pmosm_0.vbg.n49 2.25
R88926 bandgapmd_0.bg_pmosm_0.vbg.n51 bandgapmd_0.bg_pmosm_0.vbg.n43 2.25
R88927 bandgapmd_0.bg_pmosm_0.vbg.n53 bandgapmd_0.bg_pmosm_0.vbg.n52 2.25
R88928 bandgapmd_0.bg_pmosm_0.vbg.n66 bandgapmd_0.bg_pmosm_0.vbg.n40 2.25
R88929 bandgapmd_0.bg_pmosm_0.vbg.n68 bandgapmd_0.bg_pmosm_0.vbg.n67 2.25
R88930 bandgapmd_0.bg_pmosm_0.vbg.n61 bandgapmd_0.bg_pmosm_0.vbg.n41 2.25
R88931 bandgapmd_0.bg_pmosm_0.vbg.n63 bandgapmd_0.bg_pmosm_0.vbg.n62 2.25
R88932 bandgapmd_0.bg_pmosm_0.vbg.n70 bandgapmd_0.bg_pmosm_0.vbg.n69 1.776
R88933 bandgapmd_0.bg_resm_0.vbg bandgapmd_0.vbg 1.748
R88934 bandgapmd_0.bg_pmosm_0.vbg.n18 bandgapmd_0.bg_pmosm_0.vbg.n17 1.577
R88935 bandgapmd_0.bg_pmosm_0.vbg.n39 bandgapmd_0.bg_stupm_0.vbg 1.548
R88936 bandgapmd_0.bg_pmosm_0.vbg.n38 bandgapmd_0.bg_pmosm_0.vbg.n37 1.522
R88937 bandgapmd_0.bg_pmosm_0.vbg.n25 bandgapmd_0.bg_pmosm_0.vbg 1.217
R88938 bandgapmd_0.bg_pmosm_0.vbg.n54 bandgapmd_0.bg_pmosm_0.vbg.n53 1.178
R88939 bandgapmd_0.bg_pmosm_0.vbg.n64 bandgapmd_0.bg_pmosm_0.vbg.n63 1.137
R88940 bandgapmd_0.bg_pmosm_0.vbg.n49 bandgapmd_0.bg_pmosm_0.vbg.n48 1.135
R88941 bandgapmd_0.bg_pmosm_0.vbg.n39 bandgapmd_0.bg_pmosm_0.vbg.n32 1.135
R88942 bandgapmd_0.bg_pmosm_0.vbg.n59 bandgapmd_0.bg_pmosm_0.vbg.n58 1.13
R88943 bandgapmd_0.bg_pmosm_0.vbg.n12 bandgapmd_0.bg_pmosm_0.vbg.n11 1.066
R88944 bandgapmd_0.bg_stupm_0.vbg bandgapmd_0.bg_pmosm_0.vbg.n38 1.063
R88945 bandgapmd_0.bg_pmosm_0.vbg.n38 bandgapmd_0.bg_pmosm_0.vbg.n33 1.005
R88946 bandgapmd_0.bg_pmosm_0.vbg.n18 bandgapmd_0.bg_pmosm_0.vbg.n8 0.994
R88947 bandgapmd_0.bg_pmosm_0.vbg.n36 bandgapmd_0.bg_pmosm_0.vbg.n35 0.988
R88948 bandgapmd_0.bg_pmosm_0.vbg.n19 bandgapmd_0.bg_pmosm_0.vbg.n9 0.752
R88949 bandgapmd_0.bg_pmosm_0.vbg.n70 bandgapmd_0.bg_pmosm_0.vbg.n39 0.555
R88950 bandgapmd_0.bg_resm_0.vbg bandgapmd_0.bg_pmosm_0.vbg.t2 0.389
R88951 bandgapmd_0.bg_pmosm_0.vbg.n16 bandgapmd_0.bg_pmosm_0.vbg.n15 0.336
R88952 bandgapmd_0.bg_pmosm_0.vbg.n24 bandgapmd_0.bg_pmosm_0.vbg.n20 0.333
R88953 bandgapmd_0.bg_pmosm_0.vbg.n29 bandgapmd_0.bg_pmosm_0.vbg.n4 0.194
R88954 bandgapmd_0.bg_pmosm_0.vbg.n29 bandgapmd_0.bg_pmosm_0.vbg.n3 0.18
R88955 bandgapmd_0.bg_pmosm_0.vbg.n3 bandgapmd_0.bg_pmosm_0.vbg.n1 0.177
R88956 bandgapmd_0.bg_pmosm_0.vbg.n24 bandgapmd_0.bg_pmosm_0.vbg.n21 0.175
R88957 bandgapmd_0.bg_pmosm_0.vbg.n24 bandgapmd_0.bg_pmosm_0.vbg.n2 0.163
R88958 bandgapmd_0.bg_pmosm_0.vbg.n69 bandgapmd_0.bg_pmosm_0.vbg.t7 0.147
R88959 bandgapmd_0.bg_pmosm_0.vbg.n14 bandgapmd_0.bg_pmosm_0.vbg.n6 0.135
R88960 bandgapmd_0.bg_pmosm_0.vbg.n29 bandgapmd_0.bg_pmosm_0.vbg.n2 0.134
R88961 bandgapmd_0.bg_pmosm_0.vbg.n29 bandgapmd_0.bg_pmosm_0.vbg.n20 0.125
R88962 bandgapmd_0.bg_pmosm_0.vbg.n7 bandgapmd_0.bg_pmosm_0.vbg.n5 0.125
R88963 bandgapmd_0.bg_pmosm_0.vbg.n71 bandgapmd_0.bg_pmosm_0.vbg.n70 0.091
R88964 bandgapmd_0.bg_pmosm_0.vbg.n4 bandgapmd_0.bg_pmosm_0.vbg.n1 0.086
R88965 bandgapmd_0.bg_pmosm_0.vbg.n49 bandgapmd_0.bg_pmosm_0.vbg.n43 0.081
R88966 bandgapmd_0.bg_pmosm_0.vbg.n53 bandgapmd_0.bg_pmosm_0.vbg.n43 0.081
R88967 bandgapmd_0.bg_pmosm_0.vbg.n54 bandgapmd_0.bg_pmosm_0.vbg.n42 0.081
R88968 bandgapmd_0.bg_pmosm_0.vbg.n58 bandgapmd_0.bg_pmosm_0.vbg.n42 0.081
R88969 bandgapmd_0.bg_pmosm_0.vbg.n59 bandgapmd_0.bg_pmosm_0.vbg.n41 0.081
R88970 bandgapmd_0.bg_pmosm_0.vbg.n63 bandgapmd_0.bg_pmosm_0.vbg.n41 0.081
R88971 bandgapmd_0.bg_pmosm_0.vbg.n64 bandgapmd_0.bg_pmosm_0.vbg.n40 0.081
R88972 bandgapmd_0.bg_pmosm_0.vbg.n68 bandgapmd_0.bg_pmosm_0.vbg.n40 0.081
R88973 bandgapmd_0.bg_pmosm_0.vbg.n30 bandgapmd_0.bg_pmosm_0.vbg.n29 0.078
R88974 bandgapmd_0.bg_pmosm_0.vbg.n12 bandgapmd_0.bg_pmosm_0.vbg.n9 0.074
R88975 bandgapmd_0.bg_pmosm_0.vbg.n29 bandgapmd_0.bg_pmosm_0.vbg.n28 0.06
R88976 bandgapmd_0.bg_pmosm_0.vbg.n26 bandgapmd_0.bg_pmosm_0.vbg.n25 0.058
R88977 bandgapmd_0.bg_pmosm_0.vbg.n20 bandgapmd_0.bg_pmosm_0.vbg.n8 0.057
R88978 bandgapmd_0.bg_pmosm_0.vbg.n7 bandgapmd_0.bg_pmosm_0.vbg.n3 0.052
R88979 bandgapmd_0.bg_pmosm_0.vbg.n37 bandgapmd_0.bg_pmosm_0.vbg.n34 0.049
R88980 bandgapmd_0.bg_pmosm_0.vbg.n45 ldomc_0.vref 0.042
R88981 bandgapmd_0.bg_pmosm_0.vbg.n48 ldomc_0.vref 0.039
R88982 bandgapmd_0.bg_pmosm_0.vbg.n31 bandgapmd_0.bg_pmosm_0.vbg.n1 0.037
R88983 bandgapmd_0.vbg bandgapmd_0.bg_pmosm_0.vbg.n71 0.035
R88984 bandgapmd_0.bg_pmosm_0.vbg.n11 bandgapmd_0.bg_pmosm_0.vbg.n10 0.034
R88985 bandgapmd_0.bg_pmosm_0.vbg.n71 bandgapmd_0.vbg 0.033
R88986 bandgapmd_0.bg_pmosm_0.vbg.n28 bandgapmd_0.bg_pmosm_0.vbg.n21 0.032
R88987 bandgapmd_0.bg_pmosm_0.vbg.n15 bandgapmd_0.bg_pmosm_0.vbg.n2 0.028
R88988 bandgapmd_0.bg_pmosm_0.vbg.n14 bandgapmd_0.bg_pmosm_0.vbg.n4 0.025
R88989 bandgapmd_0.bg_pmosm_0.vbg.n66 bandgapmd_0.bg_pmosm_0.vbg.n65 0.024
R88990 bandgapmd_0.bg_pmosm_0.vbg.n67 bandgapmd_0.bg_pmosm_0.vbg.n66 0.024
R88991 bandgapmd_0.bg_pmosm_0.vbg.n51 bandgapmd_0.bg_pmosm_0.vbg.n50 0.024
R88992 bandgapmd_0.bg_pmosm_0.vbg.n52 bandgapmd_0.bg_pmosm_0.vbg.n51 0.024
R88993 bandgapmd_0.bg_pmosm_0.vbg.n56 bandgapmd_0.bg_pmosm_0.vbg.n55 0.024
R88994 bandgapmd_0.bg_pmosm_0.vbg.n57 bandgapmd_0.bg_pmosm_0.vbg.n56 0.024
R88995 bandgapmd_0.bg_pmosm_0.vbg.n61 bandgapmd_0.bg_pmosm_0.vbg.n60 0.024
R88996 bandgapmd_0.bg_pmosm_0.vbg.n62 bandgapmd_0.bg_pmosm_0.vbg.n61 0.024
R88997 bandgapmd_0.bg_pmosm_0.vbg.n23 bandgapmd_0.bg_pmosm_0.vbg.n22 0.023
R88998 bandgapmd_0.bg_pmosm_0.vbg.n22 bandgapmd_0.bg_pmosm_0.vbg.n0 0.022
R88999 bandgapmd_0.bg_pmosm_0.vbg.n44 ldomc_0.otaldom_0.pdiffm_0.inn 0.02
R89000 bandgapmd_0.bg_pmosm_0.vbg.n27 bandgapmd_0.bg_pmosm_0.vbg.n23 0.019
R89001 bandgapmd_0.bg_pmosm_0.vbg.n34 bandgapmd_0.bg_pmosm_0.vbg.n33 0.018
R89002 bandgapmd_0.bg_pmosm_0.vbg.n31 bandgapmd_0.bg_pmosm_0.vbg.n30 0.018
R89003 ldomc_0.otaldom_0.vref bandgapmd_0.bg_pmosm_0.vbg.n46 0.013
R89004 bandgapmd_0.bg_pmosm_0.vbg.n35 bandgapmd_0.bg_pmosm_0.vbg.n34 0.012
R89005 bandgapmd_0.bg_pmosm_0.vbg.n47 ldomc_0.otaldom_0.vref 0.011
R89006 bandgapmd_0.bg_pmosm_0.vbg.n8 bandgapmd_0.bg_pmosm_0.vbg.n7 0.01
R89007 bandgapmd_0.bg_pmosm_0.vbg.n29 bandgapmd_0.bg_pmosm_0.vbg.n6 0.01
R89008 bandgapmd_0.bg_pmosm_0.vbg.n29 bandgapmd_0.bg_pmosm_0.vbg.n5 0.01
R89009 bandgapmd_0.bg_pmosm_0.vbg.n27 bandgapmd_0.bg_pmosm_0.vbg.n26 0.007
R89010 bandgapmd_0.bg_pmosm_0.vbg.n13 bandgapmd_0.bg_pmosm_0.vbg.n12 0.006
R89011 bandgapmd_0.bg_pmosm_0.vbg.n15 bandgapmd_0.bg_pmosm_0.vbg.n14 0.005
R89012 bandgapmd_0.bg_pmosm_0.vbg.n46 ldomc_0.otaldom_0.pdiffm_0.inn 0.004
R89013 bandgapmd_0.bg_pmosm_0.vbg.n32 bandgapmd_0.bg_pmosm_0.vbg.n0 0.004
R89014 bandgapmd_0.otam_1.pcascodeupm_0.o1.n26 bandgapmd_0.otam_1.pcascodeupm_0.o1.n25 28.935
R89015 bandgapmd_0.otam_1.pcascodeupm_0.o1.n22 bandgapmd_0.otam_1.pcascodeupm_0.o1.n13 3.81
R89016 bandgapmd_0.otam_1.pcascodeupm_0.o1.n45 bandgapmd_0.otam_1.pcascodeupm_0.o1.t6 13.847
R89017 bandgapmd_0.otam_1.pcascodeupm_0.o1.n45 bandgapmd_0.otam_1.pcascodeupm_0.o1.t2 13.847
R89018 bandgapmd_0.otam_1.pcascodeupm_0.o1.n21 bandgapmd_0.otam_1.pcascodeupm_0.o1.t13 13.847
R89019 bandgapmd_0.otam_1.pcascodeupm_0.o1.n21 bandgapmd_0.otam_1.pcascodeupm_0.o1.t8 13.847
R89020 bandgapmd_0.otam_1.pcascodeupm_0.o1.n30 bandgapmd_0.otam_1.pcascodeupm_0.o1.t14 13.847
R89021 bandgapmd_0.otam_1.pcascodeupm_0.o1.n30 bandgapmd_0.otam_1.pcascodeupm_0.o1.t10 13.847
R89022 bandgapmd_0.otam_1.pcascodeupm_0.o1.n24 bandgapmd_0.otam_1.pcascodeupm_0.o1.t15 13.847
R89023 bandgapmd_0.otam_1.pcascodeupm_0.o1.n24 bandgapmd_0.otam_1.pcascodeupm_0.o1.t12 13.847
R89024 bandgapmd_0.otam_1.pcascodeupm_0.o1.n34 bandgapmd_0.otam_1.pcascodeupm_0.o1.t9 13.847
R89025 bandgapmd_0.otam_1.pcascodeupm_0.o1.n34 bandgapmd_0.otam_1.pcascodeupm_0.o1.t11 13.847
R89026 bandgapmd_0.otam_1.pcascodeupm_0.o1.n17 bandgapmd_0.otam_1.pcascodeupm_0.o1.t0 13.847
R89027 bandgapmd_0.otam_1.pcascodeupm_0.o1.n17 bandgapmd_0.otam_1.pcascodeupm_0.o1.t3 13.847
R89028 bandgapmd_0.otam_1.pcascodeupm_0.o1.n14 bandgapmd_0.otam_1.pcascodeupm_0.o1.t5 13.847
R89029 bandgapmd_0.otam_1.pcascodeupm_0.o1.n14 bandgapmd_0.otam_1.pcascodeupm_0.o1.t1 13.847
R89030 bandgapmd_0.otam_1.pcascodeupm_0.o1.n38 bandgapmd_0.otam_1.pcascodeupm_0.o1.t4 13.847
R89031 bandgapmd_0.otam_1.pcascodeupm_0.o1.n38 bandgapmd_0.otam_1.pcascodeupm_0.o1.t7 13.847
R89032 bandgapmd_0.otam_1.pcascodeupm_0.o1.n15 bandgapmd_0.otam_1.pcascodeupm_0.o1.n14 10.912
R89033 bandgapmd_0.otam_1.pcascodeupm_0.o1.n26 bandgapmd_0.otam_1.pcascodeupm_0.o1.n19 7.268
R89034 bandgapmd_0.otam_1.pcascodeupm_0.o1.n1 bandgapmd_0.otam_1.pcascodeupm_0.o1.n17 6.977
R89035 bandgapmd_0.otam_1.pcascodeupm_0.o1.n46 bandgapmd_0.otam_1.pcascodeupm_0.o1.n45 6.881
R89036 bandgapmd_0.otam_1.pcascodeupm_0.o1.n3 bandgapmd_0.otam_1.pcascodeupm_0.o1.n38 6.881
R89037 bandgapmd_0.otam_1.pcascodeupm_0.o1.n13 bandgapmd_0.otam_1.pcascodeupm_0.o1.n21 6.768
R89038 bandgapmd_0.otam_1.pcascodeupm_0.o1.n25 bandgapmd_0.otam_1.pcascodeupm_0.o1.n24 6.249
R89039 bandgapmd_0.otam_1.pcascodeupm_0.o1.n31 bandgapmd_0.otam_1.pcascodeupm_0.o1.n30 5.76
R89040 bandgapmd_0.otam_1.pcascodeupm_0.o1.n2 bandgapmd_0.otam_1.pcascodeupm_0.o1.n42 5.698
R89041 bandgapmd_0.otam_1.pcascodeupm_0.o1.n50 bandgapmd_0.otam_1.pcascodeupm_0.o1.n49 5.646
R89042 bandgapmd_0.otam_1.pcascodeupm_0.o1.n40 bandgapmd_0.otam_1.pcascodeupm_0.o1.n39 5.646
R89043 bandgapmd_0.otam_1.pcascodeupm_0.o1.n21 bandgapmd_0.otam_1.pcascodeupm_0.o1.n20 5.621
R89044 bandgapmd_0.otam_1.pcascodeupm_0.o1.n35 bandgapmd_0.otam_1.pcascodeupm_0.o1.n34 5.6
R89045 bandgapmd_0.otam_1.pcascodeupm_0.o1.n24 bandgapmd_0.otam_1.pcascodeupm_0.o1.n19 4.664
R89046 bandgapmd_0.otam_1.pcascodeupm_0.o1.n26 bandgapmd_0.otam_1.pcascodeupm_0.o1.n8 1.507
R89047 bandgapmd_0.otam_1.pcascodeupm_0.o1.n11 bandgapmd_0.otam_1.pcascodeupm_0.o1.n13 0.083
R89048 bandgapmd_0.otam_1.pcascodeupm_0.o1.n8 bandgapmd_0.otam_1.pcascodeupm_0.o1.n7 0.024
R89049 bandgapmd_0.otam_1.pcascodeupm_0.o1.n27 bandgapmd_0.otam_1.pcascodeupm_0.o1.n8 0.022
R89050 bandgapmd_0.otam_1.pcascodeupm_0.o1.n1 bandgapmd_0.otam_1.pcascodeupm_0.o1.n16 4.5
R89051 bandgapmd_0.otam_1.pcascodeupm_0.o1.n51 bandgapmd_0.otam_1.pcascodeupm_0.o1.n44 4.5
R89052 bandgapmd_0.otam_1.pcascodeupm_0.o1.n51 bandgapmd_0.otam_1.pcascodeupm_0.o1.n50 4.5
R89053 bandgapmd_0.otam_1.pcascodeupm_0.o1.n3 bandgapmd_0.otam_1.pcascodeupm_0.o1.n37 4.5
R89054 bandgapmd_0.otam_1.pcascodeupm_0.o1.n3 bandgapmd_0.otam_1.pcascodeupm_0.o1.n40 4.5
R89055 bandgapmd_0.otam_1.pcascodeupm_0.o1.n22 bandgapmd_0.otam_1.pcascodeupm_0.o1.n20 4.384
R89056 bandgapmd_0.otam_1.pcascodeupm_0.o1 bandgapmd_0.otam_1.pcascodeupm_0.o1.n53 3.614
R89057 bandgapmd_0.otam_1.pcascodeupm_0.o1.n5 bandgapmd_0.otam_1.pcascodeupm_0.o1.n29 3.03
R89058 bandgapmd_0.otam_1.pcascodeupm_0.o1.n1 bandgapmd_0.otam_1.pcascodeupm_0.o1.n18 2.693
R89059 bandgapmd_0.otam_1.pcascodeupm_0.o1.n9 bandgapmd_0.otam_1.pcascodeupm_0.o1.n27 0.77
R89060 bandgapmd_0.otam_1.pcascodeupm_0.o1.n2 bandgapmd_0.otam_1.pcascodeupm_0.o1.n43 2.252
R89061 bandgapmd_0.otam_1.pcascodeupm_0.o1.n15 bandgapmd_0.otam_1.pcascodeupm_0.o1.n1 2.252
R89062 bandgapmd_0.otam_1.pcascodeupm_0.o1.n2 bandgapmd_0.otam_1.pcascodeupm_0.o1.n51 2.25
R89063 bandgapmd_0.otam_1.pcascodeupm_0.o1.n2 bandgapmd_0.otam_1.pcascodeupm_0.o1.n52 2.25
R89064 bandgapmd_0.otam_1.pcascodeupm_0.o1.n19 bandgapmd_0.otam_1.pcascodeupm_0.o1.n6 2.182
R89065 bandgapmd_0.otam_1.pcascodeupm_0.o1.n3 bandgapmd_0.otam_1.pcascodeupm_0.o1.n10 2.087
R89066 bandgapmd_0.otam_1.pcascodeupm_0.o1.n23 bandgapmd_0.otam_1.pcascodeupm_0.o1.n12 2.664
R89067 bandgapmd_0.otam_1.pcascodeupm_0.o1.n53 bandgapmd_0.otam_1.pcascodeupm_0.o1.n35 1.377
R89068 bandgapmd_0.otam_1.pcascodeupm_0.o1 bandgapmd_0.otam_1.pcascodeupm_0.o1.n15 1.236
R89069 bandgapmd_0.otam_1.pcascodeupm_0.o1.n7 bandgapmd_0.otam_1.pcascodeupm_0.o1.n23 1.143
R89070 bandgapmd_0.otam_1.pmoslm_0.o1 bandgapmd_0.otam_1.pcascodeupm_0.o1.n9 1.137
R89071 bandgapmd_0.otam_1.pcascodeupm_0.o1.n20 bandgapmd_0.otam_1.pcascodeupm_0.o1.n11 1.033
R89072 bandgapmd_0.otam_1.pcascodeupm_0.o1.n5 bandgapmd_0.otam_1.pcascodeupm_0.o1.n31 0.999
R89073 bandgapmd_0.otam_1.pcascodeupm_0.o1.n32 bandgapmd_0.otam_1.pmoslm_0.o1 0.89
R89074 bandgapmd_0.otam_1.pcascodeupm_0.o1.n42 bandgapmd_0.otam_1.pcascodeupm_0.o1.n41 0.866
R89075 bandgapmd_0.otam_1.pcascodeupm_0.o1.n12 bandgapmd_0.otam_1.pcascodeupm_0.o1.n11 0.008
R89076 bandgapmd_0.otam_1.pcascodeupm_0.o1.n32 bandgapmd_0.otam_1.pcascodeupm_0.o1.n5 0.766
R89077 bandgapmd_0.otam_1.pcascodeupm_0.o1.n25 bandgapmd_0.otam_1.pcascodeupm_0.o1.n7 0.623
R89078 bandgapmd_0.otam_1.pcascodeupm_0.o1.n41 bandgapmd_0.otam_1.pcascodeupm_0.o1.n36 0.613
R89079 bandgapmd_0.otam_1.pcascodeupm_0.o1.n41 bandgapmd_0.otam_1.pcascodeupm_0.o1.n3 0.589
R89080 bandgapmd_0.otam_1.pcascodeupm_0.o1.n35 bandgapmd_0.otam_1.pcascodeupm_0.o1.n33 0.345
R89081 bandgapmd_0.otam_1.pcascodeupm_0.o1.n27 bandgapmd_0.otam_1.pcascodeupm_0.o1.n6 0.125
R89082 bandgapmd_0.otam_1.pcascodeupm_0.o1.n48 bandgapmd_0.otam_1.pcascodeupm_0.o1.n47 0.108
R89083 bandgapmd_0.otam_1.pcascodeupm_0.o1.n48 bandgapmd_0.otam_1.pcascodeupm_0.o1.n46 0.102
R89084 bandgapmd_0.otam_1.pcascodeupm_0.o1.n33 bandgapmd_0.otam_1.pcascodeupm_0.o1.n32 0.097
R89085 bandgapmd_0.otam_1.pcascodeupm_0.o1.n7 bandgapmd_0.otam_1.pcascodeupm_0.o1.n6 0.056
R89086 bandgapmd_0.otam_1.pcascodeupm_0.o1.n23 bandgapmd_0.otam_1.pcascodeupm_0.o1.n9 0.099
R89087 bandgapmd_0.otam_1.pcascodeupm_0.o1.n51 bandgapmd_0.otam_1.pcascodeupm_0.o1.n48 0.033
R89088 bandgapmd_0.otam_1.pcascodeupm_0.o1.n12 bandgapmd_0.otam_1.pcascodeupm_0.o1.n22 9.321
R89089 bandgapmd_0.otam_1.pcascodeupm_0.o1.n53 bandgapmd_0.otam_1.pcascodeupm_0.o1.n2 0.795
R89090 bandgapmd_0.otam_1.pcascodeupm_0.o1.n5 bandgapmd_0.otam_1.pcascodeupm_0.o1.n28 0.626
R89091 bandgapmd_0.otam_1.pcascodeupm_0.o1.n1 bandgapmd_0.otam_1.pcascodeupm_0.o1.n0 0.333
R89092 bandgapmd_0.otam_1.pcascodeupm_0.o1.n3 bandgapmd_0.otam_1.pcascodeupm_0.o1.n4 0.243
R89093 bandgapmd_0.bg_pmosm_0.comp.n2 bandgapmd_0.bg_pmosm_0.comp.t2 6.923
R89094 bandgapmd_0.bg_pmosm_0.comp.n2 bandgapmd_0.bg_pmosm_0.comp.t1 6.923
R89095 bandgapmd_0.bg_pmosm_0.comp.n7 bandgapmd_0.bg_pmosm_0.comp.n6 5.783
R89096 bandgapmd_0.bg_pmosm_0.comp.n30 bandgapmd_0.bg_pmosm_0.comp.n29 2.813
R89097 bandgapmd_0.bg_pmosm_0.comp.n23 bandgapmd_0.bg_pmosm_0.comp.n22 2.341
R89098 bandgapmd_0.bg_pmosm_0.comp.n20 bandgapmd_0.bg_pmosm_0.comp.n17 1.635
R89099 bandgapmd_0.bg_pmosm_0.comp.n15 bandgapmd_0.bg_pmosm_0.comp.n7 1.569
R89100 bandgapmd_0.bg_pmosm_0.comp.n5 bandgapmd_0.bg_pmosm_0.comp.n4 1.556
R89101 bandgapmd_0.bg_resm_0.comp bandgapmd_0.bg_pmosm_0.comp.n30 1.19
R89102 bandgapmd_0.bg_pmosm_0.comp.n23 bandgapmd_0.bg_pmosm_0.comp 0.626
R89103 bandgapmd_0.bg_pmosm_0.comp.n7 bandgapmd_0.bg_pmosm_0.comp.n2 0.554
R89104 bandgapmd_0.bg_pmosm_0.comp.n31 bandgapmd_0.bg_pmosm_0.comp.t0 0.388
R89105 bandgapmd_0.bg_pmosm_0.comp.n4 bandgapmd_0.bg_pmosm_0.comp.n3 0.376
R89106 bandgapmd_0.bg_pmosm_0.comp.n22 bandgapmd_0.bg_pmosm_0.comp.n21 0.32
R89107 bandgapmd_0.bg_pmosm_0.comp.n22 bandgapmd_0.bg_pmosm_0.comp.n1 0.182
R89108 bandgapmd_0.bg_pmosm_0.comp.n22 bandgapmd_0.bg_pmosm_0.comp.n16 0.163
R89109 bandgapmd_0.bg_pmosm_0.comp.n13 bandgapmd_0.bg_pmosm_0.comp.n12 0.086
R89110 bandgapmd_0.bg_pmosm_0.comp.n10 bandgapmd_0.bg_pmosm_0.comp.n8 0.081
R89111 bandgapmd_0.bg_pmosm_0.comp.n14 bandgapmd_0.bg_pmosm_0.comp.n10 0.072
R89112 bandgapmd_0.bg_pmosm_0.comp.n24 bandgapmd_0.bg_pmosm_0.comp.n23 0.062
R89113 bandgapmd_0.bg_pmosm_0.comp.n21 bandgapmd_0.bg_pmosm_0.comp.n20 0.055
R89114 bandgapmd_0.bg_pmosm_0.comp.n19 bandgapmd_0.bg_pmosm_0.comp.n18 0.05
R89115 bandgapmd_0.bg_pmosm_0.comp.n10 bandgapmd_0.bg_pmosm_0.comp.n9 0.041
R89116 bandgapmd_0.bg_pmosm_0.comp.n12 bandgapmd_0.bg_pmosm_0.comp.n11 0.038
R89117 bandgapmd_0.bg_pmosm_0.comp.n1 bandgapmd_0.bg_pmosm_0.comp.n0 0.033
R89118 bandgapmd_0.bg_pmosm_0.comp.n16 bandgapmd_0.bg_pmosm_0.comp.n15 0.028
R89119 bandgapmd_0.bg_pmosm_0.comp.n27 bandgapmd_0.bg_pmosm_0.comp.n26 0.025
R89120 bandgapmd_0.bg_pmosm_0.comp.n28 bandgapmd_0.bg_pmosm_0.comp.n27 0.024
R89121 bandgapmd_0.bg_pmosm_0.comp.n6 bandgapmd_0.bg_pmosm_0.comp.n5 0.023
R89122 bandgapmd_0.bg_pmosm_0.comp.n26 bandgapmd_0.bg_pmosm_0.comp.n25 0.02
R89123 bandgapmd_0.bg_pmosm_0.comp.n15 bandgapmd_0.bg_pmosm_0.comp.n14 0.015
R89124 bandgapmd_0.bg_pmosm_0.comp.n14 bandgapmd_0.bg_pmosm_0.comp.n13 0.014
R89125 bandgapmd_0.bg_pmosm_0.comp.n20 bandgapmd_0.bg_pmosm_0.comp.n19 0.01
R89126 bandgapmd_0.bg_pmosm_0.comp.n25 bandgapmd_0.bg_pmosm_0.comp.n24 0.007
R89127 bandgapmd_0.bg_resm_0.comp bandgapmd_0.bg_pmosm_0.comp.n31 0.006
R89128 bandgapmd_0.bg_pmosm_0.comp.n29 bandgapmd_0.bg_pmosm_0.comp.n28 0.004
R89129 biasbgr.n627 biasbgr.n624 28.481
R89130 biasbgr.n808 biasbgr.n805 28.481
R89131 biasbgr.n344 biasbgr.n341 28.481
R89132 biasbgr.n525 biasbgr.n522 28.481
R89133 biasbgr.n242 biasbgr.n239 28.481
R89134 biasbgr.n100 biasbgr.n99 28.481
R89135 biasbgr.n618 biasbgr.n617 13.176
R89136 biasbgr.n799 biasbgr.n798 13.176
R89137 biasbgr.n335 biasbgr.n334 13.176
R89138 biasbgr.n516 biasbgr.n515 13.176
R89139 biasbgr.n233 biasbgr.n232 13.176
R89140 biasbgr.n91 biasbgr.n90 13.176
R89141 biasbgr.n707 biasbgr.t2 12.05
R89142 biasbgr.n424 biasbgr.t5 12.05
R89143 biasbgr.n142 biasbgr.t4 12.05
R89144 biasbgr.n0 biasbgr.t0 12.05
R89145 biasbgr.n886 biasbgr.n879 9.3
R89146 biasbgr.n279 biasbgr.n278 9.3
R89147 biasbgr.n268 biasbgr.n267 9.3
R89148 biasbgr.n257 biasbgr.n256 9.3
R89149 biasbgr.n246 biasbgr.n245 9.3
R89150 biasbgr.n234 biasbgr.n233 9.3
R89151 biasbgr.n227 biasbgr.n226 9.3
R89152 biasbgr.n226 biasbgr.n225 9.3
R89153 biasbgr.n209 biasbgr.n208 9.3
R89154 biasbgr.n187 biasbgr.n186 9.3
R89155 biasbgr.n165 biasbgr.n164 9.3
R89156 biasbgr.n150 biasbgr.n149 9.3
R89157 biasbgr.n149 biasbgr.n148 9.3
R89158 biasbgr.n154 biasbgr.n153 9.3
R89159 biasbgr.n152 biasbgr.n151 9.3
R89160 biasbgr.n163 biasbgr.n162 9.3
R89161 biasbgr.n161 biasbgr.n160 9.3
R89162 biasbgr.n160 biasbgr.n159 9.3
R89163 biasbgr.n172 biasbgr.n171 9.3
R89164 biasbgr.n171 biasbgr.n170 9.3
R89165 biasbgr.n176 biasbgr.n175 9.3
R89166 biasbgr.n174 biasbgr.n173 9.3
R89167 biasbgr.n185 biasbgr.n184 9.3
R89168 biasbgr.n183 biasbgr.n182 9.3
R89169 biasbgr.n182 biasbgr.n181 9.3
R89170 biasbgr.n194 biasbgr.n193 9.3
R89171 biasbgr.n193 biasbgr.n192 9.3
R89172 biasbgr.n198 biasbgr.n197 9.3
R89173 biasbgr.n196 biasbgr.n195 9.3
R89174 biasbgr.n207 biasbgr.n206 9.3
R89175 biasbgr.n205 biasbgr.n204 9.3
R89176 biasbgr.n204 biasbgr.n203 9.3
R89177 biasbgr.n216 biasbgr.n215 9.3
R89178 biasbgr.n215 biasbgr.n214 9.3
R89179 biasbgr.n220 biasbgr.n219 9.3
R89180 biasbgr.n218 biasbgr.n217 9.3
R89181 biasbgr.n229 biasbgr.n228 9.3
R89182 biasbgr.n231 biasbgr.n230 9.3
R89183 biasbgr.n244 biasbgr.n243 9.3
R89184 biasbgr.n243 biasbgr.n242 9.3
R89185 biasbgr.n236 biasbgr.n235 9.3
R89186 biasbgr.n248 biasbgr.n247 9.3
R89187 biasbgr.n255 biasbgr.n254 9.3
R89188 biasbgr.n254 biasbgr.n253 9.3
R89189 biasbgr.n266 biasbgr.n265 9.3
R89190 biasbgr.n265 biasbgr.n264 9.3
R89191 biasbgr.n259 biasbgr.n258 9.3
R89192 biasbgr.n270 biasbgr.n269 9.3
R89193 biasbgr.n277 biasbgr.n276 9.3
R89194 biasbgr.n276 biasbgr.n275 9.3
R89195 biasbgr.n283 biasbgr.n282 9.3
R89196 biasbgr.n281 biasbgr.n280 9.3
R89197 biasbgr.n562 biasbgr.n561 9.3
R89198 biasbgr.n551 biasbgr.n550 9.3
R89199 biasbgr.n540 biasbgr.n539 9.3
R89200 biasbgr.n529 biasbgr.n528 9.3
R89201 biasbgr.n517 biasbgr.n516 9.3
R89202 biasbgr.n510 biasbgr.n509 9.3
R89203 biasbgr.n509 biasbgr.n508 9.3
R89204 biasbgr.n492 biasbgr.n491 9.3
R89205 biasbgr.n470 biasbgr.n469 9.3
R89206 biasbgr.n448 biasbgr.n447 9.3
R89207 biasbgr.n414 biasbgr.n413 9.3
R89208 biasbgr.n403 biasbgr.n402 9.3
R89209 biasbgr.n392 biasbgr.n391 9.3
R89210 biasbgr.n381 biasbgr.n380 9.3
R89211 biasbgr.n370 biasbgr.n369 9.3
R89212 biasbgr.n359 biasbgr.n358 9.3
R89213 biasbgr.n348 biasbgr.n347 9.3
R89214 biasbgr.n336 biasbgr.n335 9.3
R89215 biasbgr.n322 biasbgr.n321 9.3
R89216 biasbgr.n300 biasbgr.n299 9.3
R89217 biasbgr.n285 biasbgr.n284 9.3
R89218 biasbgr.n289 biasbgr.n288 9.3
R89219 biasbgr.n287 biasbgr.n286 9.3
R89220 biasbgr.n298 biasbgr.n297 9.3
R89221 biasbgr.n296 biasbgr.n295 9.3
R89222 biasbgr.n295 biasbgr.n294 9.3
R89223 biasbgr.n307 biasbgr.n306 9.3
R89224 biasbgr.n306 biasbgr.n305 9.3
R89225 biasbgr.n311 biasbgr.n310 9.3
R89226 biasbgr.n309 biasbgr.n308 9.3
R89227 biasbgr.n320 biasbgr.n319 9.3
R89228 biasbgr.n318 biasbgr.n317 9.3
R89229 biasbgr.n317 biasbgr.n316 9.3
R89230 biasbgr.n329 biasbgr.n328 9.3
R89231 biasbgr.n328 biasbgr.n327 9.3
R89232 biasbgr.n333 biasbgr.n332 9.3
R89233 biasbgr.n331 biasbgr.n330 9.3
R89234 biasbgr.n338 biasbgr.n337 9.3
R89235 biasbgr.n346 biasbgr.n345 9.3
R89236 biasbgr.n345 biasbgr.n344 9.3
R89237 biasbgr.n357 biasbgr.n356 9.3
R89238 biasbgr.n356 biasbgr.n355 9.3
R89239 biasbgr.n350 biasbgr.n349 9.3
R89240 biasbgr.n361 biasbgr.n360 9.3
R89241 biasbgr.n368 biasbgr.n367 9.3
R89242 biasbgr.n367 biasbgr.n366 9.3
R89243 biasbgr.n379 biasbgr.n378 9.3
R89244 biasbgr.n378 biasbgr.n377 9.3
R89245 biasbgr.n372 biasbgr.n371 9.3
R89246 biasbgr.n383 biasbgr.n382 9.3
R89247 biasbgr.n390 biasbgr.n389 9.3
R89248 biasbgr.n389 biasbgr.n388 9.3
R89249 biasbgr.n401 biasbgr.n400 9.3
R89250 biasbgr.n400 biasbgr.n399 9.3
R89251 biasbgr.n394 biasbgr.n393 9.3
R89252 biasbgr.n405 biasbgr.n404 9.3
R89253 biasbgr.n412 biasbgr.n411 9.3
R89254 biasbgr.n411 biasbgr.n410 9.3
R89255 biasbgr.n423 biasbgr.n422 9.3
R89256 biasbgr.n422 biasbgr.n421 9.3
R89257 biasbgr.n416 biasbgr.n415 9.3
R89258 biasbgr.n433 biasbgr.n432 9.3
R89259 biasbgr.n432 biasbgr.n431 9.3
R89260 biasbgr.n437 biasbgr.n436 9.3
R89261 biasbgr.n435 biasbgr.n434 9.3
R89262 biasbgr.n446 biasbgr.n445 9.3
R89263 biasbgr.n444 biasbgr.n443 9.3
R89264 biasbgr.n443 biasbgr.n442 9.3
R89265 biasbgr.n455 biasbgr.n454 9.3
R89266 biasbgr.n454 biasbgr.n453 9.3
R89267 biasbgr.n459 biasbgr.n458 9.3
R89268 biasbgr.n457 biasbgr.n456 9.3
R89269 biasbgr.n468 biasbgr.n467 9.3
R89270 biasbgr.n466 biasbgr.n465 9.3
R89271 biasbgr.n465 biasbgr.n464 9.3
R89272 biasbgr.n477 biasbgr.n476 9.3
R89273 biasbgr.n476 biasbgr.n475 9.3
R89274 biasbgr.n481 biasbgr.n480 9.3
R89275 biasbgr.n479 biasbgr.n478 9.3
R89276 biasbgr.n490 biasbgr.n489 9.3
R89277 biasbgr.n488 biasbgr.n487 9.3
R89278 biasbgr.n487 biasbgr.n486 9.3
R89279 biasbgr.n499 biasbgr.n498 9.3
R89280 biasbgr.n498 biasbgr.n497 9.3
R89281 biasbgr.n503 biasbgr.n502 9.3
R89282 biasbgr.n501 biasbgr.n500 9.3
R89283 biasbgr.n512 biasbgr.n511 9.3
R89284 biasbgr.n514 biasbgr.n513 9.3
R89285 biasbgr.n527 biasbgr.n526 9.3
R89286 biasbgr.n526 biasbgr.n525 9.3
R89287 biasbgr.n519 biasbgr.n518 9.3
R89288 biasbgr.n531 biasbgr.n530 9.3
R89289 biasbgr.n538 biasbgr.n537 9.3
R89290 biasbgr.n537 biasbgr.n536 9.3
R89291 biasbgr.n549 biasbgr.n548 9.3
R89292 biasbgr.n548 biasbgr.n547 9.3
R89293 biasbgr.n542 biasbgr.n541 9.3
R89294 biasbgr.n553 biasbgr.n552 9.3
R89295 biasbgr.n560 biasbgr.n559 9.3
R89296 biasbgr.n559 biasbgr.n558 9.3
R89297 biasbgr.n566 biasbgr.n565 9.3
R89298 biasbgr.n564 biasbgr.n563 9.3
R89299 biasbgr.n12 biasbgr.n11 9.3
R89300 biasbgr.n23 biasbgr.n22 9.3
R89301 biasbgr.n34 biasbgr.n33 9.3
R89302 biasbgr.n45 biasbgr.n44 9.3
R89303 biasbgr.n56 biasbgr.n55 9.3
R89304 biasbgr.n67 biasbgr.n66 9.3
R89305 biasbgr.n78 biasbgr.n77 9.3
R89306 biasbgr.n89 biasbgr.n88 9.3
R89307 biasbgr.n102 biasbgr.n101 9.3
R89308 biasbgr.n101 biasbgr.n100 9.3
R89309 biasbgr.n115 biasbgr.n114 9.3
R89310 biasbgr.n137 biasbgr.n136 9.3
R89311 biasbgr.n139 biasbgr.n138 9.3
R89312 biasbgr.n141 biasbgr.n140 9.3
R89313 biasbgr.n135 biasbgr.n134 9.3
R89314 biasbgr.n134 biasbgr.n133 9.3
R89315 biasbgr.n126 biasbgr.n125 9.3
R89316 biasbgr.n128 biasbgr.n127 9.3
R89317 biasbgr.n117 biasbgr.n116 9.3
R89318 biasbgr.n124 biasbgr.n123 9.3
R89319 biasbgr.n123 biasbgr.n122 9.3
R89320 biasbgr.n113 biasbgr.n112 9.3
R89321 biasbgr.n112 biasbgr.n111 9.3
R89322 biasbgr.n104 biasbgr.n103 9.3
R89323 biasbgr.n106 biasbgr.n105 9.3
R89324 biasbgr.n94 biasbgr.n93 9.3
R89325 biasbgr.n92 biasbgr.n91 9.3
R89326 biasbgr.n85 biasbgr.n84 9.3
R89327 biasbgr.n84 biasbgr.n83 9.3
R89328 biasbgr.n87 biasbgr.n86 9.3
R89329 biasbgr.n76 biasbgr.n75 9.3
R89330 biasbgr.n74 biasbgr.n73 9.3
R89331 biasbgr.n73 biasbgr.n72 9.3
R89332 biasbgr.n63 biasbgr.n62 9.3
R89333 biasbgr.n62 biasbgr.n61 9.3
R89334 biasbgr.n65 biasbgr.n64 9.3
R89335 biasbgr.n54 biasbgr.n53 9.3
R89336 biasbgr.n52 biasbgr.n51 9.3
R89337 biasbgr.n51 biasbgr.n50 9.3
R89338 biasbgr.n41 biasbgr.n40 9.3
R89339 biasbgr.n40 biasbgr.n39 9.3
R89340 biasbgr.n43 biasbgr.n42 9.3
R89341 biasbgr.n32 biasbgr.n31 9.3
R89342 biasbgr.n30 biasbgr.n29 9.3
R89343 biasbgr.n29 biasbgr.n28 9.3
R89344 biasbgr.n19 biasbgr.n18 9.3
R89345 biasbgr.n18 biasbgr.n17 9.3
R89346 biasbgr.n21 biasbgr.n20 9.3
R89347 biasbgr.n10 biasbgr.n9 9.3
R89348 biasbgr.n8 biasbgr.n7 9.3
R89349 biasbgr.n7 biasbgr.n6 9.3
R89350 biasbgr.n845 biasbgr.n844 9.3
R89351 biasbgr.n834 biasbgr.n833 9.3
R89352 biasbgr.n823 biasbgr.n822 9.3
R89353 biasbgr.n812 biasbgr.n811 9.3
R89354 biasbgr.n800 biasbgr.n799 9.3
R89355 biasbgr.n793 biasbgr.n792 9.3
R89356 biasbgr.n792 biasbgr.n791 9.3
R89357 biasbgr.n775 biasbgr.n774 9.3
R89358 biasbgr.n753 biasbgr.n752 9.3
R89359 biasbgr.n731 biasbgr.n730 9.3
R89360 biasbgr.n697 biasbgr.n696 9.3
R89361 biasbgr.n686 biasbgr.n685 9.3
R89362 biasbgr.n675 biasbgr.n674 9.3
R89363 biasbgr.n664 biasbgr.n663 9.3
R89364 biasbgr.n653 biasbgr.n652 9.3
R89365 biasbgr.n642 biasbgr.n641 9.3
R89366 biasbgr.n631 biasbgr.n630 9.3
R89367 biasbgr.n619 biasbgr.n618 9.3
R89368 biasbgr.n605 biasbgr.n604 9.3
R89369 biasbgr.n583 biasbgr.n582 9.3
R89370 biasbgr.n568 biasbgr.n567 9.3
R89371 biasbgr.n572 biasbgr.n571 9.3
R89372 biasbgr.n570 biasbgr.n569 9.3
R89373 biasbgr.n581 biasbgr.n580 9.3
R89374 biasbgr.n579 biasbgr.n578 9.3
R89375 biasbgr.n578 biasbgr.n577 9.3
R89376 biasbgr.n590 biasbgr.n589 9.3
R89377 biasbgr.n589 biasbgr.n588 9.3
R89378 biasbgr.n594 biasbgr.n593 9.3
R89379 biasbgr.n592 biasbgr.n591 9.3
R89380 biasbgr.n603 biasbgr.n602 9.3
R89381 biasbgr.n601 biasbgr.n600 9.3
R89382 biasbgr.n600 biasbgr.n599 9.3
R89383 biasbgr.n612 biasbgr.n611 9.3
R89384 biasbgr.n611 biasbgr.n610 9.3
R89385 biasbgr.n616 biasbgr.n615 9.3
R89386 biasbgr.n614 biasbgr.n613 9.3
R89387 biasbgr.n621 biasbgr.n620 9.3
R89388 biasbgr.n629 biasbgr.n628 9.3
R89389 biasbgr.n628 biasbgr.n627 9.3
R89390 biasbgr.n640 biasbgr.n639 9.3
R89391 biasbgr.n639 biasbgr.n638 9.3
R89392 biasbgr.n633 biasbgr.n632 9.3
R89393 biasbgr.n644 biasbgr.n643 9.3
R89394 biasbgr.n651 biasbgr.n650 9.3
R89395 biasbgr.n650 biasbgr.n649 9.3
R89396 biasbgr.n662 biasbgr.n661 9.3
R89397 biasbgr.n661 biasbgr.n660 9.3
R89398 biasbgr.n655 biasbgr.n654 9.3
R89399 biasbgr.n666 biasbgr.n665 9.3
R89400 biasbgr.n673 biasbgr.n672 9.3
R89401 biasbgr.n672 biasbgr.n671 9.3
R89402 biasbgr.n684 biasbgr.n683 9.3
R89403 biasbgr.n683 biasbgr.n682 9.3
R89404 biasbgr.n677 biasbgr.n676 9.3
R89405 biasbgr.n688 biasbgr.n687 9.3
R89406 biasbgr.n695 biasbgr.n694 9.3
R89407 biasbgr.n694 biasbgr.n693 9.3
R89408 biasbgr.n706 biasbgr.n705 9.3
R89409 biasbgr.n705 biasbgr.n704 9.3
R89410 biasbgr.n699 biasbgr.n698 9.3
R89411 biasbgr.n716 biasbgr.n715 9.3
R89412 biasbgr.n715 biasbgr.n714 9.3
R89413 biasbgr.n720 biasbgr.n719 9.3
R89414 biasbgr.n718 biasbgr.n717 9.3
R89415 biasbgr.n729 biasbgr.n728 9.3
R89416 biasbgr.n727 biasbgr.n726 9.3
R89417 biasbgr.n726 biasbgr.n725 9.3
R89418 biasbgr.n738 biasbgr.n737 9.3
R89419 biasbgr.n737 biasbgr.n736 9.3
R89420 biasbgr.n742 biasbgr.n741 9.3
R89421 biasbgr.n740 biasbgr.n739 9.3
R89422 biasbgr.n751 biasbgr.n750 9.3
R89423 biasbgr.n749 biasbgr.n748 9.3
R89424 biasbgr.n748 biasbgr.n747 9.3
R89425 biasbgr.n760 biasbgr.n759 9.3
R89426 biasbgr.n759 biasbgr.n758 9.3
R89427 biasbgr.n764 biasbgr.n763 9.3
R89428 biasbgr.n762 biasbgr.n761 9.3
R89429 biasbgr.n773 biasbgr.n772 9.3
R89430 biasbgr.n771 biasbgr.n770 9.3
R89431 biasbgr.n770 biasbgr.n769 9.3
R89432 biasbgr.n782 biasbgr.n781 9.3
R89433 biasbgr.n781 biasbgr.n780 9.3
R89434 biasbgr.n786 biasbgr.n785 9.3
R89435 biasbgr.n784 biasbgr.n783 9.3
R89436 biasbgr.n795 biasbgr.n794 9.3
R89437 biasbgr.n797 biasbgr.n796 9.3
R89438 biasbgr.n810 biasbgr.n809 9.3
R89439 biasbgr.n809 biasbgr.n808 9.3
R89440 biasbgr.n802 biasbgr.n801 9.3
R89441 biasbgr.n814 biasbgr.n813 9.3
R89442 biasbgr.n821 biasbgr.n820 9.3
R89443 biasbgr.n820 biasbgr.n819 9.3
R89444 biasbgr.n832 biasbgr.n831 9.3
R89445 biasbgr.n831 biasbgr.n830 9.3
R89446 biasbgr.n825 biasbgr.n824 9.3
R89447 biasbgr.n836 biasbgr.n835 9.3
R89448 biasbgr.n843 biasbgr.n842 9.3
R89449 biasbgr.n842 biasbgr.n841 9.3
R89450 biasbgr.n849 biasbgr.n848 9.3
R89451 biasbgr.n847 biasbgr.n846 9.3
R89452 biasbgr.n856 biasbgr.n855 9.3
R89453 biasbgr.n863 biasbgr.n862 9.3
R89454 biasbgr.n866 biasbgr.n865 9.3
R89455 biasbgr.n861 biasbgr.n860 9.3
R89456 biasbgr.n859 biasbgr.n858 9.3
R89457 biasbgr.n854 biasbgr.n853 9.3
R89458 biasbgr.n425 biasbgr.n424 8.764
R89459 biasbgr.n708 biasbgr.n707 8.764
R89460 biasbgr.n610 biasbgr.n609 8.763
R89461 biasbgr.n627 biasbgr.n626 8.763
R89462 biasbgr.n791 biasbgr.n790 8.763
R89463 biasbgr.n808 biasbgr.n807 8.763
R89464 biasbgr.n327 biasbgr.n326 8.763
R89465 biasbgr.n344 biasbgr.n343 8.763
R89466 biasbgr.n508 biasbgr.n507 8.763
R89467 biasbgr.n525 biasbgr.n524 8.763
R89468 biasbgr.n225 biasbgr.n224 8.763
R89469 biasbgr.n242 biasbgr.n241 8.763
R89470 biasbgr.n100 biasbgr.n98 8.763
R89471 biasbgr.n83 biasbgr.n82 8.763
R89472 biasbgr.n703 biasbgr.n702 8.215
R89473 biasbgr.n713 biasbgr.n712 8.215
R89474 biasbgr.n420 biasbgr.n419 8.215
R89475 biasbgr.n430 biasbgr.n429 8.215
R89476 biasbgr.n147 biasbgr.n146 8.215
R89477 biasbgr.n5 biasbgr.n4 8.215
R89478 biasbgr.n599 biasbgr.n598 7.668
R89479 biasbgr.n638 biasbgr.n637 7.668
R89480 biasbgr.n780 biasbgr.n779 7.668
R89481 biasbgr.n819 biasbgr.n818 7.668
R89482 biasbgr.n316 biasbgr.n315 7.668
R89483 biasbgr.n355 biasbgr.n354 7.668
R89484 biasbgr.n497 biasbgr.n496 7.668
R89485 biasbgr.n536 biasbgr.n535 7.668
R89486 biasbgr.n214 biasbgr.n213 7.668
R89487 biasbgr.n253 biasbgr.n252 7.668
R89488 biasbgr.n111 biasbgr.n110 7.668
R89489 biasbgr.n72 biasbgr.n71 7.668
R89490 biasbgr.n692 biasbgr.n691 7.12
R89491 biasbgr.n724 biasbgr.n723 7.12
R89492 biasbgr.n409 biasbgr.n408 7.12
R89493 biasbgr.n441 biasbgr.n440 7.12
R89494 biasbgr.n158 biasbgr.n157 7.12
R89495 biasbgr.n16 biasbgr.n15 7.12
R89496 biasbgr.n1 biasbgr.n0 6.915
R89497 biasbgr.n143 biasbgr.n142 6.914
R89498 biasbgr.n588 biasbgr.n587 6.572
R89499 biasbgr.n649 biasbgr.n648 6.572
R89500 biasbgr.n769 biasbgr.n768 6.572
R89501 biasbgr.n830 biasbgr.n829 6.572
R89502 biasbgr.n305 biasbgr.n304 6.572
R89503 biasbgr.n366 biasbgr.n365 6.572
R89504 biasbgr.n486 biasbgr.n485 6.572
R89505 biasbgr.n547 biasbgr.n546 6.572
R89506 biasbgr.n203 biasbgr.n202 6.572
R89507 biasbgr.n264 biasbgr.n263 6.572
R89508 biasbgr.n122 biasbgr.n121 6.572
R89509 biasbgr.n61 biasbgr.n60 6.572
R89510 biasbgr.n681 biasbgr.n680 6.025
R89511 biasbgr.n735 biasbgr.n734 6.025
R89512 biasbgr.n398 biasbgr.n397 6.025
R89513 biasbgr.n452 biasbgr.n451 6.025
R89514 biasbgr.n169 biasbgr.n168 6.025
R89515 biasbgr.n27 biasbgr.n26 6.025
R89516 biasbgr.n611 biasbgr.n607 6.023
R89517 biasbgr.n628 biasbgr.n623 6.023
R89518 biasbgr.n792 biasbgr.n788 6.023
R89519 biasbgr.n809 biasbgr.n804 6.023
R89520 biasbgr.n328 biasbgr.n324 6.023
R89521 biasbgr.n345 biasbgr.n340 6.023
R89522 biasbgr.n509 biasbgr.n505 6.023
R89523 biasbgr.n526 biasbgr.n521 6.023
R89524 biasbgr.n226 biasbgr.n222 6.023
R89525 biasbgr.n243 biasbgr.n238 6.023
R89526 biasbgr.n101 biasbgr.n96 6.023
R89527 biasbgr.n84 biasbgr.n80 6.023
R89528 biasbgr.n701 biasbgr.n700 5.647
R89529 biasbgr.n711 biasbgr.n710 5.647
R89530 biasbgr.n418 biasbgr.n417 5.647
R89531 biasbgr.n428 biasbgr.n427 5.647
R89532 biasbgr.n145 biasbgr.n144 5.647
R89533 biasbgr.n3 biasbgr.n2 5.647
R89534 biasbgr.n577 biasbgr.n576 5.477
R89535 biasbgr.n660 biasbgr.n659 5.477
R89536 biasbgr.n758 biasbgr.n757 5.477
R89537 biasbgr.n841 biasbgr.n840 5.477
R89538 biasbgr.n294 biasbgr.n293 5.477
R89539 biasbgr.n377 biasbgr.n376 5.477
R89540 biasbgr.n475 biasbgr.n474 5.477
R89541 biasbgr.n558 biasbgr.n557 5.477
R89542 biasbgr.n192 biasbgr.n191 5.477
R89543 biasbgr.n275 biasbgr.n274 5.477
R89544 biasbgr.n133 biasbgr.n132 5.477
R89545 biasbgr.n50 biasbgr.n49 5.477
R89546 biasbgr.n868 biasbgr.n867 5.343
R89547 biasbgr.n852 biasbgr.n851 5.28
R89548 biasbgr.n600 biasbgr.n596 5.27
R89549 biasbgr.n639 biasbgr.n635 5.27
R89550 biasbgr.n781 biasbgr.n777 5.27
R89551 biasbgr.n820 biasbgr.n816 5.27
R89552 biasbgr.n317 biasbgr.n313 5.27
R89553 biasbgr.n356 biasbgr.n352 5.27
R89554 biasbgr.n498 biasbgr.n494 5.27
R89555 biasbgr.n537 biasbgr.n533 5.27
R89556 biasbgr.n215 biasbgr.n211 5.27
R89557 biasbgr.n254 biasbgr.n250 5.27
R89558 biasbgr.n112 biasbgr.n108 5.27
R89559 biasbgr.n73 biasbgr.n69 5.27
R89560 biasbgr.n670 biasbgr.n669 4.929
R89561 biasbgr.n746 biasbgr.n745 4.929
R89562 biasbgr.n387 biasbgr.n386 4.929
R89563 biasbgr.n463 biasbgr.n462 4.929
R89564 biasbgr.n180 biasbgr.n179 4.929
R89565 biasbgr.n38 biasbgr.n37 4.929
R89566 biasbgr.n690 biasbgr.n689 4.894
R89567 biasbgr.n722 biasbgr.n721 4.894
R89568 biasbgr.n407 biasbgr.n406 4.894
R89569 biasbgr.n439 biasbgr.n438 4.894
R89570 biasbgr.n156 biasbgr.n155 4.894
R89571 biasbgr.n14 biasbgr.n13 4.894
R89572 biasbgr.n426 biasbgr.n425 4.65
R89573 biasbgr.n709 biasbgr.n708 4.65
R89574 biasbgr.n869 biasbgr.n868 4.65
R89575 biasbgr.n589 biasbgr.n585 4.517
R89576 biasbgr.n650 biasbgr.n646 4.517
R89577 biasbgr.n770 biasbgr.n766 4.517
R89578 biasbgr.n831 biasbgr.n827 4.517
R89579 biasbgr.n306 biasbgr.n302 4.517
R89580 biasbgr.n367 biasbgr.n363 4.517
R89581 biasbgr.n487 biasbgr.n483 4.517
R89582 biasbgr.n548 biasbgr.n544 4.517
R89583 biasbgr.n204 biasbgr.n200 4.517
R89584 biasbgr.n265 biasbgr.n261 4.517
R89585 biasbgr.n123 biasbgr.n119 4.517
R89586 biasbgr.n62 biasbgr.n58 4.517
R89587 biasbgr.n886 biasbgr.n872 4.47
R89588 biasbgr.n671 biasbgr.n670 4.381
R89589 biasbgr.n747 biasbgr.n746 4.381
R89590 biasbgr.n388 biasbgr.n387 4.381
R89591 biasbgr.n464 biasbgr.n463 4.381
R89592 biasbgr.n181 biasbgr.n180 4.381
R89593 biasbgr.n39 biasbgr.n38 4.381
R89594 biasbgr.n872 biasbgr.n871 4.214
R89595 biasbgr.n679 biasbgr.n678 4.141
R89596 biasbgr.n733 biasbgr.n732 4.141
R89597 biasbgr.n396 biasbgr.n395 4.141
R89598 biasbgr.n450 biasbgr.n449 4.141
R89599 biasbgr.n167 biasbgr.n166 4.141
R89600 biasbgr.n25 biasbgr.n24 4.141
R89601 biasbgr.n576 biasbgr.n575 3.834
R89602 biasbgr.n659 biasbgr.n658 3.834
R89603 biasbgr.n757 biasbgr.n756 3.834
R89604 biasbgr.n840 biasbgr.n839 3.834
R89605 biasbgr.n293 biasbgr.n292 3.834
R89606 biasbgr.n376 biasbgr.n375 3.834
R89607 biasbgr.n474 biasbgr.n473 3.834
R89608 biasbgr.n557 biasbgr.n556 3.834
R89609 biasbgr.n191 biasbgr.n190 3.834
R89610 biasbgr.n274 biasbgr.n273 3.834
R89611 biasbgr.n132 biasbgr.n131 3.834
R89612 biasbgr.n49 biasbgr.n48 3.834
R89613 biasbgr.n578 biasbgr.n574 3.764
R89614 biasbgr.n661 biasbgr.n657 3.764
R89615 biasbgr.n759 biasbgr.n755 3.764
R89616 biasbgr.n842 biasbgr.n838 3.764
R89617 biasbgr.n295 biasbgr.n291 3.764
R89618 biasbgr.n378 biasbgr.n374 3.764
R89619 biasbgr.n476 biasbgr.n472 3.764
R89620 biasbgr.n559 biasbgr.n555 3.764
R89621 biasbgr.n193 biasbgr.n189 3.764
R89622 biasbgr.n276 biasbgr.n272 3.764
R89623 biasbgr.n134 biasbgr.n130 3.764
R89624 biasbgr.n51 biasbgr.n47 3.764
R89625 biasbgr.n150 biasbgr.n143 3.409
R89626 biasbgr.n8 biasbgr.n1 3.408
R89627 biasbgr.n668 biasbgr.n667 3.388
R89628 biasbgr.n744 biasbgr.n743 3.388
R89629 biasbgr.n385 biasbgr.n384 3.388
R89630 biasbgr.n461 biasbgr.n460 3.388
R89631 biasbgr.n178 biasbgr.n177 3.388
R89632 biasbgr.n36 biasbgr.n35 3.388
R89633 biasbgr.n883 biasbgr.t3 3.306
R89634 biasbgr.n883 biasbgr.t1 3.306
R89635 biasbgr.n682 biasbgr.n681 3.286
R89636 biasbgr.n736 biasbgr.n735 3.286
R89637 biasbgr.n399 biasbgr.n398 3.286
R89638 biasbgr.n453 biasbgr.n452 3.286
R89639 biasbgr.n170 biasbgr.n169 3.286
R89640 biasbgr.n28 biasbgr.n27 3.286
R89641 biasbgr.n672 biasbgr.n668 3.011
R89642 biasbgr.n748 biasbgr.n744 3.011
R89643 biasbgr.n389 biasbgr.n385 3.011
R89644 biasbgr.n465 biasbgr.n461 3.011
R89645 biasbgr.n182 biasbgr.n178 3.011
R89646 biasbgr.n40 biasbgr.n36 3.011
R89647 biasbgr.n587 biasbgr.n586 2.738
R89648 biasbgr.n648 biasbgr.n647 2.738
R89649 biasbgr.n768 biasbgr.n767 2.738
R89650 biasbgr.n829 biasbgr.n828 2.738
R89651 biasbgr.n304 biasbgr.n303 2.738
R89652 biasbgr.n365 biasbgr.n364 2.738
R89653 biasbgr.n485 biasbgr.n484 2.738
R89654 biasbgr.n546 biasbgr.n545 2.738
R89655 biasbgr.n202 biasbgr.n201 2.738
R89656 biasbgr.n263 biasbgr.n262 2.738
R89657 biasbgr.n121 biasbgr.n120 2.738
R89658 biasbgr.n60 biasbgr.n59 2.738
R89659 biasbgr.n574 biasbgr.n573 2.635
R89660 biasbgr.n657 biasbgr.n656 2.635
R89661 biasbgr.n755 biasbgr.n754 2.635
R89662 biasbgr.n838 biasbgr.n837 2.635
R89663 biasbgr.n291 biasbgr.n290 2.635
R89664 biasbgr.n374 biasbgr.n373 2.635
R89665 biasbgr.n472 biasbgr.n471 2.635
R89666 biasbgr.n555 biasbgr.n554 2.635
R89667 biasbgr.n189 biasbgr.n188 2.635
R89668 biasbgr.n272 biasbgr.n271 2.635
R89669 biasbgr.n130 biasbgr.n129 2.635
R89670 biasbgr.n47 biasbgr.n46 2.635
R89671 biasbgr.n683 biasbgr.n679 2.258
R89672 biasbgr.n737 biasbgr.n733 2.258
R89673 biasbgr.n400 biasbgr.n396 2.258
R89674 biasbgr.n454 biasbgr.n450 2.258
R89675 biasbgr.n171 biasbgr.n167 2.258
R89676 biasbgr.n29 biasbgr.n25 2.258
R89677 biasbgr.n693 biasbgr.n692 2.19
R89678 biasbgr.n725 biasbgr.n724 2.19
R89679 biasbgr.n410 biasbgr.n409 2.19
R89680 biasbgr.n442 biasbgr.n441 2.19
R89681 biasbgr.n159 biasbgr.n158 2.19
R89682 biasbgr.n17 biasbgr.n16 2.19
R89683 biasbgr.n585 biasbgr.n584 1.882
R89684 biasbgr.n646 biasbgr.n645 1.882
R89685 biasbgr.n766 biasbgr.n765 1.882
R89686 biasbgr.n827 biasbgr.n826 1.882
R89687 biasbgr.n302 biasbgr.n301 1.882
R89688 biasbgr.n363 biasbgr.n362 1.882
R89689 biasbgr.n483 biasbgr.n482 1.882
R89690 biasbgr.n544 biasbgr.n543 1.882
R89691 biasbgr.n200 biasbgr.n199 1.882
R89692 biasbgr.n261 biasbgr.n260 1.882
R89693 biasbgr.n119 biasbgr.n118 1.882
R89694 biasbgr.n58 biasbgr.n57 1.882
R89695 biasbgr.n598 biasbgr.n597 1.643
R89696 biasbgr.n637 biasbgr.n636 1.643
R89697 biasbgr.n779 biasbgr.n778 1.643
R89698 biasbgr.n818 biasbgr.n817 1.643
R89699 biasbgr.n315 biasbgr.n314 1.643
R89700 biasbgr.n354 biasbgr.n353 1.643
R89701 biasbgr.n496 biasbgr.n495 1.643
R89702 biasbgr.n535 biasbgr.n534 1.643
R89703 biasbgr.n213 biasbgr.n212 1.643
R89704 biasbgr.n252 biasbgr.n251 1.643
R89705 biasbgr.n110 biasbgr.n109 1.643
R89706 biasbgr.n71 biasbgr.n70 1.643
R89707 biasbgr.n887 biasbgr.n886 1.517
R89708 biasbgr.n694 biasbgr.n690 1.505
R89709 biasbgr.n726 biasbgr.n722 1.505
R89710 biasbgr.n411 biasbgr.n407 1.505
R89711 biasbgr.n443 biasbgr.n439 1.505
R89712 biasbgr.n160 biasbgr.n156 1.505
R89713 biasbgr.n18 biasbgr.n14 1.505
R89714 biasbgr.n884 biasbgr.n883 1.467
R89715 biasbgr.n596 biasbgr.n595 1.129
R89716 biasbgr.n635 biasbgr.n634 1.129
R89717 biasbgr.n777 biasbgr.n776 1.129
R89718 biasbgr.n816 biasbgr.n815 1.129
R89719 biasbgr.n313 biasbgr.n312 1.129
R89720 biasbgr.n352 biasbgr.n351 1.129
R89721 biasbgr.n494 biasbgr.n493 1.129
R89722 biasbgr.n533 biasbgr.n532 1.129
R89723 biasbgr.n211 biasbgr.n210 1.129
R89724 biasbgr.n250 biasbgr.n249 1.129
R89725 biasbgr.n108 biasbgr.n107 1.129
R89726 biasbgr.n69 biasbgr.n68 1.129
R89727 biasbgr.n704 biasbgr.n703 1.095
R89728 biasbgr.n714 biasbgr.n713 1.095
R89729 biasbgr.n421 biasbgr.n420 1.095
R89730 biasbgr.n431 biasbgr.n430 1.095
R89731 biasbgr.n148 biasbgr.n147 1.095
R89732 biasbgr.n6 biasbgr.n5 1.095
R89733 biasbgr.n705 biasbgr.n701 0.752
R89734 biasbgr.n715 biasbgr.n711 0.752
R89735 biasbgr.n422 biasbgr.n418 0.752
R89736 biasbgr.n432 biasbgr.n428 0.752
R89737 biasbgr.n149 biasbgr.n145 0.752
R89738 biasbgr.n7 biasbgr.n3 0.752
R89739 biasbgr.n885 biasbgr.n884 0.562
R89740 biasbgr.n609 biasbgr.n608 0.547
R89741 biasbgr.n626 biasbgr.n625 0.547
R89742 biasbgr.n790 biasbgr.n789 0.547
R89743 biasbgr.n807 biasbgr.n806 0.547
R89744 biasbgr.n326 biasbgr.n325 0.547
R89745 biasbgr.n343 biasbgr.n342 0.547
R89746 biasbgr.n507 biasbgr.n506 0.547
R89747 biasbgr.n524 biasbgr.n523 0.547
R89748 biasbgr.n224 biasbgr.n223 0.547
R89749 biasbgr.n241 biasbgr.n240 0.547
R89750 biasbgr.n98 biasbgr.n97 0.547
R89751 biasbgr.n82 biasbgr.n81 0.547
R89752 bandgapmd_0.otam_1.bias biasbgr.n889 0.537
R89753 biasbgr.n858 biasbgr.n857 0.461
R89754 biasbgr.n865 biasbgr.n864 0.43
R89755 biasbgr.n607 biasbgr.n606 0.376
R89756 biasbgr.n623 biasbgr.n622 0.376
R89757 biasbgr.n788 biasbgr.n787 0.376
R89758 biasbgr.n804 biasbgr.n803 0.376
R89759 biasbgr.n324 biasbgr.n323 0.376
R89760 biasbgr.n340 biasbgr.n339 0.376
R89761 biasbgr.n505 biasbgr.n504 0.376
R89762 biasbgr.n521 biasbgr.n520 0.376
R89763 biasbgr.n222 biasbgr.n221 0.376
R89764 biasbgr.n238 biasbgr.n237 0.376
R89765 biasbgr.n96 biasbgr.n95 0.376
R89766 biasbgr.n80 biasbgr.n79 0.376
R89767 biasbgr.n285 biasbgr.n283 0.323
R89768 biasbgr.n568 biasbgr.n566 0.323
R89769 biasbgr bandgapmd_0.bias 0.268
R89770 bandgapmd_0.otam_1.bias biasbgr 0.202
R89771 biasbgr.n852 biasbgr.n850 0.144
R89772 biasbgr.n234 biasbgr.n231 0.128
R89773 biasbgr.n336 biasbgr.n333 0.128
R89774 biasbgr.n426 biasbgr.n423 0.128
R89775 biasbgr.n433 biasbgr.n426 0.128
R89776 biasbgr.n517 biasbgr.n514 0.128
R89777 biasbgr.n92 biasbgr.n89 0.128
R89778 biasbgr.n619 biasbgr.n616 0.128
R89779 biasbgr.n709 biasbgr.n706 0.128
R89780 biasbgr.n716 biasbgr.n709 0.128
R89781 biasbgr.n800 biasbgr.n797 0.128
R89782 biasbgr.n161 biasbgr.n154 0.097
R89783 biasbgr.n172 biasbgr.n165 0.097
R89784 biasbgr.n183 biasbgr.n176 0.097
R89785 biasbgr.n194 biasbgr.n187 0.097
R89786 biasbgr.n205 biasbgr.n198 0.097
R89787 biasbgr.n216 biasbgr.n209 0.097
R89788 biasbgr.n227 biasbgr.n220 0.097
R89789 biasbgr.n246 biasbgr.n244 0.097
R89790 biasbgr.n257 biasbgr.n255 0.097
R89791 biasbgr.n268 biasbgr.n266 0.097
R89792 biasbgr.n279 biasbgr.n277 0.097
R89793 biasbgr.n296 biasbgr.n289 0.097
R89794 biasbgr.n307 biasbgr.n300 0.097
R89795 biasbgr.n318 biasbgr.n311 0.097
R89796 biasbgr.n329 biasbgr.n322 0.097
R89797 biasbgr.n348 biasbgr.n346 0.097
R89798 biasbgr.n359 biasbgr.n357 0.097
R89799 biasbgr.n370 biasbgr.n368 0.097
R89800 biasbgr.n381 biasbgr.n379 0.097
R89801 biasbgr.n392 biasbgr.n390 0.097
R89802 biasbgr.n403 biasbgr.n401 0.097
R89803 biasbgr.n414 biasbgr.n412 0.097
R89804 biasbgr.n444 biasbgr.n437 0.097
R89805 biasbgr.n455 biasbgr.n448 0.097
R89806 biasbgr.n466 biasbgr.n459 0.097
R89807 biasbgr.n477 biasbgr.n470 0.097
R89808 biasbgr.n488 biasbgr.n481 0.097
R89809 biasbgr.n499 biasbgr.n492 0.097
R89810 biasbgr.n510 biasbgr.n503 0.097
R89811 biasbgr.n529 biasbgr.n527 0.097
R89812 biasbgr.n540 biasbgr.n538 0.097
R89813 biasbgr.n551 biasbgr.n549 0.097
R89814 biasbgr.n562 biasbgr.n560 0.097
R89815 biasbgr.n137 biasbgr.n135 0.097
R89816 biasbgr.n126 biasbgr.n124 0.097
R89817 biasbgr.n115 biasbgr.n113 0.097
R89818 biasbgr.n104 biasbgr.n102 0.097
R89819 biasbgr.n85 biasbgr.n78 0.097
R89820 biasbgr.n74 biasbgr.n67 0.097
R89821 biasbgr.n63 biasbgr.n56 0.097
R89822 biasbgr.n52 biasbgr.n45 0.097
R89823 biasbgr.n41 biasbgr.n34 0.097
R89824 biasbgr.n30 biasbgr.n23 0.097
R89825 biasbgr.n19 biasbgr.n12 0.097
R89826 biasbgr.n579 biasbgr.n572 0.097
R89827 biasbgr.n590 biasbgr.n583 0.097
R89828 biasbgr.n601 biasbgr.n594 0.097
R89829 biasbgr.n612 biasbgr.n605 0.097
R89830 biasbgr.n631 biasbgr.n629 0.097
R89831 biasbgr.n642 biasbgr.n640 0.097
R89832 biasbgr.n653 biasbgr.n651 0.097
R89833 biasbgr.n664 biasbgr.n662 0.097
R89834 biasbgr.n675 biasbgr.n673 0.097
R89835 biasbgr.n686 biasbgr.n684 0.097
R89836 biasbgr.n697 biasbgr.n695 0.097
R89837 biasbgr.n727 biasbgr.n720 0.097
R89838 biasbgr.n738 biasbgr.n731 0.097
R89839 biasbgr.n749 biasbgr.n742 0.097
R89840 biasbgr.n760 biasbgr.n753 0.097
R89841 biasbgr.n771 biasbgr.n764 0.097
R89842 biasbgr.n782 biasbgr.n775 0.097
R89843 biasbgr.n793 biasbgr.n786 0.097
R89844 biasbgr.n812 biasbgr.n810 0.097
R89845 biasbgr.n823 biasbgr.n821 0.097
R89846 biasbgr.n834 biasbgr.n832 0.097
R89847 biasbgr.n845 biasbgr.n843 0.097
R89848 biasbgr.n886 biasbgr.n876 0.088
R89849 biasbgr.n854 biasbgr.n852 0.084
R89850 biasbgr.n850 biasbgr.n141 0.077
R89851 biasbgr.n886 biasbgr.n881 0.075
R89852 biasbgr.n861 biasbgr.n859 0.073
R89853 biasbgr.n869 biasbgr.n866 0.073
R89854 biasbgr.n878 biasbgr.n877 0.071
R89855 biasbgr.n850 biasbgr.n849 0.069
R89856 biasbgr.n874 biasbgr.n873 0.065
R89857 biasbgr.n887 biasbgr 0.061
R89858 biasbgr.n886 biasbgr.n870 0.033
R89859 biasbgr.n886 biasbgr.n885 0.033
R89860 biasbgr.n229 biasbgr.n227 0.029
R89861 biasbgr.n244 biasbgr.n236 0.029
R89862 biasbgr.n331 biasbgr.n329 0.029
R89863 biasbgr.n346 biasbgr.n338 0.029
R89864 biasbgr.n512 biasbgr.n510 0.029
R89865 biasbgr.n527 biasbgr.n519 0.029
R89866 biasbgr.n102 biasbgr.n94 0.029
R89867 biasbgr.n87 biasbgr.n85 0.029
R89868 biasbgr.n614 biasbgr.n612 0.029
R89869 biasbgr.n629 biasbgr.n621 0.029
R89870 biasbgr.n795 biasbgr.n793 0.029
R89871 biasbgr.n810 biasbgr.n802 0.029
R89872 biasbgr.n154 biasbgr.n152 0.027
R89873 biasbgr.n416 biasbgr.n414 0.027
R89874 biasbgr.n437 biasbgr.n435 0.027
R89875 biasbgr.n12 biasbgr.n10 0.027
R89876 biasbgr.n699 biasbgr.n697 0.027
R89877 biasbgr.n720 biasbgr.n718 0.027
R89878 biasbgr.n218 biasbgr.n216 0.025
R89879 biasbgr.n255 biasbgr.n248 0.025
R89880 biasbgr.n320 biasbgr.n318 0.025
R89881 biasbgr.n357 biasbgr.n350 0.025
R89882 biasbgr.n501 biasbgr.n499 0.025
R89883 biasbgr.n538 biasbgr.n531 0.025
R89884 biasbgr.n113 biasbgr.n106 0.025
R89885 biasbgr.n76 biasbgr.n74 0.025
R89886 biasbgr.n603 biasbgr.n601 0.025
R89887 biasbgr.n640 biasbgr.n633 0.025
R89888 biasbgr.n784 biasbgr.n782 0.025
R89889 biasbgr.n821 biasbgr.n814 0.025
R89890 biasbgr.n165 biasbgr.n163 0.023
R89891 biasbgr.n405 biasbgr.n403 0.023
R89892 biasbgr.n448 biasbgr.n446 0.023
R89893 biasbgr.n23 biasbgr.n21 0.023
R89894 biasbgr.n688 biasbgr.n686 0.023
R89895 biasbgr.n731 biasbgr.n729 0.023
R89896 biasbgr.n207 biasbgr.n205 0.022
R89897 biasbgr.n266 biasbgr.n259 0.022
R89898 biasbgr.n309 biasbgr.n307 0.022
R89899 biasbgr.n368 biasbgr.n361 0.022
R89900 biasbgr.n490 biasbgr.n488 0.022
R89901 biasbgr.n549 biasbgr.n542 0.022
R89902 biasbgr.n124 biasbgr.n117 0.022
R89903 biasbgr.n65 biasbgr.n63 0.022
R89904 biasbgr.n592 biasbgr.n590 0.022
R89905 biasbgr.n651 biasbgr.n644 0.022
R89906 biasbgr.n773 biasbgr.n771 0.022
R89907 biasbgr.n832 biasbgr.n825 0.022
R89908 biasbgr.n176 biasbgr.n174 0.02
R89909 biasbgr.n394 biasbgr.n392 0.02
R89910 biasbgr.n459 biasbgr.n457 0.02
R89911 biasbgr.n34 biasbgr.n32 0.02
R89912 biasbgr.n677 biasbgr.n675 0.02
R89913 biasbgr.n742 biasbgr.n740 0.02
R89914 biasbgr.n196 biasbgr.n194 0.018
R89915 biasbgr.n277 biasbgr.n270 0.018
R89916 biasbgr.n298 biasbgr.n296 0.018
R89917 biasbgr.n379 biasbgr.n372 0.018
R89918 biasbgr.n479 biasbgr.n477 0.018
R89919 biasbgr.n560 biasbgr.n553 0.018
R89920 biasbgr.n135 biasbgr.n128 0.018
R89921 biasbgr.n54 biasbgr.n52 0.018
R89922 biasbgr.n581 biasbgr.n579 0.018
R89923 biasbgr.n662 biasbgr.n655 0.018
R89924 biasbgr.n762 biasbgr.n760 0.018
R89925 biasbgr.n843 biasbgr.n836 0.018
R89926 biasbgr.n187 biasbgr.n185 0.016
R89927 biasbgr.n281 biasbgr.n279 0.016
R89928 biasbgr.n289 biasbgr.n287 0.016
R89929 biasbgr.n383 biasbgr.n381 0.016
R89930 biasbgr.n470 biasbgr.n468 0.016
R89931 biasbgr.n564 biasbgr.n562 0.016
R89932 biasbgr.n139 biasbgr.n137 0.016
R89933 biasbgr.n45 biasbgr.n43 0.016
R89934 biasbgr.n572 biasbgr.n570 0.016
R89935 biasbgr.n666 biasbgr.n664 0.016
R89936 biasbgr.n753 biasbgr.n751 0.016
R89937 biasbgr.n847 biasbgr.n845 0.016
R89938 biasbgr.n859 biasbgr.n856 0.015
R89939 biasbgr.n886 biasbgr.n878 0.014
R89940 biasbgr.n881 biasbgr.n880 0.014
R89941 biasbgr.n185 biasbgr.n183 0.014
R89942 biasbgr.n283 biasbgr.n281 0.014
R89943 biasbgr.n287 biasbgr.n285 0.014
R89944 biasbgr.n390 biasbgr.n383 0.014
R89945 biasbgr.n468 biasbgr.n466 0.014
R89946 biasbgr.n566 biasbgr.n564 0.014
R89947 biasbgr.n141 biasbgr.n139 0.014
R89948 biasbgr.n43 biasbgr.n41 0.014
R89949 biasbgr.n570 biasbgr.n568 0.014
R89950 biasbgr.n673 biasbgr.n666 0.014
R89951 biasbgr.n751 biasbgr.n749 0.014
R89952 biasbgr.n849 biasbgr.n847 0.014
R89953 biasbgr.n888 biasbgr.n887 0.014
R89954 biasbgr.n886 biasbgr.n874 0.013
R89955 biasbgr.n198 biasbgr.n196 0.012
R89956 biasbgr.n270 biasbgr.n268 0.012
R89957 biasbgr.n300 biasbgr.n298 0.012
R89958 biasbgr.n372 biasbgr.n370 0.012
R89959 biasbgr.n481 biasbgr.n479 0.012
R89960 biasbgr.n553 biasbgr.n551 0.012
R89961 biasbgr.n128 biasbgr.n126 0.012
R89962 biasbgr.n56 biasbgr.n54 0.012
R89963 biasbgr.n583 biasbgr.n581 0.012
R89964 biasbgr.n655 biasbgr.n653 0.012
R89965 biasbgr.n764 biasbgr.n762 0.012
R89966 biasbgr.n836 biasbgr.n834 0.012
R89967 biasbgr.n866 biasbgr.n863 0.012
R89968 biasbgr.n174 biasbgr.n172 0.011
R89969 biasbgr.n401 biasbgr.n394 0.011
R89970 biasbgr.n457 biasbgr.n455 0.011
R89971 biasbgr.n32 biasbgr.n30 0.011
R89972 biasbgr.n684 biasbgr.n677 0.011
R89973 biasbgr.n740 biasbgr.n738 0.011
R89974 biasbgr.n863 biasbgr.n861 0.011
R89975 biasbgr.n889 biasbgr.n888 0.011
R89976 biasbgr.n209 biasbgr.n207 0.009
R89977 biasbgr.n259 biasbgr.n257 0.009
R89978 biasbgr.n311 biasbgr.n309 0.009
R89979 biasbgr.n361 biasbgr.n359 0.009
R89980 biasbgr.n492 biasbgr.n490 0.009
R89981 biasbgr.n542 biasbgr.n540 0.009
R89982 biasbgr.n117 biasbgr.n115 0.009
R89983 biasbgr.n67 biasbgr.n65 0.009
R89984 biasbgr.n594 biasbgr.n592 0.009
R89985 biasbgr.n644 biasbgr.n642 0.009
R89986 biasbgr.n775 biasbgr.n773 0.009
R89987 biasbgr.n825 biasbgr.n823 0.009
R89988 biasbgr.n886 biasbgr.n869 0.009
R89989 biasbgr.n876 biasbgr.n875 0.009
R89990 biasbgr.n885 biasbgr.n882 0.008
R89991 biasbgr.n856 biasbgr.n854 0.008
R89992 biasbgr.n163 biasbgr.n161 0.007
R89993 biasbgr.n412 biasbgr.n405 0.007
R89994 biasbgr.n446 biasbgr.n444 0.007
R89995 biasbgr.n21 biasbgr.n19 0.007
R89996 biasbgr.n695 biasbgr.n688 0.007
R89997 biasbgr.n729 biasbgr.n727 0.007
R89998 biasbgr.n220 biasbgr.n218 0.005
R89999 biasbgr.n248 biasbgr.n246 0.005
R90000 biasbgr.n322 biasbgr.n320 0.005
R90001 biasbgr.n350 biasbgr.n348 0.005
R90002 biasbgr.n503 biasbgr.n501 0.005
R90003 biasbgr.n531 biasbgr.n529 0.005
R90004 biasbgr.n106 biasbgr.n104 0.005
R90005 biasbgr.n78 biasbgr.n76 0.005
R90006 biasbgr.n605 biasbgr.n603 0.005
R90007 biasbgr.n633 biasbgr.n631 0.005
R90008 biasbgr.n786 biasbgr.n784 0.005
R90009 biasbgr.n814 biasbgr.n812 0.005
R90010 biasbgr.n152 biasbgr.n150 0.003
R90011 biasbgr.n423 biasbgr.n416 0.003
R90012 biasbgr.n435 biasbgr.n433 0.003
R90013 biasbgr.n10 biasbgr.n8 0.003
R90014 biasbgr.n706 biasbgr.n699 0.003
R90015 biasbgr.n718 biasbgr.n716 0.003
R90016 biasbgr.n231 biasbgr.n229 0.001
R90017 biasbgr.n236 biasbgr.n234 0.001
R90018 biasbgr.n333 biasbgr.n331 0.001
R90019 biasbgr.n338 biasbgr.n336 0.001
R90020 biasbgr.n514 biasbgr.n512 0.001
R90021 biasbgr.n519 biasbgr.n517 0.001
R90022 biasbgr.n94 biasbgr.n92 0.001
R90023 biasbgr.n89 biasbgr.n87 0.001
R90024 biasbgr.n616 biasbgr.n614 0.001
R90025 biasbgr.n621 biasbgr.n619 0.001
R90026 biasbgr.n797 biasbgr.n795 0.001
R90027 biasbgr.n802 biasbgr.n800 0.001
R90028 biasldo.n627 biasldo.n624 28.481
R90029 biasldo.n808 biasldo.n805 28.481
R90030 biasldo.n344 biasldo.n341 28.481
R90031 biasldo.n525 biasldo.n522 28.481
R90032 biasldo.n242 biasldo.n239 28.481
R90033 biasldo.n100 biasldo.n99 28.481
R90034 biasldo.n618 biasldo.n617 13.176
R90035 biasldo.n799 biasldo.n798 13.176
R90036 biasldo.n335 biasldo.n334 13.176
R90037 biasldo.n516 biasldo.n515 13.176
R90038 biasldo.n233 biasldo.n232 13.176
R90039 biasldo.n91 biasldo.n90 13.176
R90040 biasldo.n707 biasldo.t2 12.05
R90041 biasldo.n424 biasldo.t4 12.05
R90042 biasldo.n142 biasldo.t5 12.05
R90043 biasldo.n0 biasldo.t0 12.05
R90044 biasldo.n886 biasldo.n879 9.3
R90045 biasldo.n279 biasldo.n278 9.3
R90046 biasldo.n268 biasldo.n267 9.3
R90047 biasldo.n257 biasldo.n256 9.3
R90048 biasldo.n246 biasldo.n245 9.3
R90049 biasldo.n234 biasldo.n233 9.3
R90050 biasldo.n227 biasldo.n226 9.3
R90051 biasldo.n226 biasldo.n225 9.3
R90052 biasldo.n209 biasldo.n208 9.3
R90053 biasldo.n187 biasldo.n186 9.3
R90054 biasldo.n165 biasldo.n164 9.3
R90055 biasldo.n150 biasldo.n149 9.3
R90056 biasldo.n149 biasldo.n148 9.3
R90057 biasldo.n154 biasldo.n153 9.3
R90058 biasldo.n152 biasldo.n151 9.3
R90059 biasldo.n163 biasldo.n162 9.3
R90060 biasldo.n161 biasldo.n160 9.3
R90061 biasldo.n160 biasldo.n159 9.3
R90062 biasldo.n172 biasldo.n171 9.3
R90063 biasldo.n171 biasldo.n170 9.3
R90064 biasldo.n176 biasldo.n175 9.3
R90065 biasldo.n174 biasldo.n173 9.3
R90066 biasldo.n185 biasldo.n184 9.3
R90067 biasldo.n183 biasldo.n182 9.3
R90068 biasldo.n182 biasldo.n181 9.3
R90069 biasldo.n194 biasldo.n193 9.3
R90070 biasldo.n193 biasldo.n192 9.3
R90071 biasldo.n198 biasldo.n197 9.3
R90072 biasldo.n196 biasldo.n195 9.3
R90073 biasldo.n207 biasldo.n206 9.3
R90074 biasldo.n205 biasldo.n204 9.3
R90075 biasldo.n204 biasldo.n203 9.3
R90076 biasldo.n216 biasldo.n215 9.3
R90077 biasldo.n215 biasldo.n214 9.3
R90078 biasldo.n220 biasldo.n219 9.3
R90079 biasldo.n218 biasldo.n217 9.3
R90080 biasldo.n229 biasldo.n228 9.3
R90081 biasldo.n231 biasldo.n230 9.3
R90082 biasldo.n244 biasldo.n243 9.3
R90083 biasldo.n243 biasldo.n242 9.3
R90084 biasldo.n236 biasldo.n235 9.3
R90085 biasldo.n248 biasldo.n247 9.3
R90086 biasldo.n255 biasldo.n254 9.3
R90087 biasldo.n254 biasldo.n253 9.3
R90088 biasldo.n266 biasldo.n265 9.3
R90089 biasldo.n265 biasldo.n264 9.3
R90090 biasldo.n259 biasldo.n258 9.3
R90091 biasldo.n270 biasldo.n269 9.3
R90092 biasldo.n277 biasldo.n276 9.3
R90093 biasldo.n276 biasldo.n275 9.3
R90094 biasldo.n283 biasldo.n282 9.3
R90095 biasldo.n281 biasldo.n280 9.3
R90096 biasldo.n562 biasldo.n561 9.3
R90097 biasldo.n551 biasldo.n550 9.3
R90098 biasldo.n540 biasldo.n539 9.3
R90099 biasldo.n529 biasldo.n528 9.3
R90100 biasldo.n517 biasldo.n516 9.3
R90101 biasldo.n510 biasldo.n509 9.3
R90102 biasldo.n509 biasldo.n508 9.3
R90103 biasldo.n492 biasldo.n491 9.3
R90104 biasldo.n470 biasldo.n469 9.3
R90105 biasldo.n448 biasldo.n447 9.3
R90106 biasldo.n414 biasldo.n413 9.3
R90107 biasldo.n403 biasldo.n402 9.3
R90108 biasldo.n392 biasldo.n391 9.3
R90109 biasldo.n381 biasldo.n380 9.3
R90110 biasldo.n370 biasldo.n369 9.3
R90111 biasldo.n359 biasldo.n358 9.3
R90112 biasldo.n348 biasldo.n347 9.3
R90113 biasldo.n336 biasldo.n335 9.3
R90114 biasldo.n322 biasldo.n321 9.3
R90115 biasldo.n300 biasldo.n299 9.3
R90116 biasldo.n285 biasldo.n284 9.3
R90117 biasldo.n289 biasldo.n288 9.3
R90118 biasldo.n287 biasldo.n286 9.3
R90119 biasldo.n298 biasldo.n297 9.3
R90120 biasldo.n296 biasldo.n295 9.3
R90121 biasldo.n295 biasldo.n294 9.3
R90122 biasldo.n307 biasldo.n306 9.3
R90123 biasldo.n306 biasldo.n305 9.3
R90124 biasldo.n311 biasldo.n310 9.3
R90125 biasldo.n309 biasldo.n308 9.3
R90126 biasldo.n320 biasldo.n319 9.3
R90127 biasldo.n318 biasldo.n317 9.3
R90128 biasldo.n317 biasldo.n316 9.3
R90129 biasldo.n329 biasldo.n328 9.3
R90130 biasldo.n328 biasldo.n327 9.3
R90131 biasldo.n333 biasldo.n332 9.3
R90132 biasldo.n331 biasldo.n330 9.3
R90133 biasldo.n338 biasldo.n337 9.3
R90134 biasldo.n346 biasldo.n345 9.3
R90135 biasldo.n345 biasldo.n344 9.3
R90136 biasldo.n357 biasldo.n356 9.3
R90137 biasldo.n356 biasldo.n355 9.3
R90138 biasldo.n350 biasldo.n349 9.3
R90139 biasldo.n361 biasldo.n360 9.3
R90140 biasldo.n368 biasldo.n367 9.3
R90141 biasldo.n367 biasldo.n366 9.3
R90142 biasldo.n379 biasldo.n378 9.3
R90143 biasldo.n378 biasldo.n377 9.3
R90144 biasldo.n372 biasldo.n371 9.3
R90145 biasldo.n383 biasldo.n382 9.3
R90146 biasldo.n390 biasldo.n389 9.3
R90147 biasldo.n389 biasldo.n388 9.3
R90148 biasldo.n401 biasldo.n400 9.3
R90149 biasldo.n400 biasldo.n399 9.3
R90150 biasldo.n394 biasldo.n393 9.3
R90151 biasldo.n405 biasldo.n404 9.3
R90152 biasldo.n412 biasldo.n411 9.3
R90153 biasldo.n411 biasldo.n410 9.3
R90154 biasldo.n423 biasldo.n422 9.3
R90155 biasldo.n422 biasldo.n421 9.3
R90156 biasldo.n416 biasldo.n415 9.3
R90157 biasldo.n433 biasldo.n432 9.3
R90158 biasldo.n432 biasldo.n431 9.3
R90159 biasldo.n437 biasldo.n436 9.3
R90160 biasldo.n435 biasldo.n434 9.3
R90161 biasldo.n446 biasldo.n445 9.3
R90162 biasldo.n444 biasldo.n443 9.3
R90163 biasldo.n443 biasldo.n442 9.3
R90164 biasldo.n455 biasldo.n454 9.3
R90165 biasldo.n454 biasldo.n453 9.3
R90166 biasldo.n459 biasldo.n458 9.3
R90167 biasldo.n457 biasldo.n456 9.3
R90168 biasldo.n468 biasldo.n467 9.3
R90169 biasldo.n466 biasldo.n465 9.3
R90170 biasldo.n465 biasldo.n464 9.3
R90171 biasldo.n477 biasldo.n476 9.3
R90172 biasldo.n476 biasldo.n475 9.3
R90173 biasldo.n481 biasldo.n480 9.3
R90174 biasldo.n479 biasldo.n478 9.3
R90175 biasldo.n490 biasldo.n489 9.3
R90176 biasldo.n488 biasldo.n487 9.3
R90177 biasldo.n487 biasldo.n486 9.3
R90178 biasldo.n499 biasldo.n498 9.3
R90179 biasldo.n498 biasldo.n497 9.3
R90180 biasldo.n503 biasldo.n502 9.3
R90181 biasldo.n501 biasldo.n500 9.3
R90182 biasldo.n512 biasldo.n511 9.3
R90183 biasldo.n514 biasldo.n513 9.3
R90184 biasldo.n527 biasldo.n526 9.3
R90185 biasldo.n526 biasldo.n525 9.3
R90186 biasldo.n519 biasldo.n518 9.3
R90187 biasldo.n531 biasldo.n530 9.3
R90188 biasldo.n538 biasldo.n537 9.3
R90189 biasldo.n537 biasldo.n536 9.3
R90190 biasldo.n549 biasldo.n548 9.3
R90191 biasldo.n548 biasldo.n547 9.3
R90192 biasldo.n542 biasldo.n541 9.3
R90193 biasldo.n553 biasldo.n552 9.3
R90194 biasldo.n560 biasldo.n559 9.3
R90195 biasldo.n559 biasldo.n558 9.3
R90196 biasldo.n566 biasldo.n565 9.3
R90197 biasldo.n564 biasldo.n563 9.3
R90198 biasldo.n12 biasldo.n11 9.3
R90199 biasldo.n23 biasldo.n22 9.3
R90200 biasldo.n34 biasldo.n33 9.3
R90201 biasldo.n45 biasldo.n44 9.3
R90202 biasldo.n56 biasldo.n55 9.3
R90203 biasldo.n67 biasldo.n66 9.3
R90204 biasldo.n78 biasldo.n77 9.3
R90205 biasldo.n89 biasldo.n88 9.3
R90206 biasldo.n102 biasldo.n101 9.3
R90207 biasldo.n101 biasldo.n100 9.3
R90208 biasldo.n115 biasldo.n114 9.3
R90209 biasldo.n137 biasldo.n136 9.3
R90210 biasldo.n139 biasldo.n138 9.3
R90211 biasldo.n141 biasldo.n140 9.3
R90212 biasldo.n135 biasldo.n134 9.3
R90213 biasldo.n134 biasldo.n133 9.3
R90214 biasldo.n126 biasldo.n125 9.3
R90215 biasldo.n128 biasldo.n127 9.3
R90216 biasldo.n117 biasldo.n116 9.3
R90217 biasldo.n124 biasldo.n123 9.3
R90218 biasldo.n123 biasldo.n122 9.3
R90219 biasldo.n113 biasldo.n112 9.3
R90220 biasldo.n112 biasldo.n111 9.3
R90221 biasldo.n104 biasldo.n103 9.3
R90222 biasldo.n106 biasldo.n105 9.3
R90223 biasldo.n94 biasldo.n93 9.3
R90224 biasldo.n92 biasldo.n91 9.3
R90225 biasldo.n85 biasldo.n84 9.3
R90226 biasldo.n84 biasldo.n83 9.3
R90227 biasldo.n87 biasldo.n86 9.3
R90228 biasldo.n76 biasldo.n75 9.3
R90229 biasldo.n74 biasldo.n73 9.3
R90230 biasldo.n73 biasldo.n72 9.3
R90231 biasldo.n63 biasldo.n62 9.3
R90232 biasldo.n62 biasldo.n61 9.3
R90233 biasldo.n65 biasldo.n64 9.3
R90234 biasldo.n54 biasldo.n53 9.3
R90235 biasldo.n52 biasldo.n51 9.3
R90236 biasldo.n51 biasldo.n50 9.3
R90237 biasldo.n41 biasldo.n40 9.3
R90238 biasldo.n40 biasldo.n39 9.3
R90239 biasldo.n43 biasldo.n42 9.3
R90240 biasldo.n32 biasldo.n31 9.3
R90241 biasldo.n30 biasldo.n29 9.3
R90242 biasldo.n29 biasldo.n28 9.3
R90243 biasldo.n19 biasldo.n18 9.3
R90244 biasldo.n18 biasldo.n17 9.3
R90245 biasldo.n21 biasldo.n20 9.3
R90246 biasldo.n10 biasldo.n9 9.3
R90247 biasldo.n8 biasldo.n7 9.3
R90248 biasldo.n7 biasldo.n6 9.3
R90249 biasldo.n845 biasldo.n844 9.3
R90250 biasldo.n834 biasldo.n833 9.3
R90251 biasldo.n823 biasldo.n822 9.3
R90252 biasldo.n812 biasldo.n811 9.3
R90253 biasldo.n800 biasldo.n799 9.3
R90254 biasldo.n793 biasldo.n792 9.3
R90255 biasldo.n792 biasldo.n791 9.3
R90256 biasldo.n775 biasldo.n774 9.3
R90257 biasldo.n753 biasldo.n752 9.3
R90258 biasldo.n731 biasldo.n730 9.3
R90259 biasldo.n697 biasldo.n696 9.3
R90260 biasldo.n686 biasldo.n685 9.3
R90261 biasldo.n675 biasldo.n674 9.3
R90262 biasldo.n664 biasldo.n663 9.3
R90263 biasldo.n653 biasldo.n652 9.3
R90264 biasldo.n642 biasldo.n641 9.3
R90265 biasldo.n631 biasldo.n630 9.3
R90266 biasldo.n619 biasldo.n618 9.3
R90267 biasldo.n605 biasldo.n604 9.3
R90268 biasldo.n583 biasldo.n582 9.3
R90269 biasldo.n568 biasldo.n567 9.3
R90270 biasldo.n572 biasldo.n571 9.3
R90271 biasldo.n570 biasldo.n569 9.3
R90272 biasldo.n581 biasldo.n580 9.3
R90273 biasldo.n579 biasldo.n578 9.3
R90274 biasldo.n578 biasldo.n577 9.3
R90275 biasldo.n590 biasldo.n589 9.3
R90276 biasldo.n589 biasldo.n588 9.3
R90277 biasldo.n594 biasldo.n593 9.3
R90278 biasldo.n592 biasldo.n591 9.3
R90279 biasldo.n603 biasldo.n602 9.3
R90280 biasldo.n601 biasldo.n600 9.3
R90281 biasldo.n600 biasldo.n599 9.3
R90282 biasldo.n612 biasldo.n611 9.3
R90283 biasldo.n611 biasldo.n610 9.3
R90284 biasldo.n616 biasldo.n615 9.3
R90285 biasldo.n614 biasldo.n613 9.3
R90286 biasldo.n621 biasldo.n620 9.3
R90287 biasldo.n629 biasldo.n628 9.3
R90288 biasldo.n628 biasldo.n627 9.3
R90289 biasldo.n640 biasldo.n639 9.3
R90290 biasldo.n639 biasldo.n638 9.3
R90291 biasldo.n633 biasldo.n632 9.3
R90292 biasldo.n644 biasldo.n643 9.3
R90293 biasldo.n651 biasldo.n650 9.3
R90294 biasldo.n650 biasldo.n649 9.3
R90295 biasldo.n662 biasldo.n661 9.3
R90296 biasldo.n661 biasldo.n660 9.3
R90297 biasldo.n655 biasldo.n654 9.3
R90298 biasldo.n666 biasldo.n665 9.3
R90299 biasldo.n673 biasldo.n672 9.3
R90300 biasldo.n672 biasldo.n671 9.3
R90301 biasldo.n684 biasldo.n683 9.3
R90302 biasldo.n683 biasldo.n682 9.3
R90303 biasldo.n677 biasldo.n676 9.3
R90304 biasldo.n688 biasldo.n687 9.3
R90305 biasldo.n695 biasldo.n694 9.3
R90306 biasldo.n694 biasldo.n693 9.3
R90307 biasldo.n706 biasldo.n705 9.3
R90308 biasldo.n705 biasldo.n704 9.3
R90309 biasldo.n699 biasldo.n698 9.3
R90310 biasldo.n716 biasldo.n715 9.3
R90311 biasldo.n715 biasldo.n714 9.3
R90312 biasldo.n720 biasldo.n719 9.3
R90313 biasldo.n718 biasldo.n717 9.3
R90314 biasldo.n729 biasldo.n728 9.3
R90315 biasldo.n727 biasldo.n726 9.3
R90316 biasldo.n726 biasldo.n725 9.3
R90317 biasldo.n738 biasldo.n737 9.3
R90318 biasldo.n737 biasldo.n736 9.3
R90319 biasldo.n742 biasldo.n741 9.3
R90320 biasldo.n740 biasldo.n739 9.3
R90321 biasldo.n751 biasldo.n750 9.3
R90322 biasldo.n749 biasldo.n748 9.3
R90323 biasldo.n748 biasldo.n747 9.3
R90324 biasldo.n760 biasldo.n759 9.3
R90325 biasldo.n759 biasldo.n758 9.3
R90326 biasldo.n764 biasldo.n763 9.3
R90327 biasldo.n762 biasldo.n761 9.3
R90328 biasldo.n773 biasldo.n772 9.3
R90329 biasldo.n771 biasldo.n770 9.3
R90330 biasldo.n770 biasldo.n769 9.3
R90331 biasldo.n782 biasldo.n781 9.3
R90332 biasldo.n781 biasldo.n780 9.3
R90333 biasldo.n786 biasldo.n785 9.3
R90334 biasldo.n784 biasldo.n783 9.3
R90335 biasldo.n795 biasldo.n794 9.3
R90336 biasldo.n797 biasldo.n796 9.3
R90337 biasldo.n810 biasldo.n809 9.3
R90338 biasldo.n809 biasldo.n808 9.3
R90339 biasldo.n802 biasldo.n801 9.3
R90340 biasldo.n814 biasldo.n813 9.3
R90341 biasldo.n821 biasldo.n820 9.3
R90342 biasldo.n820 biasldo.n819 9.3
R90343 biasldo.n832 biasldo.n831 9.3
R90344 biasldo.n831 biasldo.n830 9.3
R90345 biasldo.n825 biasldo.n824 9.3
R90346 biasldo.n836 biasldo.n835 9.3
R90347 biasldo.n843 biasldo.n842 9.3
R90348 biasldo.n842 biasldo.n841 9.3
R90349 biasldo.n849 biasldo.n848 9.3
R90350 biasldo.n847 biasldo.n846 9.3
R90351 biasldo.n856 biasldo.n855 9.3
R90352 biasldo.n863 biasldo.n862 9.3
R90353 biasldo.n866 biasldo.n865 9.3
R90354 biasldo.n861 biasldo.n860 9.3
R90355 biasldo.n859 biasldo.n858 9.3
R90356 biasldo.n854 biasldo.n853 9.3
R90357 biasldo.n425 biasldo.n424 8.764
R90358 biasldo.n708 biasldo.n707 8.764
R90359 biasldo.n610 biasldo.n609 8.763
R90360 biasldo.n627 biasldo.n626 8.763
R90361 biasldo.n791 biasldo.n790 8.763
R90362 biasldo.n808 biasldo.n807 8.763
R90363 biasldo.n327 biasldo.n326 8.763
R90364 biasldo.n344 biasldo.n343 8.763
R90365 biasldo.n508 biasldo.n507 8.763
R90366 biasldo.n525 biasldo.n524 8.763
R90367 biasldo.n225 biasldo.n224 8.763
R90368 biasldo.n242 biasldo.n241 8.763
R90369 biasldo.n100 biasldo.n98 8.763
R90370 biasldo.n83 biasldo.n82 8.763
R90371 biasldo.n703 biasldo.n702 8.215
R90372 biasldo.n713 biasldo.n712 8.215
R90373 biasldo.n420 biasldo.n419 8.215
R90374 biasldo.n430 biasldo.n429 8.215
R90375 biasldo.n147 biasldo.n146 8.215
R90376 biasldo.n5 biasldo.n4 8.215
R90377 biasldo.n599 biasldo.n598 7.668
R90378 biasldo.n638 biasldo.n637 7.668
R90379 biasldo.n780 biasldo.n779 7.668
R90380 biasldo.n819 biasldo.n818 7.668
R90381 biasldo.n316 biasldo.n315 7.668
R90382 biasldo.n355 biasldo.n354 7.668
R90383 biasldo.n497 biasldo.n496 7.668
R90384 biasldo.n536 biasldo.n535 7.668
R90385 biasldo.n214 biasldo.n213 7.668
R90386 biasldo.n253 biasldo.n252 7.668
R90387 biasldo.n111 biasldo.n110 7.668
R90388 biasldo.n72 biasldo.n71 7.668
R90389 biasldo.n692 biasldo.n691 7.12
R90390 biasldo.n724 biasldo.n723 7.12
R90391 biasldo.n409 biasldo.n408 7.12
R90392 biasldo.n441 biasldo.n440 7.12
R90393 biasldo.n158 biasldo.n157 7.12
R90394 biasldo.n16 biasldo.n15 7.12
R90395 biasldo.n1 biasldo.n0 6.915
R90396 biasldo.n143 biasldo.n142 6.914
R90397 biasldo.n588 biasldo.n587 6.572
R90398 biasldo.n649 biasldo.n648 6.572
R90399 biasldo.n769 biasldo.n768 6.572
R90400 biasldo.n830 biasldo.n829 6.572
R90401 biasldo.n305 biasldo.n304 6.572
R90402 biasldo.n366 biasldo.n365 6.572
R90403 biasldo.n486 biasldo.n485 6.572
R90404 biasldo.n547 biasldo.n546 6.572
R90405 biasldo.n203 biasldo.n202 6.572
R90406 biasldo.n264 biasldo.n263 6.572
R90407 biasldo.n122 biasldo.n121 6.572
R90408 biasldo.n61 biasldo.n60 6.572
R90409 biasldo.n681 biasldo.n680 6.025
R90410 biasldo.n735 biasldo.n734 6.025
R90411 biasldo.n398 biasldo.n397 6.025
R90412 biasldo.n452 biasldo.n451 6.025
R90413 biasldo.n169 biasldo.n168 6.025
R90414 biasldo.n27 biasldo.n26 6.025
R90415 biasldo.n611 biasldo.n607 6.023
R90416 biasldo.n628 biasldo.n623 6.023
R90417 biasldo.n792 biasldo.n788 6.023
R90418 biasldo.n809 biasldo.n804 6.023
R90419 biasldo.n328 biasldo.n324 6.023
R90420 biasldo.n345 biasldo.n340 6.023
R90421 biasldo.n509 biasldo.n505 6.023
R90422 biasldo.n526 biasldo.n521 6.023
R90423 biasldo.n226 biasldo.n222 6.023
R90424 biasldo.n243 biasldo.n238 6.023
R90425 biasldo.n101 biasldo.n96 6.023
R90426 biasldo.n84 biasldo.n80 6.023
R90427 biasldo.n701 biasldo.n700 5.647
R90428 biasldo.n711 biasldo.n710 5.647
R90429 biasldo.n418 biasldo.n417 5.647
R90430 biasldo.n428 biasldo.n427 5.647
R90431 biasldo.n145 biasldo.n144 5.647
R90432 biasldo.n3 biasldo.n2 5.647
R90433 biasldo.n577 biasldo.n576 5.477
R90434 biasldo.n660 biasldo.n659 5.477
R90435 biasldo.n758 biasldo.n757 5.477
R90436 biasldo.n841 biasldo.n840 5.477
R90437 biasldo.n294 biasldo.n293 5.477
R90438 biasldo.n377 biasldo.n376 5.477
R90439 biasldo.n475 biasldo.n474 5.477
R90440 biasldo.n558 biasldo.n557 5.477
R90441 biasldo.n192 biasldo.n191 5.477
R90442 biasldo.n275 biasldo.n274 5.477
R90443 biasldo.n133 biasldo.n132 5.477
R90444 biasldo.n50 biasldo.n49 5.477
R90445 biasldo.n868 biasldo.n867 5.343
R90446 biasldo.n852 biasldo.n851 5.28
R90447 biasldo.n600 biasldo.n596 5.27
R90448 biasldo.n639 biasldo.n635 5.27
R90449 biasldo.n781 biasldo.n777 5.27
R90450 biasldo.n820 biasldo.n816 5.27
R90451 biasldo.n317 biasldo.n313 5.27
R90452 biasldo.n356 biasldo.n352 5.27
R90453 biasldo.n498 biasldo.n494 5.27
R90454 biasldo.n537 biasldo.n533 5.27
R90455 biasldo.n215 biasldo.n211 5.27
R90456 biasldo.n254 biasldo.n250 5.27
R90457 biasldo.n112 biasldo.n108 5.27
R90458 biasldo.n73 biasldo.n69 5.27
R90459 biasldo.n670 biasldo.n669 4.929
R90460 biasldo.n746 biasldo.n745 4.929
R90461 biasldo.n387 biasldo.n386 4.929
R90462 biasldo.n463 biasldo.n462 4.929
R90463 biasldo.n180 biasldo.n179 4.929
R90464 biasldo.n38 biasldo.n37 4.929
R90465 biasldo.n690 biasldo.n689 4.894
R90466 biasldo.n722 biasldo.n721 4.894
R90467 biasldo.n407 biasldo.n406 4.894
R90468 biasldo.n439 biasldo.n438 4.894
R90469 biasldo.n156 biasldo.n155 4.894
R90470 biasldo.n14 biasldo.n13 4.894
R90471 biasldo.n426 biasldo.n425 4.65
R90472 biasldo.n709 biasldo.n708 4.65
R90473 biasldo.n869 biasldo.n868 4.65
R90474 biasldo.n589 biasldo.n585 4.517
R90475 biasldo.n650 biasldo.n646 4.517
R90476 biasldo.n770 biasldo.n766 4.517
R90477 biasldo.n831 biasldo.n827 4.517
R90478 biasldo.n306 biasldo.n302 4.517
R90479 biasldo.n367 biasldo.n363 4.517
R90480 biasldo.n487 biasldo.n483 4.517
R90481 biasldo.n548 biasldo.n544 4.517
R90482 biasldo.n204 biasldo.n200 4.517
R90483 biasldo.n265 biasldo.n261 4.517
R90484 biasldo.n123 biasldo.n119 4.517
R90485 biasldo.n62 biasldo.n58 4.517
R90486 biasldo.n886 biasldo.n872 4.47
R90487 biasldo.n671 biasldo.n670 4.381
R90488 biasldo.n747 biasldo.n746 4.381
R90489 biasldo.n388 biasldo.n387 4.381
R90490 biasldo.n464 biasldo.n463 4.381
R90491 biasldo.n181 biasldo.n180 4.381
R90492 biasldo.n39 biasldo.n38 4.381
R90493 biasldo.n872 biasldo.n871 4.214
R90494 biasldo.n679 biasldo.n678 4.141
R90495 biasldo.n733 biasldo.n732 4.141
R90496 biasldo.n396 biasldo.n395 4.141
R90497 biasldo.n450 biasldo.n449 4.141
R90498 biasldo.n167 biasldo.n166 4.141
R90499 biasldo.n25 biasldo.n24 4.141
R90500 biasldo.n576 biasldo.n575 3.834
R90501 biasldo.n659 biasldo.n658 3.834
R90502 biasldo.n757 biasldo.n756 3.834
R90503 biasldo.n840 biasldo.n839 3.834
R90504 biasldo.n293 biasldo.n292 3.834
R90505 biasldo.n376 biasldo.n375 3.834
R90506 biasldo.n474 biasldo.n473 3.834
R90507 biasldo.n557 biasldo.n556 3.834
R90508 biasldo.n191 biasldo.n190 3.834
R90509 biasldo.n274 biasldo.n273 3.834
R90510 biasldo.n132 biasldo.n131 3.834
R90511 biasldo.n49 biasldo.n48 3.834
R90512 biasldo.n578 biasldo.n574 3.764
R90513 biasldo.n661 biasldo.n657 3.764
R90514 biasldo.n759 biasldo.n755 3.764
R90515 biasldo.n842 biasldo.n838 3.764
R90516 biasldo.n295 biasldo.n291 3.764
R90517 biasldo.n378 biasldo.n374 3.764
R90518 biasldo.n476 biasldo.n472 3.764
R90519 biasldo.n559 biasldo.n555 3.764
R90520 biasldo.n193 biasldo.n189 3.764
R90521 biasldo.n276 biasldo.n272 3.764
R90522 biasldo.n134 biasldo.n130 3.764
R90523 biasldo.n51 biasldo.n47 3.764
R90524 biasldo.n150 biasldo.n143 3.409
R90525 biasldo.n8 biasldo.n1 3.408
R90526 biasldo.n668 biasldo.n667 3.388
R90527 biasldo.n744 biasldo.n743 3.388
R90528 biasldo.n385 biasldo.n384 3.388
R90529 biasldo.n461 biasldo.n460 3.388
R90530 biasldo.n178 biasldo.n177 3.388
R90531 biasldo.n36 biasldo.n35 3.388
R90532 biasldo.n883 biasldo.t3 3.306
R90533 biasldo.n883 biasldo.t1 3.306
R90534 biasldo.n682 biasldo.n681 3.286
R90535 biasldo.n736 biasldo.n735 3.286
R90536 biasldo.n399 biasldo.n398 3.286
R90537 biasldo.n453 biasldo.n452 3.286
R90538 biasldo.n170 biasldo.n169 3.286
R90539 biasldo.n28 biasldo.n27 3.286
R90540 biasldo.n672 biasldo.n668 3.011
R90541 biasldo.n748 biasldo.n744 3.011
R90542 biasldo.n389 biasldo.n385 3.011
R90543 biasldo.n465 biasldo.n461 3.011
R90544 biasldo.n182 biasldo.n178 3.011
R90545 biasldo.n40 biasldo.n36 3.011
R90546 biasldo.n587 biasldo.n586 2.738
R90547 biasldo.n648 biasldo.n647 2.738
R90548 biasldo.n768 biasldo.n767 2.738
R90549 biasldo.n829 biasldo.n828 2.738
R90550 biasldo.n304 biasldo.n303 2.738
R90551 biasldo.n365 biasldo.n364 2.738
R90552 biasldo.n485 biasldo.n484 2.738
R90553 biasldo.n546 biasldo.n545 2.738
R90554 biasldo.n202 biasldo.n201 2.738
R90555 biasldo.n263 biasldo.n262 2.738
R90556 biasldo.n121 biasldo.n120 2.738
R90557 biasldo.n60 biasldo.n59 2.738
R90558 biasldo.n574 biasldo.n573 2.635
R90559 biasldo.n657 biasldo.n656 2.635
R90560 biasldo.n755 biasldo.n754 2.635
R90561 biasldo.n838 biasldo.n837 2.635
R90562 biasldo.n291 biasldo.n290 2.635
R90563 biasldo.n374 biasldo.n373 2.635
R90564 biasldo.n472 biasldo.n471 2.635
R90565 biasldo.n555 biasldo.n554 2.635
R90566 biasldo.n189 biasldo.n188 2.635
R90567 biasldo.n272 biasldo.n271 2.635
R90568 biasldo.n130 biasldo.n129 2.635
R90569 biasldo.n47 biasldo.n46 2.635
R90570 biasldo.n683 biasldo.n679 2.258
R90571 biasldo.n737 biasldo.n733 2.258
R90572 biasldo.n400 biasldo.n396 2.258
R90573 biasldo.n454 biasldo.n450 2.258
R90574 biasldo.n171 biasldo.n167 2.258
R90575 biasldo.n29 biasldo.n25 2.258
R90576 biasldo.n693 biasldo.n692 2.19
R90577 biasldo.n725 biasldo.n724 2.19
R90578 biasldo.n410 biasldo.n409 2.19
R90579 biasldo.n442 biasldo.n441 2.19
R90580 biasldo.n159 biasldo.n158 2.19
R90581 biasldo.n17 biasldo.n16 2.19
R90582 biasldo.n585 biasldo.n584 1.882
R90583 biasldo.n646 biasldo.n645 1.882
R90584 biasldo.n766 biasldo.n765 1.882
R90585 biasldo.n827 biasldo.n826 1.882
R90586 biasldo.n302 biasldo.n301 1.882
R90587 biasldo.n363 biasldo.n362 1.882
R90588 biasldo.n483 biasldo.n482 1.882
R90589 biasldo.n544 biasldo.n543 1.882
R90590 biasldo.n200 biasldo.n199 1.882
R90591 biasldo.n261 biasldo.n260 1.882
R90592 biasldo.n119 biasldo.n118 1.882
R90593 biasldo.n58 biasldo.n57 1.882
R90594 biasldo.n598 biasldo.n597 1.643
R90595 biasldo.n637 biasldo.n636 1.643
R90596 biasldo.n779 biasldo.n778 1.643
R90597 biasldo.n818 biasldo.n817 1.643
R90598 biasldo.n315 biasldo.n314 1.643
R90599 biasldo.n354 biasldo.n353 1.643
R90600 biasldo.n496 biasldo.n495 1.643
R90601 biasldo.n535 biasldo.n534 1.643
R90602 biasldo.n213 biasldo.n212 1.643
R90603 biasldo.n252 biasldo.n251 1.643
R90604 biasldo.n110 biasldo.n109 1.643
R90605 biasldo.n71 biasldo.n70 1.643
R90606 biasldo.n889 biasldo.n886 1.517
R90607 biasldo.n694 biasldo.n690 1.505
R90608 biasldo.n726 biasldo.n722 1.505
R90609 biasldo.n411 biasldo.n407 1.505
R90610 biasldo.n443 biasldo.n439 1.505
R90611 biasldo.n160 biasldo.n156 1.505
R90612 biasldo.n18 biasldo.n14 1.505
R90613 biasldo.n884 biasldo.n883 1.467
R90614 biasldo.n596 biasldo.n595 1.129
R90615 biasldo.n635 biasldo.n634 1.129
R90616 biasldo.n777 biasldo.n776 1.129
R90617 biasldo.n816 biasldo.n815 1.129
R90618 biasldo.n313 biasldo.n312 1.129
R90619 biasldo.n352 biasldo.n351 1.129
R90620 biasldo.n494 biasldo.n493 1.129
R90621 biasldo.n533 biasldo.n532 1.129
R90622 biasldo.n211 biasldo.n210 1.129
R90623 biasldo.n250 biasldo.n249 1.129
R90624 biasldo.n108 biasldo.n107 1.129
R90625 biasldo.n69 biasldo.n68 1.129
R90626 biasldo.n704 biasldo.n703 1.095
R90627 biasldo.n714 biasldo.n713 1.095
R90628 biasldo.n421 biasldo.n420 1.095
R90629 biasldo.n431 biasldo.n430 1.095
R90630 biasldo.n148 biasldo.n147 1.095
R90631 biasldo.n6 biasldo.n5 1.095
R90632 biasldo.n705 biasldo.n701 0.752
R90633 biasldo.n715 biasldo.n711 0.752
R90634 biasldo.n422 biasldo.n418 0.752
R90635 biasldo.n432 biasldo.n428 0.752
R90636 biasldo.n149 biasldo.n145 0.752
R90637 biasldo.n7 biasldo.n3 0.752
R90638 biasldo.n885 biasldo.n884 0.562
R90639 biasldo.n609 biasldo.n608 0.547
R90640 biasldo.n626 biasldo.n625 0.547
R90641 biasldo.n790 biasldo.n789 0.547
R90642 biasldo.n807 biasldo.n806 0.547
R90643 biasldo.n326 biasldo.n325 0.547
R90644 biasldo.n343 biasldo.n342 0.547
R90645 biasldo.n507 biasldo.n506 0.547
R90646 biasldo.n524 biasldo.n523 0.547
R90647 biasldo.n224 biasldo.n223 0.547
R90648 biasldo.n241 biasldo.n240 0.547
R90649 biasldo.n98 biasldo.n97 0.547
R90650 biasldo.n82 biasldo.n81 0.547
R90651 biasldo.n858 biasldo.n857 0.461
R90652 biasldo.n865 biasldo.n864 0.43
R90653 biasldo.n607 biasldo.n606 0.376
R90654 biasldo.n623 biasldo.n622 0.376
R90655 biasldo.n788 biasldo.n787 0.376
R90656 biasldo.n804 biasldo.n803 0.376
R90657 biasldo.n324 biasldo.n323 0.376
R90658 biasldo.n340 biasldo.n339 0.376
R90659 biasldo.n505 biasldo.n504 0.376
R90660 biasldo.n521 biasldo.n520 0.376
R90661 biasldo.n222 biasldo.n221 0.376
R90662 biasldo.n238 biasldo.n237 0.376
R90663 biasldo.n96 biasldo.n95 0.376
R90664 biasldo.n80 biasldo.n79 0.376
R90665 biasldo.n285 biasldo.n283 0.323
R90666 biasldo.n568 biasldo.n566 0.323
R90667 ldomc_0.bias ldomc_0.otaldom_0.bias 0.285
R90668 biasldo.n887 ldomc_0.bias 0.251
R90669 biasldo.n852 biasldo.n850 0.144
R90670 biasldo.n234 biasldo.n231 0.128
R90671 biasldo.n336 biasldo.n333 0.128
R90672 biasldo.n426 biasldo.n423 0.128
R90673 biasldo.n433 biasldo.n426 0.128
R90674 biasldo.n517 biasldo.n514 0.128
R90675 biasldo.n92 biasldo.n89 0.128
R90676 biasldo.n619 biasldo.n616 0.128
R90677 biasldo.n709 biasldo.n706 0.128
R90678 biasldo.n716 biasldo.n709 0.128
R90679 biasldo.n800 biasldo.n797 0.128
R90680 biasldo.n161 biasldo.n154 0.097
R90681 biasldo.n172 biasldo.n165 0.097
R90682 biasldo.n183 biasldo.n176 0.097
R90683 biasldo.n194 biasldo.n187 0.097
R90684 biasldo.n205 biasldo.n198 0.097
R90685 biasldo.n216 biasldo.n209 0.097
R90686 biasldo.n227 biasldo.n220 0.097
R90687 biasldo.n246 biasldo.n244 0.097
R90688 biasldo.n257 biasldo.n255 0.097
R90689 biasldo.n268 biasldo.n266 0.097
R90690 biasldo.n279 biasldo.n277 0.097
R90691 biasldo.n296 biasldo.n289 0.097
R90692 biasldo.n307 biasldo.n300 0.097
R90693 biasldo.n318 biasldo.n311 0.097
R90694 biasldo.n329 biasldo.n322 0.097
R90695 biasldo.n348 biasldo.n346 0.097
R90696 biasldo.n359 biasldo.n357 0.097
R90697 biasldo.n370 biasldo.n368 0.097
R90698 biasldo.n381 biasldo.n379 0.097
R90699 biasldo.n392 biasldo.n390 0.097
R90700 biasldo.n403 biasldo.n401 0.097
R90701 biasldo.n414 biasldo.n412 0.097
R90702 biasldo.n444 biasldo.n437 0.097
R90703 biasldo.n455 biasldo.n448 0.097
R90704 biasldo.n466 biasldo.n459 0.097
R90705 biasldo.n477 biasldo.n470 0.097
R90706 biasldo.n488 biasldo.n481 0.097
R90707 biasldo.n499 biasldo.n492 0.097
R90708 biasldo.n510 biasldo.n503 0.097
R90709 biasldo.n529 biasldo.n527 0.097
R90710 biasldo.n540 biasldo.n538 0.097
R90711 biasldo.n551 biasldo.n549 0.097
R90712 biasldo.n562 biasldo.n560 0.097
R90713 biasldo.n137 biasldo.n135 0.097
R90714 biasldo.n126 biasldo.n124 0.097
R90715 biasldo.n115 biasldo.n113 0.097
R90716 biasldo.n104 biasldo.n102 0.097
R90717 biasldo.n85 biasldo.n78 0.097
R90718 biasldo.n74 biasldo.n67 0.097
R90719 biasldo.n63 biasldo.n56 0.097
R90720 biasldo.n52 biasldo.n45 0.097
R90721 biasldo.n41 biasldo.n34 0.097
R90722 biasldo.n30 biasldo.n23 0.097
R90723 biasldo.n19 biasldo.n12 0.097
R90724 biasldo.n579 biasldo.n572 0.097
R90725 biasldo.n590 biasldo.n583 0.097
R90726 biasldo.n601 biasldo.n594 0.097
R90727 biasldo.n612 biasldo.n605 0.097
R90728 biasldo.n631 biasldo.n629 0.097
R90729 biasldo.n642 biasldo.n640 0.097
R90730 biasldo.n653 biasldo.n651 0.097
R90731 biasldo.n664 biasldo.n662 0.097
R90732 biasldo.n675 biasldo.n673 0.097
R90733 biasldo.n686 biasldo.n684 0.097
R90734 biasldo.n697 biasldo.n695 0.097
R90735 biasldo.n727 biasldo.n720 0.097
R90736 biasldo.n738 biasldo.n731 0.097
R90737 biasldo.n749 biasldo.n742 0.097
R90738 biasldo.n760 biasldo.n753 0.097
R90739 biasldo.n771 biasldo.n764 0.097
R90740 biasldo.n782 biasldo.n775 0.097
R90741 biasldo.n793 biasldo.n786 0.097
R90742 biasldo.n812 biasldo.n810 0.097
R90743 biasldo.n823 biasldo.n821 0.097
R90744 biasldo.n834 biasldo.n832 0.097
R90745 biasldo.n845 biasldo.n843 0.097
R90746 biasldo.n886 biasldo.n876 0.088
R90747 biasldo.n854 biasldo.n852 0.084
R90748 biasldo.n850 biasldo.n141 0.077
R90749 biasldo.n886 biasldo.n881 0.075
R90750 biasldo.n861 biasldo.n859 0.073
R90751 biasldo.n869 biasldo.n866 0.073
R90752 biasldo.n878 biasldo.n877 0.071
R90753 biasldo.n850 biasldo.n849 0.069
R90754 biasldo.n874 biasldo.n873 0.065
R90755 biasldo biasldo.n889 0.061
R90756 biasldo.n886 biasldo.n870 0.033
R90757 biasldo.n886 biasldo.n885 0.033
R90758 biasldo.n229 biasldo.n227 0.029
R90759 biasldo.n244 biasldo.n236 0.029
R90760 biasldo.n331 biasldo.n329 0.029
R90761 biasldo.n346 biasldo.n338 0.029
R90762 biasldo.n512 biasldo.n510 0.029
R90763 biasldo.n527 biasldo.n519 0.029
R90764 biasldo.n102 biasldo.n94 0.029
R90765 biasldo.n87 biasldo.n85 0.029
R90766 biasldo.n614 biasldo.n612 0.029
R90767 biasldo.n629 biasldo.n621 0.029
R90768 biasldo.n795 biasldo.n793 0.029
R90769 biasldo.n810 biasldo.n802 0.029
R90770 biasldo.n154 biasldo.n152 0.027
R90771 biasldo.n416 biasldo.n414 0.027
R90772 biasldo.n437 biasldo.n435 0.027
R90773 biasldo.n12 biasldo.n10 0.027
R90774 biasldo.n699 biasldo.n697 0.027
R90775 biasldo.n720 biasldo.n718 0.027
R90776 biasldo.n218 biasldo.n216 0.025
R90777 biasldo.n255 biasldo.n248 0.025
R90778 biasldo.n320 biasldo.n318 0.025
R90779 biasldo.n357 biasldo.n350 0.025
R90780 biasldo.n501 biasldo.n499 0.025
R90781 biasldo.n538 biasldo.n531 0.025
R90782 biasldo.n113 biasldo.n106 0.025
R90783 biasldo.n76 biasldo.n74 0.025
R90784 biasldo.n603 biasldo.n601 0.025
R90785 biasldo.n640 biasldo.n633 0.025
R90786 biasldo.n784 biasldo.n782 0.025
R90787 biasldo.n821 biasldo.n814 0.025
R90788 biasldo.n165 biasldo.n163 0.023
R90789 biasldo.n405 biasldo.n403 0.023
R90790 biasldo.n448 biasldo.n446 0.023
R90791 biasldo.n23 biasldo.n21 0.023
R90792 biasldo.n688 biasldo.n686 0.023
R90793 biasldo.n731 biasldo.n729 0.023
R90794 biasldo.n207 biasldo.n205 0.022
R90795 biasldo.n266 biasldo.n259 0.022
R90796 biasldo.n309 biasldo.n307 0.022
R90797 biasldo.n368 biasldo.n361 0.022
R90798 biasldo.n490 biasldo.n488 0.022
R90799 biasldo.n549 biasldo.n542 0.022
R90800 biasldo.n124 biasldo.n117 0.022
R90801 biasldo.n65 biasldo.n63 0.022
R90802 biasldo.n592 biasldo.n590 0.022
R90803 biasldo.n651 biasldo.n644 0.022
R90804 biasldo.n773 biasldo.n771 0.022
R90805 biasldo.n832 biasldo.n825 0.022
R90806 biasldo.n176 biasldo.n174 0.02
R90807 biasldo.n394 biasldo.n392 0.02
R90808 biasldo.n459 biasldo.n457 0.02
R90809 biasldo.n34 biasldo.n32 0.02
R90810 biasldo.n677 biasldo.n675 0.02
R90811 biasldo.n742 biasldo.n740 0.02
R90812 biasldo.n196 biasldo.n194 0.018
R90813 biasldo.n277 biasldo.n270 0.018
R90814 biasldo.n298 biasldo.n296 0.018
R90815 biasldo.n379 biasldo.n372 0.018
R90816 biasldo.n479 biasldo.n477 0.018
R90817 biasldo.n560 biasldo.n553 0.018
R90818 biasldo.n135 biasldo.n128 0.018
R90819 biasldo.n54 biasldo.n52 0.018
R90820 biasldo.n581 biasldo.n579 0.018
R90821 biasldo.n662 biasldo.n655 0.018
R90822 biasldo.n762 biasldo.n760 0.018
R90823 biasldo.n843 biasldo.n836 0.018
R90824 biasldo.n187 biasldo.n185 0.016
R90825 biasldo.n281 biasldo.n279 0.016
R90826 biasldo.n289 biasldo.n287 0.016
R90827 biasldo.n383 biasldo.n381 0.016
R90828 biasldo.n470 biasldo.n468 0.016
R90829 biasldo.n564 biasldo.n562 0.016
R90830 biasldo.n139 biasldo.n137 0.016
R90831 biasldo.n45 biasldo.n43 0.016
R90832 biasldo.n572 biasldo.n570 0.016
R90833 biasldo.n666 biasldo.n664 0.016
R90834 biasldo.n753 biasldo.n751 0.016
R90835 biasldo.n847 biasldo.n845 0.016
R90836 biasldo.n859 biasldo.n856 0.015
R90837 biasldo.n886 biasldo.n878 0.014
R90838 biasldo.n881 biasldo.n880 0.014
R90839 biasldo.n185 biasldo.n183 0.014
R90840 biasldo.n283 biasldo.n281 0.014
R90841 biasldo.n287 biasldo.n285 0.014
R90842 biasldo.n390 biasldo.n383 0.014
R90843 biasldo.n468 biasldo.n466 0.014
R90844 biasldo.n566 biasldo.n564 0.014
R90845 biasldo.n141 biasldo.n139 0.014
R90846 biasldo.n43 biasldo.n41 0.014
R90847 biasldo.n570 biasldo.n568 0.014
R90848 biasldo.n673 biasldo.n666 0.014
R90849 biasldo.n751 biasldo.n749 0.014
R90850 biasldo.n849 biasldo.n847 0.014
R90851 biasldo.n889 biasldo.n888 0.014
R90852 biasldo.n886 biasldo.n874 0.013
R90853 biasldo.n198 biasldo.n196 0.012
R90854 biasldo.n270 biasldo.n268 0.012
R90855 biasldo.n300 biasldo.n298 0.012
R90856 biasldo.n372 biasldo.n370 0.012
R90857 biasldo.n481 biasldo.n479 0.012
R90858 biasldo.n553 biasldo.n551 0.012
R90859 biasldo.n128 biasldo.n126 0.012
R90860 biasldo.n56 biasldo.n54 0.012
R90861 biasldo.n583 biasldo.n581 0.012
R90862 biasldo.n655 biasldo.n653 0.012
R90863 biasldo.n764 biasldo.n762 0.012
R90864 biasldo.n836 biasldo.n834 0.012
R90865 biasldo.n866 biasldo.n863 0.012
R90866 biasldo.n174 biasldo.n172 0.011
R90867 biasldo.n401 biasldo.n394 0.011
R90868 biasldo.n457 biasldo.n455 0.011
R90869 biasldo.n32 biasldo.n30 0.011
R90870 biasldo.n684 biasldo.n677 0.011
R90871 biasldo.n740 biasldo.n738 0.011
R90872 biasldo.n863 biasldo.n861 0.011
R90873 biasldo.n888 biasldo.n887 0.011
R90874 biasldo.n209 biasldo.n207 0.009
R90875 biasldo.n259 biasldo.n257 0.009
R90876 biasldo.n311 biasldo.n309 0.009
R90877 biasldo.n361 biasldo.n359 0.009
R90878 biasldo.n492 biasldo.n490 0.009
R90879 biasldo.n542 biasldo.n540 0.009
R90880 biasldo.n117 biasldo.n115 0.009
R90881 biasldo.n67 biasldo.n65 0.009
R90882 biasldo.n594 biasldo.n592 0.009
R90883 biasldo.n644 biasldo.n642 0.009
R90884 biasldo.n775 biasldo.n773 0.009
R90885 biasldo.n825 biasldo.n823 0.009
R90886 biasldo.n886 biasldo.n869 0.009
R90887 biasldo.n876 biasldo.n875 0.009
R90888 biasldo.n885 biasldo.n882 0.008
R90889 biasldo.n856 biasldo.n854 0.008
R90890 biasldo.n163 biasldo.n161 0.007
R90891 biasldo.n412 biasldo.n405 0.007
R90892 biasldo.n446 biasldo.n444 0.007
R90893 biasldo.n21 biasldo.n19 0.007
R90894 biasldo.n695 biasldo.n688 0.007
R90895 biasldo.n729 biasldo.n727 0.007
R90896 biasldo.n220 biasldo.n218 0.005
R90897 biasldo.n248 biasldo.n246 0.005
R90898 biasldo.n322 biasldo.n320 0.005
R90899 biasldo.n350 biasldo.n348 0.005
R90900 biasldo.n503 biasldo.n501 0.005
R90901 biasldo.n531 biasldo.n529 0.005
R90902 biasldo.n106 biasldo.n104 0.005
R90903 biasldo.n78 biasldo.n76 0.005
R90904 biasldo.n605 biasldo.n603 0.005
R90905 biasldo.n633 biasldo.n631 0.005
R90906 biasldo.n786 biasldo.n784 0.005
R90907 biasldo.n814 biasldo.n812 0.005
R90908 biasldo.n152 biasldo.n150 0.003
R90909 biasldo.n423 biasldo.n416 0.003
R90910 biasldo.n435 biasldo.n433 0.003
R90911 biasldo.n10 biasldo.n8 0.003
R90912 biasldo.n706 biasldo.n699 0.003
R90913 biasldo.n718 biasldo.n716 0.003
R90914 biasldo.n231 biasldo.n229 0.001
R90915 biasldo.n236 biasldo.n234 0.001
R90916 biasldo.n333 biasldo.n331 0.001
R90917 biasldo.n338 biasldo.n336 0.001
R90918 biasldo.n514 biasldo.n512 0.001
R90919 biasldo.n519 biasldo.n517 0.001
R90920 biasldo.n94 biasldo.n92 0.001
R90921 biasldo.n89 biasldo.n87 0.001
R90922 biasldo.n616 biasldo.n614 0.001
R90923 biasldo.n621 biasldo.n619 0.001
R90924 biasldo.n797 biasldo.n795 0.001
R90925 biasldo.n802 biasldo.n800 0.001
R90926 ldomc_0.otaldom_0.pcascodeupm_0.o2.n7 ldomc_0.otaldom_0.pcascodeupm_0.o2.t6 13.847
R90927 ldomc_0.otaldom_0.pcascodeupm_0.o2.n7 ldomc_0.otaldom_0.pcascodeupm_0.o2.t4 13.847
R90928 ldomc_0.otaldom_0.pcascodeupm_0.o2.n9 ldomc_0.otaldom_0.pcascodeupm_0.o2.t1 13.847
R90929 ldomc_0.otaldom_0.pcascodeupm_0.o2.n9 ldomc_0.otaldom_0.pcascodeupm_0.o2.t2 13.847
R90930 ldomc_0.otaldom_0.pcascodeupm_0.o2.n25 ldomc_0.otaldom_0.pcascodeupm_0.o2.t5 13.847
R90931 ldomc_0.otaldom_0.pcascodeupm_0.o2.n25 ldomc_0.otaldom_0.pcascodeupm_0.o2.t3 13.847
R90932 ldomc_0.otaldom_0.pcascodeupm_0.o2.n15 ldomc_0.otaldom_0.pcascodeupm_0.o2.t12 13.847
R90933 ldomc_0.otaldom_0.pcascodeupm_0.o2.n15 ldomc_0.otaldom_0.pcascodeupm_0.o2.t9 13.847
R90934 ldomc_0.otaldom_0.pcascodeupm_0.o2.n14 ldomc_0.otaldom_0.pcascodeupm_0.o2.t14 13.847
R90935 ldomc_0.otaldom_0.pcascodeupm_0.o2.n14 ldomc_0.otaldom_0.pcascodeupm_0.o2.t15 13.847
R90936 ldomc_0.otaldom_0.pcascodeupm_0.o2.n20 ldomc_0.otaldom_0.pcascodeupm_0.o2.t8 13.847
R90937 ldomc_0.otaldom_0.pcascodeupm_0.o2.n20 ldomc_0.otaldom_0.pcascodeupm_0.o2.t13 13.847
R90938 ldomc_0.otaldom_0.pcascodeupm_0.o2.n16 ldomc_0.otaldom_0.pcascodeupm_0.o2.t10 13.847
R90939 ldomc_0.otaldom_0.pcascodeupm_0.o2.n16 ldomc_0.otaldom_0.pcascodeupm_0.o2.t11 13.847
R90940 ldomc_0.otaldom_0.pcascodeupm_0.o2.n12 ldomc_0.otaldom_0.pcascodeupm_0.o2.t0 13.847
R90941 ldomc_0.otaldom_0.pcascodeupm_0.o2.n12 ldomc_0.otaldom_0.pcascodeupm_0.o2.t7 13.847
R90942 ldomc_0.otaldom_0.pcascodeupm_0.o2.n3 ldomc_0.otaldom_0.pcascodeupm_0.o2.n7 6.881
R90943 ldomc_0.otaldom_0.pcascodeupm_0.o2.n22 ldomc_0.otaldom_0.pcascodeupm_0.o2.n20 6.852
R90944 ldomc_0.otaldom_0.pcascodeupm_0.o2.n2 ldomc_0.otaldom_0.pcascodeupm_0.o2.n9 5.97
R90945 ldomc_0.otaldom_0.pcascodeupm_0.o2.n13 ldomc_0.otaldom_0.pcascodeupm_0.o2.n12 5.76
R90946 ldomc_0.otaldom_0.pcascodeupm_0.o2.n0 ldomc_0.otaldom_0.pcascodeupm_0.o2.n19 5.681
R90947 ldomc_0.otaldom_0.pcascodeupm_0.o2.n26 ldomc_0.otaldom_0.pcascodeupm_0.o2.n25 5.621
R90948 ldomc_0.otaldom_0.pcascodeupm_0.o2.n17 ldomc_0.otaldom_0.pcascodeupm_0.o2.n16 5.536
R90949 ldomc_0.otaldom_0.pcascodeupm_0.o2.n22 ldomc_0.otaldom_0.pcascodeupm_0.o2.n21 4.5
R90950 ldomc_0.otaldom_0.pcascodeupm_0.o2.n8 ldomc_0.otaldom_0.pcascodeupm_0.o2.n27 4.5
R90951 ldomc_0.otaldom_0.pcascodeupm_0.o2.n3 ldomc_0.otaldom_0.pcascodeupm_0.o2.n29 4.5
R90952 ldomc_0.otaldom_0.pcascodeupm_0.o2.n23 ldomc_0.otaldom_0.pcascodeupm_0.o2 3.322
R90953 ldomc_0.otaldom_0.pcascodeupm_0.o2.n4 ldomc_0.otaldom_0.pcascodeupm_0.o2.n11 3.03
R90954 ldomc_0.otaldom_0.pcascodeupm_0.o2.n5 ldomc_0.otaldom_0.pcascodeupm_0.o2.n18 3.029
R90955 ldomc_0.otaldom_0.pcascodeupm_0.o2.n3 ldomc_0.otaldom_0.pcascodeupm_0.o2.n28 2.181
R90956 ldomc_0.otaldom_0.pcascodeupm_0.o2.n1 ldomc_0.otaldom_0.pcascodeupm_0.o2.n23 2.04
R90957 ldomc_0.otaldom_0.pcascodeupm_0.o2.n30 ldomc_0.otaldom_0.pcascodeupm_0.o2.n1 2.039
R90958 ldomc_0.otaldom_0.pcascodeupm_0.o2 ldomc_0.otaldom_0.pcascodeupm_0.o2.n6 1.557
R90959 ldomc_0.otaldom_0.pcascodeupm_0.o2.n15 ldomc_0.otaldom_0.pcascodeupm_0.o2.n6 3.983
R90960 ldomc_0.otaldom_0.pcascodeupm_0.o2.n5 ldomc_0.otaldom_0.pcascodeupm_0.o2.n17 1.309
R90961 ldomc_0.otaldom_0.pmosrm_0.o2 ldomc_0.otaldom_0.pcascodeupm_0.o2.n30 1.243
R90962 ldomc_0.otaldom_0.pcascodeupm_0.o2.n8 ldomc_0.otaldom_0.pcascodeupm_0.o2.n26 1.033
R90963 ldomc_0.otaldom_0.pcascodeupm_0.o2.n4 ldomc_0.otaldom_0.pcascodeupm_0.o2.n13 0.999
R90964 ldomc_0.otaldom_0.pmosrm_0.o2 ldomc_0.otaldom_0.pcascodeupm_0.o2.n2 0.882
R90965 ldomc_0.otaldom_0.pcascodeupm_0.o2.n0 ldomc_0.otaldom_0.pcascodeupm_0.o2.n22 0.756
R90966 ldomc_0.otaldom_0.pcascodeupm_0.o2.n8 ldomc_0.otaldom_0.pcascodeupm_0.o2.n24 0.613
R90967 ldomc_0.otaldom_0.pcascodeupm_0.o2.n6 ldomc_0.otaldom_0.pcascodeupm_0.o2.n14 9.628
R90968 ldomc_0.otaldom_0.pcascodeupm_0.o2.n30 ldomc_0.otaldom_0.pcascodeupm_0.o2.n3 1.216
R90969 ldomc_0.otaldom_0.pcascodeupm_0.o2.n19 ldomc_0.otaldom_0.pcascodeupm_0.o2.n5 0.923
R90970 ldomc_0.otaldom_0.pcascodeupm_0.o2.n1 ldomc_0.otaldom_0.pcascodeupm_0.o2.n8 0.865
R90971 ldomc_0.otaldom_0.pcascodeupm_0.o2.n2 ldomc_0.otaldom_0.pcascodeupm_0.o2.n4 0.862
R90972 ldomc_0.otaldom_0.pcascodeupm_0.o2.n23 ldomc_0.otaldom_0.pcascodeupm_0.o2.n0 0.805
R90973 ldomc_0.otaldom_0.pcascodeupm_0.o2.n4 ldomc_0.otaldom_0.pcascodeupm_0.o2.n10 0.626
R90974 trim[0] trim[0].t0 125.051
R90975 bandgapmd_0.trim[0] trim[0] 0.087
R90976 bandgapmd_0.trim[0] trim[0] 0.037
R90977 trim[1] trim[1].t0 125.208
R90978 trim[1] bandgapmd_0.trim[1] 0.045
R90979 trim[11] trim[11].t0 125.202
R90980 bandgapmd_0.trim[11] trim[11] 0.073
R90981 bandgapmd_0.trim[11] trim[11] 0.003
R90982 trim[2] trim[2].t0 125.035
R90983 bandgapmd_0.trim[2] trim[2] 0.16
R90984 bandgapmd_0.trim[2] trim[2] 0.01
R90985 trim[4] trim[4].t0 125.067
R90986 bandgapmd_0.trim[4] trim[4] 0.097
R90987 bandgapmd_0.trim[4] trim[4] 0.039
R90988 bandgapmd_0.trim[14] trim[14].t0 125.017
R90989 bandgapmd_0.trim[14] trim[14] 0.03
R90990 bandgapmd_0.trim[5] trim[5].t0 125.171
R90991 bandgapmd_0.trim[5] trim[5] 0.027
R90992 trim[10] trim[10].t0 125.088
R90993 bandgapmd_0.trim[10] trim[10] 0.096
R90994 bandgapmd_0.trim[10] trim[10] 0.026
R90995 trim[9] trim[9].t0 125.169
R90996 bandgapmd_0.trim[9] trim[9] 0.057
R90997 bandgapmd_0.trim[9] trim[9] 0.012
R90998 trim[15] trim[15].t0 125.107
R90999 bandgapmd_0.trim[15] trim[15] 0.065
R91000 bandgapmd_0.trim[15] trim[15] 0.002
R91001 trim[13] trim[13].t0 125.162
R91002 bandgapmd_0.trim[13] trim[13] 0.067
R91003 bandgapmd_0.trim[13] trim[13] 0.015
R91004 trim[6] trim[6].t0 125.065
R91005 bandgapmd_0.trim[6] trim[6] 0.121
R91006 trim[6].n0 trim[6] 0.028
R91007 trim[6].n0 trim[6] 0.027
R91008 bandgapmd_0.trim[6] trim[6].n0 0.006
R91009 bandgapmd_0.trim[3] trim[3].t0 125.202
R91010 bandgapmd_0.trim[3] trim[3] 0.003
R91011 trim[8] trim[8].t0 125.094
R91012 trim[7] trim[7].t0 125.199
R91013 bandgapmd_0.trim[7] trim[7] 0.043
R91014 bandgapmd_0.trim[7] trim[7] 0.009
R91015 bandgapmd_0.trim[12] trim[12].t0 125.056
R91016 trim[12].n0 trim[12] 0.095
R91017 trim[12] bandgapmd_0.trim[12] 0.012
R91018 bandgapmd_0.trim[12] trim[12] 0.011
R91019 trim[12].n0 trim[12] 0.003
R91020 trim[12] trim[12].n0 0.002
C0 a_8764_8048# ldomc_0.otaldom_0.pcsm_0.vbp1 0.00fF
C1 bandgapmd_0.otam_1.pdiffm_0.inn a_n17534_4148# 0.01fF
C2 a_n17534_4148# bandgapmd_0.bg_resm_0.trimup 0.05fF
C3 a_n11912_5108# bandgapmd_0.bg_pmosm_0.comp 0.00fF
C4 a_n11678_5108# bandgapmd_0.bg_pmosm_0.vbg 0.00fF
C5 a_n18594_4148# a_n17534_4148# 0.16fF
C6 vdd ldomc_0.otaldom_0.nmoslm_0.outp 1.51fF
C7 vdd ldomc_0.otaldom_0.pcsm_0.vbn2 8.11fF
C8 vdd bandgapmd_0.otam_1.pmosrm_0.bias1 217.11fF
C9 trim[6] a_n21356_2676# 0.00fF
C10 a_n19218_2674# trim[9] 0.00fF
C11 trim[0] trim[4] 0.00fF
C12 bandgapmd_0.otam_1.pdiffm_0.inp a_n17534_4148# 0.00fF
C13 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pcascodeupm_0.o2 6.82fF
C14 vdd ldomc_0.otaldom_0.pcsm_0.diff 29.15fF
C15 a_n22428_2672# trim[5] 0.11fF
C16 a_n15188_2076# a_n14486_2076# 0.00fF
C17 ldomc_0.otaldom_0.pcsm_0.vbp1 bandgapmd_0.bg_pmosm_0.vbg 0.06fF
C18 bandgapmd_0.bg_trimmup_0.bot trim[4] 0.43fF
C19 a_n23894_4148# a_n24544_2674# 0.03fF
C20 a_n22834_4148# a_n21774_4148# 0.16fF
C21 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.nmosbn1m_0.vbn1 0.00fF
C22 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 a_n14954_5108# 0.00fF
C23 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pcascodeupm_0.o1 0.52fF
C24 bandgapmd_0.otam_1.pdiffm_0.inn trim[8] 0.04fF
C25 a_n20714_4148# trim[12] 0.00fF
C26 trim[10] a_n19654_4148# 0.06fF
C27 ldomc_0.otaldom_0.pmosrm_0.bias1 bandgapmd_0.bg_pmosm_0.vbg 0.70fF
C28 ldomc_0.otaldom_0.pdiffm_0.inp biasldo 0.01fF
C29 a_n14954_5108# a_n12614_5108# 0.00fF
C30 a_n14720_5108# a_n12848_5108# 0.00fF
C31 a_8644_10248# a_8884_10248# 0.63fF
C32 vdd bandgapmd_0.bg_trimmup_0.bot 1.30fF
C33 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.nmosrm_0.outn 5.58fF
C34 a_n11678_5108# bandgapmd_0.bg_pmosm_0.comp 0.00fF
C35 a_n11444_2076# a_n11210_2076# 1.03fF
C36 out a_8404_8048# 0.65fF
C37 out ldomc_0.otaldom_0.pcsm_0.vbn2 0.00fF
C38 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pcascodeupm_0.vg 0.77fF
C39 bandgapmd_0.otam_1.pdiffm_0.inp trim[8] 0.00fF
C40 trim[7] trim[11] 0.00fF
C41 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 0.19fF
C42 trim[12] a_n19218_2674# 0.00fF
C43 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcascodeupm_0.o1 0.00fF
C44 vdd ldomc_0.otaldom_0.pcsm_0.vbp1 19.21fF
C45 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.nmoslm_0.outp 0.00fF
C46 bandgapmd_0.bg_resm_0.trimup a_n13550_2076# 0.72fF
C47 out ldomc_0.otaldom_0.pcsm_0.diff 0.00fF
C48 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pcsm_0.vbn2 5.09fF
C49 a_n7846_4436# bandgapmd_0.bg_stupm_0.vs2 0.52fF
C50 a_n21774_4148# a_n21356_2676# 0.05fF
C51 a_n19218_2674# trim[11] 0.11fF
C52 trim[2] a_n23894_4148# 0.08fF
C53 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.nmosrm_0.outn 0.58fF
C54 a_n17534_4148# trim[15] 0.00fF
C55 vdd ldomc_0.otaldom_0.pmosrm_0.bias1 216.63fF
C56 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcascodeupm_0.vg 0.00fF
C57 trim[6] trim[8] 0.03fF
C58 a_n22428_2672# trim[7] 0.02fF
C59 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 a_n14720_5108# 0.00fF
C60 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.nmoslm_0.outp 2.69fF
C61 bandgapmd_0.bg_trimmup_0.bot a_n22834_4148# 0.23fF
C62 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcsm_0.vbn2 2.09fF
C63 ldomc_0.otaldom_0.pdiffm_0.inp a_8404_8048# 0.90fF
C64 bandgapmd_0.otam_1.pdiffm_0.inn a_n14954_5108# 0.01fF
C65 bandgapmd_0.bg_trimmup_0.bot trim[14] 0.44fF
C66 a_n21356_2676# a_n20290_2674# 0.16fF
C67 bandgapmd_0.otam_1.pdiffm_0.inn a_n20714_4148# 0.01fF
C68 out a_8524_8048# 0.03fF
C69 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 a_n12848_5108# 0.00fF
C70 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcsm_0.diff 4.96fF
C71 out ldomc_0.otaldom_0.pcsm_0.vbp1 0.00fF
C72 bandgapmd_0.otam_1.pdiffm_0.inp a_n14954_5108# 0.83fF
C73 a_n12848_5108# a_n12614_5108# 0.98fF
C74 bandgapmd_0.bg_resm_0.trimup a_n13316_2076# 1.16fF
C75 trim[9] trim[11] 0.04fF
C76 a_n19218_2674# bandgapmd_0.bg_resm_0.trimup 0.00fF
C77 a_n18594_4148# a_n19218_2674# 0.03fF
C78 a_n14954_5108# a_n14018_5108# 0.43fF
C79 bandgapmd_0.bg_trimmup_0.bot a_n21356_2676# 0.23fF
C80 trim[4] a_n23460_2674# 0.00fF
C81 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 biasbgr 0.54fF
C82 a_n19218_2674# trim[13] 0.02fF
C83 bandgapmd_0.bg_resm_0.trimup a_n11444_2076# 0.00fF
C84 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pmosrm_0.bias1 10.06fF
C85 bandgapmd_0.bg_trimmup_0.bot trim[3] 0.39fF
C86 bandgapmd_0.otam_1.pdiffm_0.inn trim[2] 0.05fF
C87 ldomc_0.otaldom_0.pdiffm_0.inp a_8524_8048# 0.83fF
C88 trim[6] a_n20714_4148# 0.00fF
C89 a_n21774_4148# trim[8] 0.00fF
C90 a_n22428_2672# trim[9] 0.00fF
C91 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pcsm_0.vbp1 0.55fF
C92 bandgapmd_0.otam_1.pdiffm_0.inn a_n14720_5108# 0.00fF
C93 trim[10] trim[14] 0.00fF
C94 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 a_n12614_5108# 0.00fF
C95 bandgapmd_0.otam_1.pdiffm_0.inp trim[2] 0.00fF
C96 bandgapmd_0.bg_trimmup_0.bot a_n17534_4148# 0.23fF
C97 ldomc_0.otaldom_0.pdiffm_0.inp ldomc_0.otaldom_0.pmosrm_0.bias1 1.33fF
C98 bandgapmd_0.otam_1.pdiffm_0.inp a_n14720_5108# 0.03fF
C99 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.otam_1.nmosbn1m_0.vbn1 0.02fF
C100 bandgapmd_0.otam_1.nmosrm_0.outn biasbgr 0.00fF
C101 trim[8] a_n20290_2674# 0.00fF
C102 a_n15422_2076# a_n13550_2076# 0.00fF
C103 a_n14720_5108# a_n14018_5108# 0.00fF
C104 bandgapmd_0.otam_1.nmoslm_0.outp biasbgr 0.00fF
C105 trim[9] trim[13] 0.00fF
C106 bandgapmd_0.otam_1.nmosrm_0.outn bandgapmd_0.otam_1.nmosbn1m_0.vbn1 6.45fF
C107 bandgapmd_0.otam_1.pdiffm_0.inp a_n12848_5108# 0.77fF
C108 trim[2] trim[6] 0.00fF
C109 vdd bandgapmd_0.bg_pmosm_0.vbg 22.00fF
C110 a_n22834_4148# a_n23460_2674# 0.03fF
C111 bandgapmd_0.otam_1.pdiffm_0.inn biasbgr 1.22fF
C112 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 9.34fF
C113 bandgapmd_0.otam_1.nmosrm_0.outn bandgapmd_0.otam_1.pmosrm_0.out 6.60fF
C114 a_n19218_2674# trim[15] 0.00fF
C115 a_n14018_5108# a_n12848_5108# 0.06fF
C116 vdd a_n14486_2076# 0.01fF
C117 bandgapmd_0.bg_trimmup_0.bot trim[8] 0.39fF
C118 bandgapmd_0.otam_1.pdiffm_0.inn a_n23894_4148# 0.01fF
C119 bandgapmd_0.bg_pmosm_0.vbg bandgapmd_0.bg_pmosm_0.comp 2.83fF
C120 bandgapmd_0.bg_trimmup_0.bot trim[5] 0.38fF
C121 out a_8764_8048# 0.02fF
C122 a_n21774_4148# a_n20714_4148# 0.16fF
C123 a_n21774_4148# trim[7] 0.00fF
C124 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.nmosbn1m_0.vbn1 1.15fF
C125 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.pmosrm_0.out 0.01fF
C126 bandgapmd_0.otam_1.pdiffm_0.inp biasbgr 1.07fF
C127 bandgapmd_0.otam_1.pdiffm_0.inn trim[12] 0.04fF
C128 trim[12] a_n18594_4148# 0.13fF
C129 trim[14] a_n18160_2676# 0.00fF
C130 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.otam_1.nmosbn1m_0.vbn1 0.75fF
C131 bandgapmd_0.otam_1.nmoslm_0.outp bandgapmd_0.otam_1.nmosrm_0.outn 14.13fF
C132 a_n14486_2076# a_n14252_2076# 0.94fF
C133 a_n15188_2076# a_n13550_2076# 0.00fF
C134 bandgapmd_0.otam_1.pdiffm_0.inp trim[12] 0.00fF
C135 a_n20714_4148# a_n20290_2674# 0.05fF
C136 bandgapmd_0.otam_1.pdiffm_0.inp a_n12614_5108# 0.04fF
C137 a_n20290_2674# trim[7] 0.00fF
C138 vdd bandgapmd_0.bg_pmosm_0.comp 2.16fF
C139 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 a_n14018_5108# 0.00fF
C140 trim[11] trim[13] 0.04fF
C141 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.otam_1.pmosrm_0.out 0.00fF
C142 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.nmosrm_0.outn 2.48fF
C143 ldomc_0.otaldom_0.pdiffm_0.inp a_8764_8048# 0.73fF
C144 trim[0] a_n24544_2674# 0.00fF
C145 trim[4] a_n22834_4148# 0.06fF
C146 a_n23894_4148# trim[6] 0.00fF
C147 a_n13784_5108# a_n12848_5108# 0.00fF
C148 a_n14486_2076# a_n12380_2076# 0.00fF
C149 a_n14018_5108# a_n12614_5108# 0.00fF
C150 a_n23460_2674# trim[3] 0.11fF
C151 a_n20290_2674# a_n19218_2674# 0.16fF
C152 trim[8] trim[10] 0.04fF
C153 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.pmosrm_0.out 5.79fF
C154 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.otam_1.nmosrm_0.outn 0.43fF
C155 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.otam_1.nmoslm_0.outp 0.49fF
C156 bandgapmd_0.bg_trimmup_0.bot a_n24544_2674# 0.41fF
C157 bandgapmd_0.bg_trimmup_0.bot a_n20714_4148# 0.23fF
C158 bandgapmd_0.bg_trimmup_0.bot trim[7] 0.50fF
C159 a_n12848_5108# a_n11912_5108# 0.48fF
C160 vdd out 518.05fF
C161 vdd a_n12380_2076# 0.04fF
C162 bandgapmd_0.otam_1.pcsm_0.vbn2 biasbgr 0.17fF
C163 bandgapmd_0.otam_1.pcascodeupm_0.o2 bandgapmd_0.otam_1.nmosrm_0.outn 0.09fF
C164 bandgapmd_0.otam_1.pcascodeupm_0.o1 bandgapmd_0.otam_1.pmosrm_0.out 0.00fF
C165 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.nmosbn1m_0.vbn1 0.05fF
C166 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.otam_1.nmoslm_0.outp 2.51fF
C167 ldomc_0.otaldom_0.pdiffm_0.inp bandgapmd_0.bg_pmosm_0.vbg 6.16fF
C168 bandgapmd_0.otam_1.pdiffm_0.inn a_n18594_4148# 0.01fF
C169 bandgapmd_0.bg_trimmup_0.bot a_n19218_2674# 0.23fF
C170 vdd ldomc_0.otaldom_0.pmosrm_0.out 128.12fF
C171 a_n17534_4148# a_n18160_2676# 0.03fF
C172 bandgapmd_0.bg_resm_0.trimup trim[13] 0.00fF
C173 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.otam_1.pdiffm_0.inn 16.34fF
C174 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 7.06fF
C175 bandgapmd_0.otam_1.pcascodeupm_0.o1 bandgapmd_0.otam_1.nmosrm_0.outn 0.17fF
C176 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pmosrm_0.out 0.17fF
C177 trim[0] trim[2] 0.04fF
C178 a_n18594_4148# trim[13] 0.00fF
C179 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 a_n13784_5108# 0.00fF
C180 bandgapmd_0.otam_1.pmosrm_0.out a_n7846_4436# 0.06fF
C181 a_8164_10248# a_9124_10248# 0.01fF
C182 trim[6] a_n22428_2672# 0.00fF
C183 a_n20290_2674# trim[9] 0.11fF
C184 a_n14252_2076# a_n12380_2076# 0.00fF
C185 a_n14486_2076# a_n12146_2076# 0.00fF
C186 a_n13784_5108# a_n12614_5108# 0.00fF
C187 bandgapmd_0.otam_1.pdiffm_0.inn a_n14018_5108# 0.00fF
C188 trim[11] trim[15] 0.00fF
C189 bandgapmd_0.otam_1.pcascodeupm_0.o1 bandgapmd_0.otam_1.nmoslm_0.outp 0.01fF
C190 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pmosrm_0.out 6.46fF
C191 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.nmosrm_0.outn 2.77fF
C192 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.nmosbn1m_0.vbn1 0.08fF
C193 out a_8164_10248# 0.00fF
C194 bandgapmd_0.bg_trimmup_0.bot trim[2] 0.37fF
C195 bandgapmd_0.bg_pmosm_0.vbg bandgapmd_0.bg_stupm_0.vs2 2.30fF
C196 out a_9124_10248# 0.03fF
C197 a_n24956_4148# a_n24544_2674# 0.05fF
C198 vdd ldomc_0.otaldom_0.pdiffm_0.inp 11.32fF
C199 a_n23460_2674# trim[5] 0.02fF
C200 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 a_n11912_5108# 0.00fF
C201 bandgapmd_0.otam_1.pdiffm_0.inn trim[6] 0.04fF
C202 bandgapmd_0.otam_1.pdiffm_0.inp a_n14018_5108# 0.78fF
C203 trim[8] a_n19654_4148# 0.00fF
C204 a_n20714_4148# trim[10] 0.00fF
C205 a_n12614_5108# a_n11912_5108# 0.00fF
C206 bandgapmd_0.otam_1.pmosrm_0.bias1 biasbgr 2.71fF
C207 bandgapmd_0.otam_1.pcascodeupm_0.o1 bandgapmd_0.otam_1.pdiffm_0.inn 0.00fF
C208 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.nmoslm_0.outp 6.36fF
C209 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmosrm_0.outn 9.97fF
C210 vdd trim[3] 0.01fF
C211 vdd a_n12146_2076# 0.01fF
C212 bandgapmd_0.otam_1.pmosrm_0.out a_n11912_5108# 0.01fF
C213 bandgapmd_0.bg_trimmup_0.bot trim[9] 0.39fF
C214 a_8164_10248# a_8284_10248# 1.40fF
C215 ldomc_0.otaldom_0.pmosrm_0.out out 171.71fF
C216 bandgapmd_0.otam_1.pdiffm_0.inp trim[6] 0.00fF
C217 a_8284_10248# a_9124_10248# 0.00fF
C218 bandgapmd_0.otam_1.pcascodeupm_0.o1 bandgapmd_0.otam_1.pdiffm_0.inp 0.00fF
C219 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.nmoslm_0.outp 21.57fF
C220 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pdiffm_0.inn 0.00fF
C221 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 0.87fF
C222 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.nmosrm_0.outn 8.18fF
C223 trim[10] a_n19218_2674# 0.00fF
C224 vdd bandgapmd_0.bg_stupm_0.vs2 3.51fF
C225 a_8164_10248# ldomc_0.otaldom_0.pdiffm_0.inp 0.04fF
C226 ldomc_0.otaldom_0.pdiffm_0.inp a_9124_10248# 0.00fF
C227 bandgapmd_0.bg_resm_0.trimup trim[15] 0.26fF
C228 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.nmoslm_0.outp 8.49fF
C229 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pmosrm_0.out 9.39fF
C230 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.nmosrm_0.outn 0.00fF
C231 bandgapmd_0.otam_1.pcascodeupm_0.o1 bandgapmd_0.otam_1.pcascodeupm_0.o2 7.04fF
C232 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pdiffm_0.inp 0.00fF
C233 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pdiffm_0.inn 0.87fF
C234 trim[0] a_n23894_4148# 0.00fF
C235 a_9124_10248# a_9244_10248# 1.40fF
C236 out ldomc_0.otaldom_0.pdiffm_0.inp 109.34fF
C237 a_n21774_4148# a_n22428_2672# 0.03fF
C238 out a_9244_10248# 0.02fF
C239 trim[4] trim[8] 0.00fF
C240 a_n20290_2674# trim[11] 0.02fF
C241 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 a_n11678_5108# 0.00fF
C242 trim[13] trim[15] 0.04fF
C243 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pdiffm_0.inp 1.89fF
C244 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o2 5.07fF
C245 bandgapmd_0.bg_trimmup_0.bot a_n23894_4148# 0.19fF
C246 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inn 6.12fF
C247 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.nmoslm_0.outp 0.00fF
C248 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.nmosrm_0.outn 2.36fF
C249 bandgapmd_0.otam_1.pdiffm_0.inp a_n13784_5108# 0.04fF
C250 a_n24544_2674# a_n23460_2674# 0.16fF
C251 a_n12380_2076# a_n12146_2076# 0.92fF
C252 ldomc_0.otaldom_0.pmosrm_0.out ldomc_0.otaldom_0.pdiffm_0.inp 0.02fF
C253 a_n23460_2674# trim[7] 0.00fF
C254 bandgapmd_0.bg_trimmup_0.bot trim[12] 0.39fF
C255 bandgapmd_0.otam_1.pdiffm_0.inn a_n21774_4148# 0.01fF
C256 bandgapmd_0.otam_1.pmosrm_0.out a_n11678_5108# 0.01fF
C257 ldomc_0.otaldom_0.pdiffm_0.inp a_8284_10248# 0.02fF
C258 a_n20714_4148# a_n19654_4148# 0.16fF
C259 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pdiffm_0.inp 5.02fF
C260 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.nmoslm_0.outp 0.46fF
C261 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pdiffm_0.inn 0.04fF
C262 vdd trim[5] 0.01fF
C263 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcascodeupm_0.o2 0.01fF
C264 bandgapmd_0.otam_1.pcascodeupm_0.vg bandgapmd_0.otam_1.pcascodeupm_0.o1 20.42fF
C265 a_n14018_5108# a_n13784_5108# 1.06fF
C266 a_n14486_2076# a_n13550_2076# 0.39fF
C267 bandgapmd_0.bg_resm_0.trimup a_n15422_2076# 0.89fF
C268 bandgapmd_0.bg_trimmup_0.bot trim[11] 0.39fF
C269 bandgapmd_0.otam_1.pdiffm_0.inp a_n11912_5108# 0.32fF
C270 trim[14] a_n17534_4148# 0.06fF
C271 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcascodeupm_0.o1 0.01fF
C272 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcascodeupm_0.o2 0.00fF
C273 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pdiffm_0.inp 0.04fF
C274 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pdiffm_0.inn 0.65fF
C275 a_n19654_4148# a_n19218_2674# 0.05fF
C276 a_n14018_5108# a_n11912_5108# 0.00fF
C277 vdd a_n13550_2076# 0.05fF
C278 a_n19218_2674# a_n18160_2676# 0.16fF
C279 trim[2] a_n23460_2674# 0.00fF
C280 bandgapmd_0.otam_1.pcsm_0.vbn2 bandgapmd_0.otam_1.pcascodeupm_0.vg 4.91fF
C281 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pdiffm_0.inp 0.93fF
C282 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcascodeupm_0.o1 0.00fF
C283 a_n24956_4148# a_n23894_4148# 0.16fF
C284 bandgapmd_0.bg_trimmup_0.bot a_n22428_2672# 0.23fF
C285 bandgapmd_0.otam_1.pdiffm_0.inn trim[0] 0.04fF
C286 a_n22834_4148# trim[8] 0.00fF
C287 a_n20290_2674# trim[13] 0.00fF
C288 trim[6] a_n21774_4148# 0.06fF
C289 a_n22834_4148# trim[5] 0.00fF
C290 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o2 7.05fF
C291 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcascodeupm_0.vg 0.06fF
C292 trim[10] trim[12] 0.04fF
C293 a_n14252_2076# a_n13550_2076# 0.00fF
C294 a_n14486_2076# a_n13316_2076# 0.00fF
C295 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 biasldo 0.54fF
C296 bandgapmd_0.otam_1.pdiffm_0.inp trim[0] 0.00fF
C297 bandgapmd_0.otam_1.pdiffm_0.inn bandgapmd_0.bg_trimmup_0.bot 8.48fF
C298 bandgapmd_0.bg_trimmup_0.bot bandgapmd_0.bg_resm_0.trimup 0.86fF
C299 bandgapmd_0.bg_resm_0.trimup a_n15188_2076# 0.05fF
C300 bandgapmd_0.bg_trimmup_0.bot a_n18594_4148# 0.23fF
C301 bandgapmd_0.otam_1.pdiffm_0.inp a_n11678_5108# 0.02fF
C302 ldomc_0.otaldom_0.pcascodeupm_0.o1 ldomc_0.otaldom_0.pcascodeupm_0.o2 7.04fF
C303 vdd trim[7] 0.01fF
C304 bandgapmd_0.otam_1.pcsm_0.diff bandgapmd_0.otam_1.pcsm_0.vbn2 4.85fF
C305 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.o1 7.12fF
C306 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcascodeupm_0.vg 0.00fF
C307 bandgapmd_0.bg_trimmup_0.bot trim[13] 0.44fF
C308 ldomc_0.otaldom_0.nmosrm_0.outn biasldo 0.00fF
C309 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.bg_trimmup_0.bot 0.07fF
C310 a_n14018_5108# a_n11678_5108# 0.00fF
C311 a_n13784_5108# a_n11912_5108# 0.00fF
C312 ldomc_0.otaldom_0.pcascodeupm_0.o2 ldomc_0.otaldom_0.nmosrm_0.outn 0.09fF
C313 a_n13550_2076# a_n12380_2076# 0.38fF
C314 vdd a_n13316_2076# 0.01fF
C315 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o2 5.07fF
C316 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcascodeupm_0.vg 12.28fF
C317 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.vbn2 5.30fF
C318 trim[8] a_n21356_2676# 0.00fF
C319 trim[2] trim[4] 0.04fF
C320 a_n21356_2676# trim[5] 0.00fF
C321 ldomc_0.otaldom_0.nmoslm_0.outp biasldo 0.00fF
C322 ldomc_0.otaldom_0.nmosrm_0.outn ldomc_0.otaldom_0.nmosbn1m_0.vbn1 6.45fF
C323 ldomc_0.otaldom_0.pcascodeupm_0.o1 ldomc_0.otaldom_0.nmosrm_0.outn 0.17fF
C324 ldomc_0.otaldom_0.pcsm_0.vbn2 biasldo 0.17fF
C325 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.nmosbn1m_0.vbn1 0.05fF
C326 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.pcascodeupm_0.o1 20.42fF
C327 a_n23894_4148# a_n23460_2674# 0.05fF
C328 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcascodeupm_0.o2 0.01fF
C329 a_n12848_5108# bandgapmd_0.bg_pmosm_0.vbg 0.00fF
C330 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcsm_0.vbn2 1.95fF
C331 bandgapmd_0.otam_1.pcsm_0.vbp1 bandgapmd_0.otam_1.pcsm_0.diff 5.32fF
C332 vdd a_n11444_2076# 0.04fF
C333 trim[3] trim[5] 0.03fF
C334 bandgapmd_0.bg_trimmup_0.bot trim[6] 0.44fF
C335 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosbn1m_0.vbn1 9.34fF
C336 bandgapmd_0.otam_1.pdiffm_0.inn a_n24956_4148# 0.01fF
C337 a_8164_10248# a_8644_10248# 0.63fF
C338 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.nmosrm_0.outn 2.77fF
C339 ldomc_0.otaldom_0.pcascodeupm_0.o1 ldomc_0.otaldom_0.nmoslm_0.outp 0.01fF
C340 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 7.12fF
C341 a_n14252_2076# a_n13316_2076# 0.00fF
C342 a_8644_10248# a_9124_10248# 0.00fF
C343 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcascodeupm_0.o1 0.01fF
C344 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcascodeupm_0.o2 0.00fF
C345 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcsm_0.diff 2.65fF
C346 bandgapmd_0.otam_1.pdiffm_0.inn trim[10] 0.05fF
C347 trim[10] a_n18594_4148# 0.00fF
C348 a_n19654_4148# trim[12] 0.00fF
C349 out a_8644_10248# 0.01fF
C350 ldomc_0.otaldom_0.nmoslm_0.outp ldomc_0.otaldom_0.nmosrm_0.outn 14.13fF
C351 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmosrm_0.outn 9.69fF
C352 ldomc_0.otaldom_0.pcascodeupm_0.vg ldomc_0.otaldom_0.nmoslm_0.outp 6.36fF
C353 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.nmosbn1m_0.vbn1 0.08fF
C354 trim[12] a_n18160_2676# 0.00fF
C355 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.pcascodeupm_0.vg 4.91fF
C356 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcascodeupm_0.o1 0.00fF
C357 a_n13316_2076# a_n12380_2076# 0.00fF
C358 a_n13550_2076# a_n12146_2076# 0.00fF
C359 vdd trim[9] 0.01fF
C360 bandgapmd_0.otam_1.pmosrm_0.bias1 bandgapmd_0.otam_1.pcsm_0.vbp1 4.29fF
C361 bandgapmd_0.otam_1.pdiffm_0.inp trim[10] 0.00fF
C362 a_n19654_4148# trim[11] 0.00fF
C363 bandgapmd_0.bg_trimmup_0.bot trim[15] 0.39fF
C364 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.nmosrm_0.outn 7.84fF
C365 a_n18160_2676# trim[11] 0.00fF
C366 ldomc_0.otaldom_0.pcsm_0.vbn2 ldomc_0.otaldom_0.nmoslm_0.outp 21.56fF
C367 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 bandgapmd_0.bg_pmosm_0.vbg 0.00fF
C368 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcascodeupm_0.vg 0.06fF
C369 a_n23460_2674# a_n22428_2672# 0.16fF
C370 a_n20714_4148# a_n21356_2676# 0.03fF
C371 a_n12614_5108# bandgapmd_0.bg_pmosm_0.vbg 0.00fF
C372 a_n11912_5108# a_n11678_5108# 0.94fF
C373 a_n12380_2076# a_n11444_2076# 0.45fF
C374 a_n12848_5108# bandgapmd_0.bg_pmosm_0.comp 0.00fF
C375 trim[2] a_n22834_4148# 0.00fF
C376 a_n21356_2676# trim[7] 0.03fF
C377 vdd a_n11210_2076# 0.01fF
C378 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.nmoslm_0.outp 8.19fF
C379 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.bg_pmosm_0.vbg 6.39fF
C380 a_8404_8048# ldomc_0.otaldom_0.pcsm_0.diff 0.01fF
C381 ldomc_0.otaldom_0.pdiffm_0.inp a_8644_10248# 0.01fF
C382 ldomc_0.otaldom_0.pcsm_0.diff ldomc_0.otaldom_0.pcsm_0.vbn2 4.72fF
C383 trim[6] trim[10] 0.00fF
C384 vdd biasbgr 0.02fF
C385 a_n24544_2674# trim[3] 0.02fF
C386 ldomc_0.otaldom_0.pmosrm_0.bias1 biasldo 2.73fF
C387 trim[3] trim[7] 0.00fF
C388 bandgapmd_0.bg_trimmup_0.bot a_n21774_4148# 0.23fF
C389 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o2 7.05fF
C390 a_n15422_2076# a_n15188_2076# 0.93fF
C391 vdd bandgapmd_0.otam_1.nmosbn1m_0.vbn1 0.37fF
C392 bandgapmd_0.otam_1.pdiffm_0.inn a_n19654_4148# 0.01fF
C393 a_n19654_4148# a_n18594_4148# 0.16fF
C394 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 0.88fF
C395 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.nmosrm_0.outn 0.00fF
C396 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcascodeupm_0.vg 0.00fF
C397 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.o1 7.12fF
C398 a_n18160_2676# bandgapmd_0.bg_resm_0.trimup 0.19fF
C399 a_n18594_4148# a_n18160_2676# 0.05fF
C400 vdd trim[11] 0.01fF
C401 vdd bandgapmd_0.otam_1.pmosrm_0.out 22.59fF
C402 a_8404_8048# a_8524_8048# 1.82fF
C403 bandgapmd_0.bg_trimmup_0.bot a_n20290_2674# 0.23fF
C404 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.nmosrm_0.outn 2.37fF
C405 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.nmoslm_0.outp 0.00fF
C406 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.vbn2 5.30fF
C407 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcascodeupm_0.vg 12.28fF
C408 a_8404_8048# ldomc_0.otaldom_0.pcsm_0.vbp1 0.00fF
C409 trim[4] a_n22428_2672# 0.00fF
C410 a_n12614_5108# bandgapmd_0.bg_pmosm_0.comp 0.00fF
C411 a_n18160_2676# trim[13] 0.03fF
C412 vdd bandgapmd_0.otam_1.nmosrm_0.outn 4.51fF
C413 bandgapmd_0.bg_trimmup_0.bot trim[0] 0.41fF
C414 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.bg_pmosm_0.comp 2.26fF
C415 a_8524_8048# ldomc_0.otaldom_0.pcsm_0.diff 0.00fF
C416 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.nmoslm_0.outp 0.45fF
C417 a_n23894_4148# a_n22834_4148# 0.16fF
C418 a_n21356_2676# trim[9] 0.02fF
C419 a_8884_10248# a_9124_10248# 0.61fF
C420 ldomc_0.otaldom_0.pcsm_0.vbp1 ldomc_0.otaldom_0.pcsm_0.diff 5.55fF
C421 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcsm_0.vbn2 2.01fF
C422 bandgapmd_0.bg_resm_0.trimup a_n14486_2076# 0.87fF
C423 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.bg_pmosm_0.vbg 0.05fF
C424 bandgapmd_0.otam_1.pdiffm_0.inn trim[4] 0.04fF
C425 a_n21774_4148# trim[10] 0.00fF
C426 trim[8] a_n20714_4148# 0.13fF
C427 out a_8884_10248# 0.01fF
C428 vdd bandgapmd_0.otam_1.nmoslm_0.outp 1.51fF
C429 trim[5] trim[7] 0.03fF
C430 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcsm_0.diff 2.31fF
C431 trim[12] trim[14] 0.03fF
C432 bandgapmd_0.otam_1.pdiffm_0.inp trim[4] 0.00fF
C433 vdd bandgapmd_0.otam_1.pdiffm_0.inn 8.77fF
C434 vdd bandgapmd_0.bg_resm_0.trimup 0.96fF
C435 a_8524_8048# ldomc_0.otaldom_0.pcsm_0.vbp1 0.00fF
C436 trim[10] a_n20290_2674# 0.00fF
C437 trim[0] a_n24956_4148# 0.06fF
C438 vdd bandgapmd_0.otam_1.pdiffm_0.inp 8.65fF
C439 vdd trim[13] 0.01fF
C440 ldomc_0.otaldom_0.pdiffm_0.inp a_8884_10248# 0.01fF
C441 a_n22834_4148# a_n22428_2672# 0.05fF
C442 a_n18160_2676# trim[15] 0.02fF
C443 trim[4] trim[6] 0.04fF
C444 a_n13550_2076# a_n13316_2076# 1.04fF
C445 a_n23894_4148# trim[3] 0.00fF
C446 bandgapmd_0.bg_resm_0.trimup a_n14252_2076# 0.06fF
C447 vdd bandgapmd_0.otam_1.pcascodeupm_0.o2 45.06fF
C448 ldomc_0.otaldom_0.pmosrm_0.bias1 ldomc_0.otaldom_0.pcsm_0.vbp1 4.27fF
C449 bandgapmd_0.bg_trimmup_0.bot a_n24956_4148# 0.27fF
C450 bandgapmd_0.otam_1.pdiffm_0.inp bandgapmd_0.bg_pmosm_0.comp 0.01fF
C451 bandgapmd_0.bg_pmosm_0.vbg a_n7846_4436# 1.34fF
C452 a_n21356_2676# trim[11] 0.00fF
C453 bandgapmd_0.bg_trimmup_0.bot trim[10] 0.45fF
C454 bandgapmd_0.otam_1.pdiffm_0.inn a_n22834_4148# 0.01fF
C455 vdd bandgapmd_0.otam_1.pcascodeupm_0.o1 30.60fF
C456 bandgapmd_0.bg_resm_0.trimup a_n12380_2076# 0.01fF
C457 trim[5] trim[9] 0.00fF
C458 bandgapmd_0.otam_1.pdiffm_0.inn trim[14] 0.03fF
C459 trim[14] bandgapmd_0.bg_resm_0.trimup 0.00fF
C460 bandgapmd_0.bg_pmosm_0.vbg ldomc_0.otaldom_0.nmosbn1m_0.vbn1 0.13fF
C461 trim[12] a_n17534_4148# 0.00fF
C462 ldomc_0.otaldom_0.pcascodeupm_0.o1 bandgapmd_0.bg_pmosm_0.vbg 0.00fF
C463 a_8404_8048# a_8764_8048# 0.00fF
C464 vdd bandgapmd_0.otam_1.pcascodeupm_0.vg 287.48fF
C465 a_n22428_2672# a_n21356_2676# 0.16fF
C466 a_n11912_5108# bandgapmd_0.bg_pmosm_0.vbg 0.45fF
C467 bandgapmd_0.otam_1.pdiffm_0.inp trim[14] 0.00fF
C468 vdd a_n7846_4436# 0.86fF
C469 bandgapmd_0.bg_pmosm_0.vbg ldomc_0.otaldom_0.nmosrm_0.outn 2.48fF
C470 ldomc_0.otaldom_0.pcascodeupm_0.vg bandgapmd_0.bg_pmosm_0.vbg 0.00fF
C471 bandgapmd_0.otam_1.pmosrm_0.out bandgapmd_0.bg_stupm_0.vs2 0.07fF
C472 vdd biasldo 0.00fF
C473 a_8764_8048# ldomc_0.otaldom_0.pcsm_0.diff 0.00fF
C474 a_n19654_4148# a_n20290_2674# 0.03fF
C475 vdd trim[15] 0.01fF
C476 vdd ldomc_0.otaldom_0.pcascodeupm_0.o2 45.06fF
C477 a_n22428_2672# trim[3] 0.00fF
C478 vdd bandgapmd_0.otam_1.pcsm_0.vbn2 8.12fF
C479 bandgapmd_0.bg_pmosm_0.comp a_n7846_4436# 0.00fF
C480 bandgapmd_0.bg_pmosm_0.vbg ldomc_0.otaldom_0.nmoslm_0.outp 0.49fF
C481 trim[2] a_n24544_2674# 0.00fF
C482 trim[4] a_n21774_4148# 0.00fF
C483 a_n22834_4148# trim[6] 0.00fF
C484 ldomc_0.otaldom_0.pcsm_0.vbn2 bandgapmd_0.bg_pmosm_0.vbg 0.89fF
C485 vdd ldomc_0.otaldom_0.nmosbn1m_0.vbn1 0.33fF
C486 a_n14954_5108# a_n14720_5108# 1.06fF
C487 a_n15422_2076# a_n14486_2076# 0.46fF
C488 bandgapmd_0.bg_trimmup_0.bot a_n23460_2674# 0.23fF
C489 vdd ldomc_0.otaldom_0.pcascodeupm_0.o1 30.59fF
C490 vdd bandgapmd_0.otam_1.pcsm_0.diff 26.49fF
C491 trim[8] trim[12] 0.00fF
C492 bandgapmd_0.bg_resm_0.trimup a_n12146_2076# 0.00fF
C493 bandgapmd_0.bg_trimmup_0.bot a_n19654_4148# 0.23fF
C494 ldomc_0.otaldom_0.pcsm_0.diff bandgapmd_0.bg_pmosm_0.vbg 4.91fF
C495 vdd ldomc_0.otaldom_0.nmosrm_0.outn 4.53fF
C496 vdd ldomc_0.otaldom_0.pcascodeupm_0.vg 286.90fF
C497 a_n14954_5108# a_n12848_5108# 0.00fF
C498 vdd bandgapmd_0.otam_1.pcsm_0.vbp1 19.77fF
C499 a_n20714_4148# trim[9] 0.00fF
C500 a_8524_8048# a_8764_8048# 0.19fF
C501 bandgapmd_0.bg_trimmup_0.bot a_n18160_2676# 0.23fF
C502 trim[7] trim[9] 0.03fF
C503 vdd a_n15422_2076# 0.01fF
C504 ldomc_0.otaldom_0.nmosbn1m_0.vbn1 vss -25.55fF
C505 ldomc_0.otaldom_0.nmosrm_0.outn vss 1.42fF
C506 ldomc_0.otaldom_0.nmoslm_0.outp vss -6.03fF
C507 bandgapmd_0.bg_stupm_0.vs2 vss 92.33fF
C508 a_n7846_4436# vss 1.08fF
C509 a_n11210_2076# vss 0.65fF
C510 a_n11444_2076# vss 1.22fF
C511 a_n11678_5108# vss 0.65fF
C512 a_n11912_5108# vss 0.67fF
C513 a_n12146_2076# vss 0.62fF
C514 a_n12380_2076# vss 0.80fF
C515 a_n12614_5108# vss 0.69fF
C516 a_n12848_5108# vss 0.80fF
C517 a_n13316_2076# vss 0.64fF
C518 a_n13550_2076# vss 0.82fF
C519 a_n13784_5108# vss 0.68fF
C520 a_n14018_5108# vss 0.83fF
C521 a_n14252_2076# vss 0.61fF
C522 a_n14486_2076# vss 0.67fF
C523 a_n14720_5108# vss 0.71fF
C524 a_n14954_5108# vss 0.76fF
C525 a_n15188_2076# vss 0.61fF
C526 a_n15422_2076# vss 1.11fF
C527 ldomc_0.otaldom_0.pcascodeupm_0.vg vss -78.53fF
C528 ldomc_0.otaldom_0.pcsm_0.vbn2 vss 325.71fF
C529 ldomc_0.otaldom_0.pcsm_0.diff vss -14.02fF
C530 bandgapmd_0.bg_resm_0.trimup vss 2.04fF
C531 a_n18160_2676# vss 1.04fF
C532 a_n19218_2674# vss 0.85fF
C533 a_n20290_2674# vss 0.88fF
C534 a_n21356_2676# vss 0.95fF
C535 a_n22428_2672# vss 0.88fF
C536 a_n23460_2674# vss 0.90fF
C537 a_n24544_2674# vss 0.88fF
C538 a_n17534_4148# vss 1.32fF
C539 a_n18594_4148# vss 0.99fF
C540 a_n19654_4148# vss 1.09fF
C541 a_n20714_4148# vss 1.03fF
C542 a_n21774_4148# vss 1.08fF
C543 a_n22834_4148# vss 1.12fF
C544 a_n23894_4148# vss 1.13fF
C545 a_n24956_4148# vss 1.30fF
C546 bandgapmd_0.bg_trimmup_0.bot vss 37.06fF
C547 ldomc_0.otaldom_0.pcsm_0.vbp1 vss -11.61fF
C548 ldomc_0.otaldom_0.pmosrm_0.bias1 vss -56.59fF
C549 a_9244_10248# vss 0.38fF
C550 a_9124_10248# vss 1.66fF
C551 a_8884_10248# vss 0.42fF
C552 a_8764_8048# vss 1.10fF
C553 a_8644_10248# vss 0.41fF
C554 a_8524_8048# vss 1.75fF
C555 a_8404_8048# vss 3.03fF
C556 a_8284_10248# vss 0.32fF
C557 ldomc_0.otaldom_0.pdiffm_0.inp vss 18.56fF
C558 a_8164_10248# vss 1.31fF
C559 bandgapmd_0.otam_1.nmosbn1m_0.vbn1 vss -25.66fF
C560 bandgapmd_0.otam_1.pmosrm_0.out vss 271.17fF
C561 bandgapmd_0.otam_1.nmoslm_0.outp vss -6.02fF
C562 bandgapmd_0.otam_1.pdiffm_0.inn vss -12.28fF
C563 bandgapmd_0.otam_1.pdiffm_0.inp vss 23.68fF
C564 bandgapmd_0.otam_1.pcascodeupm_0.o2 vss -12.22fF
C565 bandgapmd_0.otam_1.pcascodeupm_0.vg vss -78.54fF
C566 bandgapmd_0.otam_1.pcsm_0.vbn2 vss 326.02fF
C567 bandgapmd_0.otam_1.pcsm_0.diff vss -15.93fF
C568 bandgapmd_0.otam_1.pcsm_0.vbp1 vss -11.78fF
C569 bandgapmd_0.otam_1.pmosrm_0.bias1 vss -56.86fF
C570 ldomc_0.otaldom_0.pmosrm_0.out vss 13.66fF
C571 vdd vss -3677.03fF
C572 ldomc_0.otaldom_0.pcascodeupm_0.o2.t6 vss 0.18fF
C573 ldomc_0.otaldom_0.pcascodeupm_0.o2.t4 vss 0.18fF
C574 ldomc_0.otaldom_0.pcascodeupm_0.o2.t1 vss 0.18fF
C575 ldomc_0.otaldom_0.pcascodeupm_0.o2.t2 vss 0.18fF
C576 ldomc_0.otaldom_0.pcascodeupm_0.o2.t0 vss 0.18fF
C577 ldomc_0.otaldom_0.pcascodeupm_0.o2.t7 vss 0.18fF
C578 ldomc_0.otaldom_0.pcascodeupm_0.o2.t14 vss 0.18fF
C579 ldomc_0.otaldom_0.pcascodeupm_0.o2.t15 vss 0.18fF
C580 ldomc_0.otaldom_0.pcascodeupm_0.o2.t12 vss 0.18fF
C581 ldomc_0.otaldom_0.pcascodeupm_0.o2.t9 vss 0.18fF
C582 ldomc_0.otaldom_0.pcascodeupm_0.o2.t10 vss 0.18fF
C583 ldomc_0.otaldom_0.pcascodeupm_0.o2.t11 vss 0.18fF
C584 ldomc_0.otaldom_0.pcascodeupm_0.o2.t8 vss 0.18fF
C585 ldomc_0.otaldom_0.pcascodeupm_0.o2.t13 vss 0.18fF
C586 ldomc_0.otaldom_0.pcascodeupm_0.o2.t5 vss 0.18fF
C587 ldomc_0.otaldom_0.pcascodeupm_0.o2.t3 vss 0.18fF
C588 biasldo.t0 vss 20.49fF
C589 biasldo.t5 vss 20.49fF
C590 biasldo.t4 vss 20.49fF
C591 biasldo.t2 vss 20.49fF
C592 biasldo.t3 vss 0.21fF
C593 biasldo.t1 vss 0.21fF
C594 biasbgr.t0 vss 20.47fF
C595 biasbgr.t4 vss 20.47fF
C596 biasbgr.t5 vss 20.47fF
C597 biasbgr.t2 vss 20.47fF
C598 biasbgr.t3 vss 0.20fF
C599 biasbgr.t1 vss 0.20fF
C600 bandgapmd_0.bg_pmosm_0.comp.t2 vss 0.09fF
C601 bandgapmd_0.bg_pmosm_0.comp.t1 vss 0.09fF
C602 bandgapmd_0.bg_pmosm_0.comp.t0 vss 1.37fF
C603 bandgapmd_0.otam_1.pcascodeupm_0.o1.t5 vss 0.16fF
C604 bandgapmd_0.otam_1.pcascodeupm_0.o1.t1 vss 0.16fF
C605 bandgapmd_0.otam_1.pcascodeupm_0.o1.t0 vss 0.16fF
C606 bandgapmd_0.otam_1.pcascodeupm_0.o1.t3 vss 0.16fF
C607 bandgapmd_0.otam_1.pcascodeupm_0.o1.t13 vss 0.16fF
C608 bandgapmd_0.otam_1.pcascodeupm_0.o1.t8 vss 0.16fF
C609 bandgapmd_0.otam_1.pcascodeupm_0.o1.t15 vss 0.16fF
C610 bandgapmd_0.otam_1.pcascodeupm_0.o1.t12 vss 0.16fF
C611 bandgapmd_0.otam_1.pcascodeupm_0.o1.t14 vss 0.16fF
C612 bandgapmd_0.otam_1.pcascodeupm_0.o1.t10 vss 0.16fF
C613 bandgapmd_0.otam_1.pcascodeupm_0.o1.t9 vss 0.16fF
C614 bandgapmd_0.otam_1.pcascodeupm_0.o1.t11 vss 0.16fF
C615 bandgapmd_0.otam_1.pcascodeupm_0.o1.t4 vss 0.16fF
C616 bandgapmd_0.otam_1.pcascodeupm_0.o1.t7 vss 0.16fF
C617 bandgapmd_0.otam_1.pcascodeupm_0.o1.t6 vss 0.16fF
C618 bandgapmd_0.otam_1.pcascodeupm_0.o1.t2 vss 0.16fF
C619 bandgapmd_0.bg_pmosm_0.vbg.t0 vss 0.04fF
C620 bandgapmd_0.bg_pmosm_0.vbg.t1 vss 0.04fF
C621 bandgapmd_0.bg_pmosm_0.vbg.t5 vss 0.09fF
C622 bandgapmd_0.bg_pmosm_0.vbg.t7 vss 6.39fF
C623 bandgapmd_0.bg_pmosm_0.vbg.t8 vss 0.37fF
C624 bandgapmd_0.bg_pmosm_0.vbg.t6 vss 0.37fF
C625 bandgapmd_0.bg_pmosm_0.vbg.t10 vss 0.37fF
C626 bandgapmd_0.bg_pmosm_0.vbg.t14 vss 0.37fF
C627 bandgapmd_0.bg_pmosm_0.vbg.t11 vss 0.37fF
C628 bandgapmd_0.bg_pmosm_0.vbg.t4 vss 0.37fF
C629 bandgapmd_0.bg_pmosm_0.vbg.t3 vss 0.37fF
C630 bandgapmd_0.bg_pmosm_0.vbg.t12 vss 0.37fF
C631 bandgapmd_0.bg_pmosm_0.vbg.t13 vss 0.37fF
C632 bandgapmd_0.bg_pmosm_0.vbg.t9 vss 0.37fF
C633 bandgapmd_0.bg_pmosm_0.vbg.t2 vss 0.55fF
C634 bandgapmd_0.bg_stupm_0.vs2.t1 vss 3.72fF
C635 bandgapmd_0.bg_stupm_0.vs2.t0 vss 3.28fF
C636 bandgapmd_0.otam_1.pdiffm_0.inp.t10 vss 0.75fF
C637 bandgapmd_0.otam_1.pdiffm_0.inp.t8 vss 0.75fF
C638 bandgapmd_0.otam_1.pdiffm_0.inp.t4 vss 0.75fF
C639 bandgapmd_0.otam_1.pdiffm_0.inp.t2 vss 0.75fF
C640 bandgapmd_0.otam_1.pdiffm_0.inp.t6 vss 0.75fF
C641 bandgapmd_0.otam_1.pdiffm_0.inp.t5 vss 0.75fF
C642 bandgapmd_0.otam_1.pdiffm_0.inp.t9 vss 0.75fF
C643 bandgapmd_0.otam_1.pdiffm_0.inp.t7 vss 0.75fF
C644 bandgapmd_0.otam_1.pdiffm_0.inp.t3 vss 0.75fF
C645 bandgapmd_0.otam_1.pdiffm_0.inp.t11 vss 0.75fF
C646 bandgapmd_0.otam_1.pdiffm_0.inp.t0 vss 1.08fF
C647 ldomc_0.otaldom_0.pcascodeupm_0.o1.t4 vss 0.16fF
C648 ldomc_0.otaldom_0.pcascodeupm_0.o1.t1 vss 0.16fF
C649 ldomc_0.otaldom_0.pcascodeupm_0.o1.t5 vss 0.16fF
C650 ldomc_0.otaldom_0.pcascodeupm_0.o1.t3 vss 0.16fF
C651 ldomc_0.otaldom_0.pcascodeupm_0.o1.t11 vss 0.16fF
C652 ldomc_0.otaldom_0.pcascodeupm_0.o1.t10 vss 0.16fF
C653 ldomc_0.otaldom_0.pcascodeupm_0.o1.t12 vss 0.16fF
C654 ldomc_0.otaldom_0.pcascodeupm_0.o1.t14 vss 0.16fF
C655 ldomc_0.otaldom_0.pcascodeupm_0.o1.t8 vss 0.16fF
C656 ldomc_0.otaldom_0.pcascodeupm_0.o1.t15 vss 0.16fF
C657 ldomc_0.otaldom_0.pcascodeupm_0.o1.t13 vss 0.16fF
C658 ldomc_0.otaldom_0.pcascodeupm_0.o1.t9 vss 0.16fF
C659 ldomc_0.otaldom_0.pcascodeupm_0.o1.t6 vss 0.16fF
C660 ldomc_0.otaldom_0.pcascodeupm_0.o1.t7 vss 0.16fF
C661 ldomc_0.otaldom_0.pcascodeupm_0.o1.t2 vss 0.16fF
C662 ldomc_0.otaldom_0.pcascodeupm_0.o1.t0 vss 0.16fF
C663 out.t61 vss 0.31fF
C664 out.t57 vss 0.31fF
C665 out.t31 vss 0.31fF
C666 out.t23 vss 0.31fF
C667 out.t65 vss 0.31fF
C668 out.t63 vss 0.31fF
C669 out.t44 vss 0.31fF
C670 out.t36 vss 0.31fF
C671 out.t48 vss 0.31fF
C672 out.t41 vss 0.31fF
C673 out.t29 vss 0.31fF
C674 out.t47 vss 0.31fF
C675 out.t59 vss 0.31fF
C676 out.t32 vss 0.31fF
C677 out.t35 vss 0.31fF
C678 out.t55 vss 0.31fF
C679 out.t53 vss 0.31fF
C680 out.t26 vss 0.31fF
C681 out.t38 vss 0.31fF
C682 out.t51 vss 0.31fF
C683 out.t24 vss 0.31fF
C684 out.t43 vss 0.31fF
C685 out.t1 vss 0.10fF
C686 out.t0 vss 0.07fF
C687 out.t14 vss 2.83fF
C688 out.t16 vss 2.83fF
C689 out.t10 vss 2.83fF
C690 out.t11 vss 2.83fF
C691 out.t13 vss 2.83fF
C692 out.t2 vss 2.83fF
C693 out.t4 vss 2.83fF
C694 out.t18 vss 2.83fF
C695 out.t7 vss 2.83fF
C696 out.t9 vss 3.31fF
C697 out.t8 vss 2.83fF
C698 out.t3 vss 2.83fF
C699 out.t17 vss 2.83fF
C700 out.t12 vss 2.83fF
C701 out.t6 vss 2.83fF
C702 out.t5 vss 2.83fF
C703 out.t20 vss 2.83fF
C704 out.t21 vss 2.83fF
C705 out.t19 vss 2.83fF
C706 out.t15 vss 3.31fF
C707 out.t69 vss 3.91fF
C708 out.t77 vss 3.99fF
C709 out.t67 vss 3.99fF
C710 out.t74 vss 3.99fF
C711 out.t73 vss 3.90fF
C712 out.t81 vss 3.91fF
C713 out.t78 vss 3.99fF
C714 out.t68 vss 3.99fF
C715 out.t76 vss 3.99fF
C716 out.t75 vss 3.90fF
C717 out.t72 vss 3.91fF
C718 out.t84 vss 3.99fF
C719 out.t70 vss 3.99fF
C720 out.t80 vss 3.99fF
C721 out.t79 vss 3.90fF
C722 out.t66 vss 3.91fF
C723 out.t85 vss 3.99fF
C724 out.t71 vss 3.99fF
C725 out.t83 vss 3.99fF
C726 out.t82 vss 4.28fF
C727 out.t40 vss 0.31fF
C728 out.t52 vss 0.31fF
C729 out.t33 vss 0.31fF
C730 out.t25 vss 0.31fF
C731 out.t27 vss 0.31fF
C732 out.t45 vss 0.31fF
C733 out.t60 vss 0.31fF
C734 out.t34 vss 0.31fF
C735 out.t37 vss 0.31fF
C736 out.t56 vss 0.31fF
C737 out.t46 vss 0.31fF
C738 out.t39 vss 0.31fF
C739 out.t54 vss 0.31fF
C740 out.t28 vss 0.31fF
C741 out.t50 vss 0.31fF
C742 out.t42 vss 0.31fF
C743 out.t30 vss 0.31fF
C744 out.t49 vss 0.31fF
C745 out.t22 vss 0.31fF
C746 out.t64 vss 0.31fF
C747 out.t62 vss 0.31fF
C748 out.t58 vss 0.31fF
C749 vdd.t52 vss 0.57fF
C750 vdd.t41 vss 0.57fF
C751 vdd.t74 vss 0.57fF
C752 vdd.t91 vss 0.57fF
C753 vdd.t229 vss 2.01fF
C754 vdd.t89 vss 0.57fF
C755 vdd.t230 vss 0.57fF
C756 vdd.t231 vss 0.57fF
C757 vdd.t40 vss 0.57fF
C758 vdd.t93 vss 0.57fF
C759 vdd.t96 vss 0.57fF
C760 vdd.t51 vss 0.57fF
C761 vdd.t86 vss 0.57fF
C762 vdd.t98 vss 0.57fF
C763 vdd.t67 vss 0.57fF
C764 vdd.t57 vss 0.57fF
C765 vdd.t313 vss 0.17fF
C766 vdd.t297 vss 0.22fF
C767 vdd.t305 vss 0.15fF
C768 vdd.t318 vss 0.01fF
C769 vdd.t332 vss 0.07fF
C770 vdd.t115 vss 0.05fF
C771 vdd.t103 vss 0.05fF
C772 vdd.t287 vss 0.22fF
C773 vdd.t130 vss 0.23fF
C774 vdd.t133 vss 0.05fF
C775 vdd.t131 vss 0.05fF
C776 vdd.t132 vss 0.06fF
C777 vdd.t329 vss 0.07fF
C778 vdd.t122 vss 0.10fF
C779 vdd.t286 vss 0.22fF
C780 vdd.t108 vss 0.31fF
C781 vdd.t331 vss 0.23fF
C782 vdd.t110 vss 0.29fF
C783 vdd.t111 vss 0.05fF
C784 vdd.t109 vss 0.05fF
C785 vdd.t112 vss 0.07fF
C786 vdd.t285 vss 0.07fF
C787 vdd.t288 vss 0.06fF
C788 vdd.t128 vss 0.22fF
C789 vdd.t135 vss 0.05fF
C790 vdd.t129 vss 0.05fF
C791 vdd.t327 vss 0.31fF
C792 vdd.t328 vss 0.23fF
C793 vdd.t136 vss 0.07fF
C794 vdd.t283 vss 0.09fF
C795 vdd.t127 vss 0.05fF
C796 vdd.t137 vss 0.05fF
C797 vdd.t126 vss 0.07fF
C798 vdd.t316 vss 0.07fF
C799 vdd.t334 vss 0.22fF
C800 vdd.t107 vss 0.05fF
C801 vdd.t121 vss 0.05fF
C802 vdd.t106 vss 0.08fF
C803 vdd.t323 vss 0.07fF
C804 vdd.t289 vss 0.31fF
C805 vdd.t320 vss 0.02fF
C806 vdd.t212 vss 0.18fF
C807 vdd.t294 vss 0.13fF
C808 vdd.t360 vss 0.09fF
C809 vdd.t308 vss 0.23fF
C810 vdd.t366 vss 0.09fF
C811 vdd.t387 vss 0.02fF
C812 vdd.t303 vss 0.21fF
C813 vdd.t353 vss 0.11fF
C814 vdd.t299 vss 0.15fF
C815 vdd.t372 vss 0.25fF
C816 vdd.t56 vss 7.01fF
C817 vdd.t82 vss 2.86fF
C818 vdd.t295 vss 0.40fF
C819 vdd.t381 vss 0.40fF
C820 vdd.t80 vss 0.08fF
C821 vdd.t362 vss 0.40fF
C822 vdd.t368 vss 0.31fF
C823 vdd.t314 vss 0.30fF
C824 vdd.t357 vss 0.31fF
C825 vdd.t310 vss 0.31fF
C826 vdd.t306 vss 0.31fF
C827 vdd.t309 vss 0.31fF
C828 vdd.t377 vss 0.05fF
C829 vdd.t298 vss 0.38fF
C830 vdd.t383 vss 0.30fF
C831 vdd.t302 vss 0.09fF
C832 vdd.t375 vss 0.31fF
C833 vdd.t291 vss 0.31fF
C834 vdd.t364 vss 0.31fF
C835 vdd.t374 vss 0.31fF
C836 vdd.t370 vss 0.32fF
C837 vdd.t386 vss 0.02fF
C838 vdd.t378 vss 0.02fF
C839 vdd.t384 vss 0.02fF
C840 vdd.t376 vss 0.02fF
C841 vdd.t365 vss 0.02fF
C842 vdd.t185 vss 0.24fF
C843 vdd.t189 vss 0.24fF
C844 vdd.t187 vss 0.02fF
C845 vdd.t188 vss 0.01fF
C846 vdd.t358 vss 0.02fF
C847 vdd.t380 vss 0.02fF
C848 vdd.t373 vss 0.02fF
C849 vdd.t382 vss 0.02fF
C850 vdd.t388 vss 0.02fF
C851 vdd.t354 vss 0.02fF
C852 vdd.t361 vss 0.02fF
C853 vdd.t224 vss 0.24fF
C854 vdd.t211 vss 0.24fF
C855 vdd.t367 vss 0.02fF
C856 vdd.t356 vss 0.02fF
C857 vdd.t363 vss 0.02fF
C858 vdd.t369 vss 0.02fF
C859 vdd.t186 vss 0.40fF
C860 vdd.t190 vss 0.07fF
C861 vdd.t385 vss 0.31fF
C862 vdd.t379 vss 0.31fF
C863 vdd.t311 vss 0.06fF
C864 vdd.t371 vss 0.40fF
C865 vdd.t359 vss 0.40fF
C866 vdd.t83 vss 0.25fF
C867 vdd.t301 vss 0.06fF
C868 vdd.t355 vss 0.17fF
C869 vdd.t304 vss 0.06fF
C870 vdd.t225 vss 0.15fF
C871 vdd.t296 vss -1.81fF
C872 vdd.t319 vss 0.21fF
C873 vdd.t324 vss 0.21fF
C874 vdd.t284 vss 0.23fF
C875 vdd.t120 vss 0.23fF
C876 vdd.t335 vss 0.31fF
C877 vdd.t118 vss 0.22fF
C878 vdd.t119 vss 0.05fF
C879 vdd.t117 vss 0.05fF
C880 vdd.t116 vss 0.07fF
C881 vdd.t134 vss 0.23fF
C882 vdd.t104 vss 0.09fF
C883 vdd.t105 vss 0.05fF
C884 vdd.t113 vss 0.05fF
C885 vdd.t330 vss 0.08fF
C886 vdd.t124 vss 0.22fF
C887 vdd.t125 vss 0.05fF
C888 vdd.t123 vss 0.05fF
C889 vdd.t290 vss 0.07fF
C890 vdd.t326 vss 0.07fF
C891 vdd.t315 vss 0.23fF
C892 vdd.t114 vss 0.31fF
C893 vdd.t102 vss 0.22fF
C894 vdd.t333 vss 0.09fF
C895 vdd.t317 vss 0.31fF
C896 vdd.t321 vss 0.23fF
C897 vdd.t322 vss 0.33fF
C898 vdd.t307 vss 0.17fF
C899 vdd.t312 vss 0.17fF
C900 vdd.t292 vss 0.17fF
C901 vdd.t293 vss 0.22fF
C902 vdd.t300 vss 0.17fF
C903 vdd.t220 vss 0.07fF
C904 vdd.t27 vss 0.32fF
C905 vdd.t336 vss 0.08fF
C906 vdd.t0 vss 0.40fF
C907 vdd.t269 vss 0.06fF
C908 vdd.t28 vss 0.09fF
C909 vdd.t341 vss 7.01fF
C910 vdd.t339 vss 2.86fF
C911 vdd.t263 vss -0.80fF
C912 vdd.t249 vss -1.82fF
C913 vdd.t181 vss 0.18fF
C914 vdd.t195 vss 0.15fF
C915 vdd.t266 vss 0.13fF
C916 vdd.t251 vss 0.23fF
C917 vdd.t34 vss 0.09fF
C918 vdd.t261 vss 0.06fF
C919 vdd.t18 vss 0.17fF
C920 vdd.t2 vss 0.02fF
C921 vdd.t260 vss 0.21fF
C922 vdd.t16 vss 0.11fF
C923 vdd.t259 vss 0.15fF
C924 vdd.t14 vss 0.25fF
C925 vdd.t337 vss 0.25fF
C926 vdd.t22 vss 0.40fF
C927 vdd.t6 vss 0.40fF
C928 vdd.t24 vss 0.40fF
C929 vdd.t252 vss 0.06fF
C930 vdd.t20 vss 0.31fF
C931 vdd.t257 vss 0.30fF
C932 vdd.t8 vss 0.31fF
C933 vdd.t270 vss 0.31fF
C934 vdd.t25 vss 0.31fF
C935 vdd.t254 vss 0.31fF
C936 vdd.t4 vss 0.31fF
C937 vdd.t271 vss 0.31fF
C938 vdd.t10 vss 0.05fF
C939 vdd.t258 vss 0.38fF
C940 vdd.t30 vss 0.30fF
C941 vdd.t264 vss 0.09fF
C942 vdd.t12 vss 0.31fF
C943 vdd.t250 vss 0.31fF
C944 vdd.t32 vss 0.31fF
C945 vdd.t23 vss 0.31fF
C946 vdd.t243 vss 0.14fF
C947 vdd.t247 vss 0.14fF
C948 vdd.t352 vss 0.14fF
C949 vdd.t350 vss 0.14fF
C950 vdd.t274 vss 0.14fF
C951 vdd.t277 vss 0.14fF
C952 vdd.t346 vss 0.03fF
C953 vdd.t344 vss 0.04fF
C954 vdd.t281 vss 0.14fF
C955 vdd.t273 vss 0.14fF
C956 vdd.t348 vss -2.79fF
C957 vdd.t347 vss 0.03fF
C958 vdd.t160 vss 0.04fF
C959 vdd.t143 vss 0.05fF
C960 vdd.t145 vss 0.05fF
C961 vdd.t155 vss 0.05fF
C962 vdd.t159 vss 0.05fF
C963 vdd.t171 vss 0.05fF
C964 vdd.t165 vss 0.05fF
C965 vdd.t170 vss 0.17fF
C966 vdd.t140 vss 0.17fF
C967 vdd.t153 vss 0.05fF
C968 vdd.t141 vss 0.05fF
C969 vdd.t244 vss 0.17fF
C970 vdd.t242 vss 0.17fF
C971 vdd.t152 vss 0.17fF
C972 vdd.t164 vss 0.04fF
C973 vdd.t154 vss 0.05fF
C974 vdd.t158 vss 0.17fF
C975 vdd.t142 vss 0.17fF
C976 vdd.t144 vss 0.17fF
C977 vdd.t168 vss 0.04fF
C978 vdd.t169 vss 0.05fF
C979 vdd.t161 vss 0.05fF
C980 vdd.t163 vss 0.05fF
C981 vdd.t147 vss 0.05fF
C982 vdd.t149 vss 0.05fF
C983 vdd.t173 vss 0.05fF
C984 vdd.t175 vss 0.05fF
C985 vdd.t167 vss 0.05fF
C986 vdd.t166 vss 0.17fF
C987 vdd.t150 vss 0.17fF
C988 vdd.t151 vss 0.05fF
C989 vdd.t157 vss 0.05fF
C990 vdd.t256 vss 0.17fF
C991 vdd.t268 vss 0.22fF
C992 vdd.t267 vss 0.17fF
C993 vdd.t272 vss 0.17fF
C994 vdd.t255 vss 0.17fF
C995 vdd.t253 vss 0.17fF
C996 vdd.t265 vss 0.22fF
C997 vdd.t262 vss 0.17fF
C998 vdd.t241 vss 0.17fF
C999 vdd.t248 vss 0.17fF
C1000 vdd.t156 vss 0.17fF
C1001 vdd.t174 vss 0.04fF
C1002 vdd.t172 vss 0.05fF
C1003 vdd.t148 vss 0.17fF
C1004 vdd.t146 vss 0.17fF
C1005 vdd.t162 vss 0.17fF
C1006 vdd.t280 vss 0.03fF
C1007 vdd.t279 vss 0.14fF
C1008 vdd.t351 vss 0.14fF
C1009 vdd.t349 vss 0.14fF
C1010 vdd.t276 vss 0.04fF
C1011 vdd.t278 vss 0.03fF
C1012 vdd.t345 vss 0.14fF
C1013 vdd.t325 vss 0.14fF
C1014 vdd.t282 vss 0.14fF
C1015 vdd.t275 vss 0.14fF
C1016 vdd.t246 vss 0.14fF
C1017 vdd.t245 vss 0.14fF
C1018 vdd.t177 vss 0.40fF
C1019 vdd.t33 vss 0.02fF
C1020 vdd.t178 vss 0.02fF
C1021 vdd.t176 vss 0.24fF
C1022 vdd.t219 vss 0.24fF
C1023 vdd.t179 vss 0.01fF
C1024 vdd.t31 vss 0.02fF
C1025 vdd.t13 vss 0.02fF
C1026 vdd.t5 vss 0.02fF
C1027 vdd.t11 vss 0.02fF
C1028 vdd.t9 vss 0.02fF
C1029 vdd.t26 vss 0.02fF
C1030 vdd.t15 vss 0.02fF
C1031 vdd.t1 vss 0.02fF
C1032 vdd.t3 vss 0.02fF
C1033 vdd.t17 vss 0.02fF
C1034 vdd.t29 vss 0.02fF
C1035 vdd.t194 vss 0.24fF
C1036 vdd.t180 vss 0.24fF
C1037 vdd.t35 vss 0.02fF
C1038 vdd.t19 vss 0.02fF
C1039 vdd.t7 vss 0.02fF
C1040 vdd.t21 vss 0.02fF
C1041 vdd.t200 vss 0.34fF
C1042 vdd.t239 vss 0.05fF
C1043 vdd.t202 vss 0.05fF
C1044 vdd.t338 vss 0.05fF
C1045 vdd.t238 vss 0.48fF
C1046 vdd.t199 vss 0.48fF
C1047 vdd.t240 vss 0.05fF
C1048 vdd.t201 vss 0.05fF
C1049 vdd.t203 vss 0.12fF
C1050 vdd.t100 vss 0.15fF
C1051 vdd.t138 vss 0.97fF
C1052 vdd.t204 vss 1.09fF
C1053 vdd.t101 vss 0.01fF
C1054 vdd.t139 vss 0.01fF
C1055 vdd.t340 vss 0.05fF
C1056 vdd.t236 vss 0.05fF
C1057 vdd.t207 vss 0.05fF
C1058 vdd.t343 vss 0.05fF
C1059 vdd.t342 vss 0.05fF
C1060 vdd.t235 vss 0.48fF
C1061 vdd.t205 vss 0.48fF
C1062 vdd.t237 vss 0.05fF
C1063 vdd.t206 vss 0.05fF
C1064 vdd.t55 vss 0.57fF
C1065 vdd.t45 vss 0.57fF
C1066 vdd.t76 vss 0.57fF
C1067 vdd.t92 vss 0.57fF
C1068 vdd.t90 vss 0.57fF
C1069 vdd.t233 vss 0.57fF
C1070 vdd.t234 vss 0.57fF
C1071 vdd.t79 vss 0.57fF
C1072 vdd.t77 vss 0.57fF
C1073 vdd.t36 vss 0.44fF
C1074 vdd.t217 vss 0.57fF
C1075 vdd.t218 vss 0.57fF
C1076 vdd.t64 vss 0.57fF
C1077 vdd.t216 vss 2.01fF
C1078 vdd.t232 vss 2.01fF
C1079 vdd.t78 vss 0.57fF
C1080 vdd.t75 vss 0.57fF
C1081 vdd.t65 vss 0.57fF
C1082 vdd.t81 vss 0.57fF
C1083 vdd.t58 vss 0.57fF
C1084 vdd.t48 vss 0.57fF
C1085 vdd.t44 vss 0.57fF
C1086 vdd.t69 vss 0.57fF
C1087 vdd.t209 vss 0.57fF
C1088 vdd.t210 vss 0.57fF
C1089 vdd.t61 vss 0.57fF
C1090 vdd.t39 vss 0.44fF
C1091 vdd.t208 vss 2.01fF
C1092 bandgapmd_0.otam_1.nmosrm_0.outn.t10 vss 0.02fF
C1093 bandgapmd_0.otam_1.nmosrm_0.outn.t12 vss 0.02fF
C1094 bandgapmd_0.otam_1.nmosrm_0.outn.t7 vss 0.02fF
C1095 bandgapmd_0.otam_1.nmosrm_0.outn.t4 vss 0.02fF
C1096 bandgapmd_0.otam_1.nmosrm_0.outn.t6 vss 0.02fF
C1097 bandgapmd_0.otam_1.nmosrm_0.outn.t8 vss 0.02fF
C1098 bandgapmd_0.otam_1.nmosrm_0.outn.t15 vss 0.02fF
C1099 bandgapmd_0.otam_1.nmosrm_0.outn.t1 vss 0.02fF
C1100 bandgapmd_0.otam_1.nmosrm_0.outn.t2 vss 0.02fF
C1101 bandgapmd_0.otam_1.nmosrm_0.outn.t9 vss 0.02fF
C1102 bandgapmd_0.otam_1.nmosrm_0.outn.t0 vss 0.02fF
C1103 bandgapmd_0.otam_1.nmosrm_0.outn.t13 vss 0.02fF
C1104 bandgapmd_0.otam_1.nmosrm_0.outn.t11 vss 0.02fF
C1105 bandgapmd_0.otam_1.nmosrm_0.outn.t14 vss 0.02fF
C1106 bandgapmd_0.otam_1.nmosrm_0.outn.t3 vss 0.02fF
C1107 bandgapmd_0.otam_1.nmosrm_0.outn.t5 vss 0.02fF
C1108 bandgapmd_0.otam_1.nmosrm_0.outn.t18 vss 0.03fF
C1109 bandgapmd_0.otam_1.nmosrm_0.outn.t17 vss 0.03fF
C1110 bandgapmd_0.otam_1.nmosrm_0.outn.t20 vss 0.03fF
C1111 bandgapmd_0.otam_1.nmosrm_0.outn.t22 vss 0.03fF
C1112 bandgapmd_0.otam_1.nmosrm_0.outn.t19 vss 0.03fF
C1113 bandgapmd_0.otam_1.nmosrm_0.outn.t21 vss 0.03fF
C1114 bandgapmd_0.otam_1.nmosrm_0.outn.t23 vss 0.03fF
C1115 bandgapmd_0.otam_1.nmosrm_0.outn.t16 vss 0.03fF
C1116 bandgapmd_0.otam_1.nmosrm_0.outn.t28 vss 0.07fF
C1117 bandgapmd_0.otam_1.nmosrm_0.outn.t25 vss 0.07fF
C1118 bandgapmd_0.otam_1.nmosrm_0.outn.t24 vss 0.07fF
C1119 bandgapmd_0.otam_1.nmosrm_0.outn.t32 vss 0.07fF
C1120 bandgapmd_0.otam_1.nmosrm_0.outn.t30 vss 0.07fF
C1121 bandgapmd_0.otam_1.nmosrm_0.outn.t31 vss 0.07fF
C1122 bandgapmd_0.otam_1.nmosrm_0.outn.t29 vss 0.07fF
C1123 bandgapmd_0.otam_1.nmosrm_0.outn.t27 vss 0.07fF
C1124 bandgapmd_0.otam_1.nmosrm_0.outn.t26 vss 0.07fF
C1125 bandgapmd_0.otam_1.nmosrm_0.outn.t33 vss 0.07fF
.ends

