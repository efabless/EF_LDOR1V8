VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_LDOR01
  CLASS BLOCK ;
  FOREIGN EF_LDOR01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END EF_LDOR01
END LIBRARY

