** sch_path: /home/ahmedreda/Project/AR_BGR/testbench/full_ldo/fullldox_v2-tb/startup.sch
**.subckt startup
C3 vo net1 47u m=1
R4 net1 vss 0.1 m=1
R5 vo net2 18 m=1
Vl net2 vss 0
.save i(vl)
x1 biasldo biasbgr vss vss vss vdd vss vss vss vss vss vss vss vss vss vss vss vss vo vdd vss fullldom

vdd2 vdd1 vss PWL(0 0 1u 0 2u 3.3)
.save i(vdd2)
vss2 vss GND 0
.save i(vss2)
Vbias net3 biasbgr 0
.save i(vbias)
vtot vdd1 vdd 0
.save i(vtot)
R3 net4 vdd 300000 m=1
Vbiasldo net4 biasldo 0
.save i(vbiasldo)
R2 net3 vdd 450000 m=1
**** begin user architecture code


.lib /home/ahmedreda/PDK/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.include fullldom.spice



.options RSHUNT=1e15
.options savecurrents
.option TEMP=27
.option TNOM=27
.control
**set filetype=binary
set filetype=ascii
set color0=white
set color1=black
set color3=blue
set xbrushwidth=5
save all
OP
tran 0.1u 0.6m 0.1u
plot  vdd vo
.endc





.GLOBAL GND
.end
